* NGSPICE file created from adc_top.ext - technology: sky130A

.subckt adc_top_postlayout result_out[0] result_out[1] result_out[2] result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8] result_out[9] result_out[10] result_out[11] result_out[12] result_out[13] result_out[14] result_out[15] 
+ VDD VSS conversion_finished_out rst_n start_conversion_in clk_vcm inp_analog inn_analog
+ config_1_in[0] config_1_in[1] config_1_in[2] config_1_in[3] config_1_in[4] config_1_in[5] config_1_in[6] config_1_in[7] config_1_in[8] config_1_in[9]
+ config_1_in[10] config_1_in[11] config_1_in[12] config_1_in[13] config_1_in[14] config_1_in[15] 
+ config_2_in[0] config_2_in[1] config_2_in[2] config_2_in[3] config_2_in[4] config_2_in[5] config_2_in[6] config_2_in[7] config_2_in[8] config_2_in[9] 
+ config_2_in[10] config_2_in[11] config_2_in[12] config_2_in[13] config_2_in[14] config_2_in[15] 
+ dummypin[0] dummypin[10] dummypin[11] dummypin[12] dummypin[13] dummypin[14] dummypin[15] dummypin[1] dummypin[2] dummypin[3] dummypin[4] dummypin[5] dummypin[6] dummypin[7] dummypin[8] dummypin[9]
+ ctopp ctopn vcm clk_dig clk_comp clk_ena ndecision_finish comp_latch
C_D0 VSS a_7717_14735# 0.01fF
C_D1 VSS a_12447_16143# 0.01fF
C_D10 VSS a_7109_29423# 0.01fF
C_D100 VSS _1184_.A2 0.01fF
C_D1000 VSS a_2007_25597# 0.01fF
C_D1001 VSS _1154_.A 0.01fF
C_D1002 VSS _1224_.X 0.01fF
C_D1003 VSS a_4259_31375# 0.01fF
C_D1004 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D1005 VSS a_2263_43719# 0.01fF
C_D1006 VSS a_9411_2215# 0.01fF
C_D1007 VSS pmat.sw 0.01fF
C_D1008 VSS a_11149_40188# 0.01fF
C_D1009 VSS a_4383_7093# 0.01fF
C_D101 VSS a_12263_50959# 0.01fF
C_D1010 VSS cgen.dlycontrol4_in[2] 0.01fF
C_D1011 VSS a_24591_28327# 0.01fF
C_D1012 VSS a_37820_30485# 0.01fF
C_D1013 VSS a_13091_7655# 0.01fF
C_D1014 VSS a_13459_28111# 0.01fF
C_D1015 VSS _1224_.X 0.01fF
C_D1016 VSS pmat.en_bit_n[0] 0.01fF
C_D1017 VSS a_1957_43567# 0.01fF
C_D1018 VSS _1179_.X 0.01fF
C_D1019 VSS a_40837_46261# 0.01fF
C_D102 VSS a_6787_47607# 0.01fF
C_D1020 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D1021 VSS a_10515_13967# 0.01fF
C_D1022 VSS a_2407_49289# 0.01fF
C_D1023 VSS a_18563_27791# 0.01fF
C_D1024 VSS a_21279_48999# 0.01fF
C_D1025 VSS a_40837_46261# 0.01fF
C_D1026 VSS a_1899_35051# 0.01fF
C_D1027 VSS a_4383_7093# 0.01fF
C_D1028 VSS a_30663_50087# 0.01fF
C_D1029 VSS a_24407_31375# 0.01fF
C_D103 VSS a_9963_28111# 0.01fF
C_D1030 VSS a_11067_16359# 0.01fF
C_D1031 VSS a_17139_30503# 0.01fF
C_D1032 VSS _1154_.A 0.01fF
C_D1033 VSS a_25879_31591# 0.01fF
C_D1034 VSS cgen.dlycontrol4_in[5] 0.01fF
C_D1035 VSS _1192_.A2 0.01fF
C_D1036 VSS a_2411_43301# 0.01fF
C_D1037 VSS a_11435_58791# 0.01fF
C_D1038 VSS a_10055_31591# 0.01fF
C_D1039 VSS nmat.col_n[30] 0.01fF
C_D104 VSS a_10239_14183# 0.01fF
C_D1040 VSS a_5081_53135# 0.01fF
C_D1041 VSS a_4075_68583# 0.01fF
C_D1042 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D1043 VSS _1194_.A2 0.01fF
C_D1044 VSS a_13091_52047# 0.01fF
C_D1045 VSS a_4128_64391# 0.01fF
C_D1046 VSS a_22153_37179# 0.01fF
C_D1047 VSS a_2407_49289# 0.01fF
C_D1048 VSS a_11067_27239# 0.01fF
C_D1049 VSS a_29937_31055# 0.01fF
C_D105 VSS a_4075_31591# 0.01fF
C_D1050 VSS nmat.sw 0.01fF
C_D1051 VSS a_11067_16359# 0.01fF
C_D1052 VSS a_10515_61839# 0.01fF
C_D1053 VSS a_33423_47695# 0.01fF
C_D1054 VSS a_2411_43301# 0.01fF
C_D1055 VSS _1196_.B1 0.01fF
C_D1056 VSS a_2411_43301# 0.01fF
C_D1057 VSS a_11067_16359# 0.01fF
C_D1058 VSS a_4075_50087# 0.01fF
C_D1059 VSS a_4719_30287# 0.01fF
C_D106 VSS _1194_.A2 0.01fF
C_D1060 VSS _1224_.X 0.01fF
C_D1061 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D1062 VSS a_10883_3303# 0.01fF
C_D1063 VSS _1196_.B1 0.01fF
C_D1064 VSS a_2419_53351# 0.01fF
C_D1065 VSS a_25879_31591# 0.01fF
C_D1066 VSS a_14887_46377# 0.01fF
C_D1067 VSS config_1_in[1] 0.01fF
C_D1068 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D1069 VSS a_10515_61839# 0.01fF
C_D107 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D1070 VSS a_5651_66975# 0.01fF
C_D1071 VSS nmat.col[29] 0.01fF
C_D1072 VSS nmat.col[15] 0.01fF
C_D1073 VSS a_8583_29199# 0.01fF
C_D1074 VSS _1154_.A 0.01fF
C_D1075 VSS nmat.en_bit_n[1] 0.01fF
C_D1076 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D1077 VSS pmat.row_n[8] 0.01fF
C_D1078 VSS a_9963_28111# 0.01fF
C_D1079 VSS a_2007_25597# 0.01fF
C_D108 VSS a_5081_53135# 0.01fF
C_D1080 VSS _1224_.X 0.01fF
C_D1081 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D1082 VSS _1192_.B1 0.01fF
C_D1083 VSS a_11067_64015# 0.01fF
C_D1084 VSS a_7939_31591# 0.01fF
C_D1085 VSS a_33423_47695# 0.01fF
C_D1086 VSS a_6559_33767# 0.01fF
C_D1087 VSS a_2835_13077# 0.01fF
C_D1088 VSS comp_latch 0.01fF
C_D1089 VSS a_6467_29415# 0.01fF
C_D109 VSS pmat.row_n[5] 0.01fF
C_D1090 VSS a_2791_57703# 0.01fF
C_D1091 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D1092 VSS cgen.dlycontrol1_in[2] 0.01fF
C_D1093 VSS _1192_.B1 0.01fF
C_D1094 VSS a_1586_50247# 0.01fF
C_D1095 VSS a_11067_16359# 0.01fF
C_D1096 VSS a_12263_50959# 0.01fF
C_D1097 VSS a_13091_28327# 0.01fF
C_D1098 VSS pmat.rowoff_n[8] 0.01fF
C_D1099 VSS a_6664_26159# 0.01fF
C_D11 VSS _1154_.X 0.01fF
C_D110 VSS a_7109_29423# 0.01fF
C_D1100 VSS a_7717_14735# 0.01fF
C_D1101 VSS pmat.rowoff_n[7] 0.01fF
C_D1102 VSS a_1586_18231# 0.01fF
C_D1103 VSS a_1591_31599# 0.01fF
C_D1104 VSS config_1_in[9] 0.01fF
C_D1105 VSS a_7415_29397# 0.01fF
C_D1106 VSS a_6664_26159# 0.01fF
C_D1107 VSS cgen.dlycontrol3_in[0] 0.01fF
C_D1108 VSS a_11067_64015# 0.01fF
C_D1109 VSS _1196_.B1 0.01fF
C_D111 VSS pmat.row_n[2] 0.01fF
C_D1110 VSS _1183_.A2 0.01fF
C_D1111 VSS a_11067_27239# 0.01fF
C_D1112 VSS a_5651_66975# 0.01fF
C_D1113 VSS cgen.dlycontrol2_in[3] 0.01fF
C_D1114 VSS a_10515_13967# 0.01fF
C_D1115 VSS a_18563_27791# 0.01fF
C_D1116 VSS nmat.rowon_n[7] 0.01fF
C_D1117 VSS a_4075_31591# 0.01fF
C_D1118 VSS clk_ena 0.01fF
C_D1119 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D112 VSS a_13641_23439# 0.01fF
C_D1120 VSS a_13091_28327# 0.01fF
C_D1121 VSS a_1923_61759# 0.01fF
C_D1122 VSS a_14287_70543# 0.01fF
C_D1123 VSS a_22199_30287# 0.01fF
C_D1124 VSS a_17842_27497# 0.01fF
C_D1125 VSS a_2791_57703# 0.01fF
C_D1126 VSS a_1586_18231# 0.01fF
C_D1127 VSS a_1586_50247# 0.01fF
C_D1128 VSS a_31675_47695# 0.01fF
C_D1129 VSS a_31675_47695# 0.01fF
C_D113 VSS a_3615_71631# 0.01fF
C_D1130 VSS config_1_in[8] 0.01fF
C_D1131 VSS nmat.rowon_n[7] 0.01fF
C_D1132 VSS nmat.col[18] 0.01fF
C_D1133 VSS a_2879_57487# 0.01fF
C_D1134 VSS config_1_in[11] 0.01fF
C_D1135 VSS a_10515_13967# 0.01fF
C_D1136 VSS cgen.dlycontrol2_in[4] 0.01fF
C_D1137 VSS a_2419_69455# 0.01fF
C_D1138 VSS clk_ena 0.01fF
C_D1139 VSS _1184_.A2 0.01fF
C_D114 VSS a_13459_28111# 0.01fF
C_D1140 VSS a_2791_57703# 0.01fF
C_D1141 VSS a_6927_30503# 0.01fF
C_D1142 VSS pmat.rowon_n[7] 0.01fF
C_D1143 VSS a_13091_28327# 0.01fF
C_D1144 VSS a_6787_47607# 0.01fF
C_D1145 VSS pmat.col[31] 0.01fF
C_D1146 VSS cgen.dlycontrol3_in[1] 0.01fF
C_D1147 VSS a_1586_50247# 0.01fF
C_D1148 VSS clk_ena 0.01fF
C_D1149 VSS a_5651_66975# 0.01fF
C_D115 VSS _1224_.X 0.01fF
C_D1150 VSS a_2263_43719# 0.01fF
C_D1151 VSS ANTENNA_fanout52_A.DIODE 0.01fF
C_D1152 VSS nmat.col[26] 0.01fF
C_D1153 VSS nmat.col[31] 0.01fF
C_D1154 VSS clk_ena 0.01fF
C_D1155 VSS a_4075_50087# 0.01fF
C_D1156 VSS a_8583_29199# 0.01fF
C_D1157 VSS _1179_.X 0.01fF
C_D1158 VSS pmat.row_n[6] 0.01fF
C_D1159 VSS a_4719_30287# 0.01fF
C_D116 VSS a_11067_30287# 0.01fF
C_D1160 VSS a_6787_47607# 0.01fF
C_D1161 VSS nmat.sw 0.01fF
C_D1162 VSS _1187_.A2 0.01fF
C_D1163 VSS nmat.col_n[12] 0.01fF
C_D1164 VSS nmat.col[24] 0.01fF
C_D1165 VSS a_28915_50959# 0.01fF
C_D1166 VSS pmat.row_n[10] 0.01fF
C_D1167 VSS config_2_in[13] 0.01fF
C_D1168 VSS a_9411_2215# 0.01fF
C_D1169 VSS a_9963_13967# 0.01fF
C_D117 VSS a_10515_13967# 0.01fF
C_D1170 VSS _1179_.X 0.01fF
C_D1171 VSS a_30663_50087# 0.01fF
C_D1172 VSS a_2411_43301# 0.01fF
C_D1173 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D1174 VSS a_30111_47911# 0.01fF
C_D1175 VSS nmat.rowon_n[7] 0.01fF
C_D1176 VSS _1194_.B1 0.01fF
C_D1177 VSS a_5651_66975# 0.01fF
C_D1178 VSS a_5351_19913# 0.01fF
C_D1179 VSS a_4719_30287# 0.01fF
C_D118 VSS a_1769_13103# 0.01fF
C_D1180 VSS a_10883_3303# 0.01fF
C_D1181 VSS a_1923_31743# 0.01fF
C_D1182 VSS a_2407_49289# 0.01fF
C_D1183 VSS nmat.col_n[19] 0.01fF
C_D1184 VSS a_5363_33551# 0.01fF
C_D1185 VSS pmat.rowon_n[7] 0.01fF
C_D1186 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D1187 VSS pmat.rowon_n[8] 0.01fF
C_D1188 VSS a_7415_29397# 0.01fF
C_D1189 VSS a_30571_50959# 0.01fF
C_D119 VSS a_4383_7093# 0.01fF
C_D1190 VSS a_4383_7093# 0.01fF
C_D1191 VSS a_1923_61759# 0.01fF
C_D1192 VSS a_6283_31591# 0.01fF
C_D1193 VSS pmat.rowoff_n[15] 0.01fF
C_D1194 VSS a_5351_19913# 0.01fF
C_D1195 VSS a_10515_13967# 0.01fF
C_D1196 VSS a_2411_43301# 0.01fF
C_D1197 VSS nmat.col_n[10] 0.01fF
C_D1198 VSS a_30571_50959# 0.01fF
C_D1199 VSS ANTENNA__1183__B1.DIODE 0.01fF
C_D12 VSS _1154_.X 0.01fF
C_D120 VSS a_10239_14183# 0.01fF
C_D1200 VSS a_10055_31591# 0.01fF
C_D1201 VSS a_13275_48783# 0.01fF
C_D1202 VSS a_9963_13967# 0.01fF
C_D1203 VSS _1194_.B1 0.01fF
C_D1204 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D1205 VSS a_30111_47911# 0.01fF
C_D1206 VSS a_24407_31375# 0.01fF
C_D1207 VSS a_6283_31591# 0.01fF
C_D1208 VSS nmat.rowon_n[14] 0.01fF
C_D1209 VSS a_25879_31591# 0.01fF
C_D121 VSS a_7109_29423# 0.01fF
C_D1210 VSS cgen.start_conv_in 0.01fF
C_D1211 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D1212 VSS a_17139_30503# 0.01fF
C_D1213 VSS a_28915_50959# 0.01fF
C_D1214 VSS a_1923_61759# 0.01fF
C_D1215 VSS pmat.row_n[14] 0.01fF
C_D1216 VSS a_1586_50247# 0.01fF
C_D1217 VSS a_25695_28111# 0.01fF
C_D1218 VSS a_21739_29415# 0.01fF
C_D1219 VSS a_6283_31591# 0.01fF
C_D122 VSS a_1586_50247# 0.01fF
C_D1220 VSS comp_latch 0.01fF
C_D1221 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D1222 VSS a_11067_30287# 0.01fF
C_D1223 VSS a_11317_36924# 0.01fF
C_D1224 VSS a_30571_50959# 0.01fF
C_D1225 VSS a_1899_35051# 0.01fF
C_D1226 VSS a_1923_61759# 0.01fF
C_D1227 VSS nmat.sw 0.01fF
C_D1228 VSS a_11067_30287# 0.01fF
C_D1229 VSS cgen.dlycontrol4_in[5] 0.01fF
C_D123 VSS a_1923_31743# 0.01fF
C_D1230 VSS a_2263_43719# 0.01fF
C_D1231 VSS a_4075_31591# 0.01fF
C_D1232 VSS pmat.en_bit_n[2] 0.01fF
C_D1233 VSS a_11317_36924# 0.01fF
C_D1234 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D1235 VSS _1194_.B1 0.01fF
C_D1236 VSS a_33423_47695# 0.01fF
C_D1237 VSS a_4383_7093# 0.01fF
C_D1238 VSS _1184_.A2 0.01fF
C_D1239 VSS nmat.sw 0.01fF
C_D124 VSS pmat.row_n[8] 0.01fF
C_D1240 VSS pmat.row_n[4] 0.01fF
C_D1241 VSS a_16311_28327# 0.01fF
C_D1242 VSS a_4075_31591# 0.01fF
C_D1243 VSS a_11067_27239# 0.01fF
C_D1244 VSS a_3339_59879# 0.01fF
C_D1245 VSS a_8491_47911# 0.01fF
C_D1246 VSS a_30111_47911# 0.01fF
C_D1247 VSS a_22199_30287# 0.01fF
C_D1248 VSS a_2046_30184# 0.01fF
C_D1249 VSS cgen.dlycontrol4_in[3] 0.01fF
C_D125 VSS a_14887_46377# 0.01fF
C_D1250 VSS _1196_.B1 0.01fF
C_D1251 VSS a_2411_43301# 0.01fF
C_D1252 VSS a_13091_52047# 0.01fF
C_D1253 VSS a_24407_31375# 0.01fF
C_D1254 VSS a_1957_43567# 0.01fF
C_D1255 VSS config_2_in[5] 0.01fF
C_D1256 VSS a_15667_27239# 0.01fF
C_D1257 VSS _1224_.X 0.01fF
C_D1258 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D1259 VSS a_2046_30184# 0.01fF
C_D126 VSS a_16311_28327# 0.01fF
C_D1260 VSS a_8491_47911# 0.01fF
C_D1261 VSS a_4075_31591# 0.01fF
C_D1262 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D1263 VSS a_2879_57487# 0.01fF
C_D1264 VSS pmat.rowon_n[7] 0.01fF
C_D1265 VSS clk_dig 0.01fF
C_D1266 VSS a_6559_33767# 0.01fF
C_D1267 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D1268 VSS a_31675_47695# 0.01fF
C_D1269 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D127 VSS comp_latch 0.01fF
C_D1270 VSS a_10873_38517# 0.01fF
C_D1271 VSS a_4259_73807# 0.01fF
C_D1272 VSS a_38851_28327# 0.01fF
C_D1273 VSS a_13091_52047# 0.01fF
C_D1274 VSS a_1769_14735# 0.01fF
C_D1275 VSS a_1586_18231# 0.01fF
C_D1276 VSS a_6664_26159# 0.01fF
C_D1277 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D1278 VSS a_30663_50087# 0.01fF
C_D1279 VSS a_1781_9308# 0.01fF
C_D128 VSS a_10883_3303# 0.01fF
C_D1280 VSS a_21739_29415# 0.01fF
C_D1281 VSS a_41731_49525# 0.01fF
C_D1282 VSS a_24867_53135# 0.01fF
C_D1283 VSS a_4383_7093# 0.01fF
C_D1284 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D1285 VSS a_5363_70543# 0.01fF
C_D1286 VSS a_2046_30184# 0.01fF
C_D1287 VSS a_15667_27239# 0.01fF
C_D1288 VSS a_2791_57703# 0.01fF
C_D1289 VSS a_4991_69831# 0.01fF
C_D129 VSS a_12116_40871# 0.01fF
C_D1290 VSS _1154_.A 0.01fF
C_D1291 VSS a_40837_46261# 0.01fF
C_D1292 VSS nmat.rowon_n[7] 0.01fF
C_D1293 VSS a_8583_29199# 0.01fF
C_D1294 VSS a_21739_29415# 0.01fF
C_D1295 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D1296 VSS a_9963_13967# 0.01fF
C_D1297 VSS a_2648_29397# 0.01fF
C_D1298 VSS a_1899_35051# 0.01fF
C_D1299 VSS a_30663_50087# 0.01fF
C_D13 VSS a_4128_64391# 0.01fF
C_D130 VSS a_5351_19913# 0.01fF
C_D1300 VSS a_38851_28327# 0.01fF
C_D1301 VSS a_2419_53351# 0.01fF
C_D1302 VSS a_17842_27497# 0.01fF
C_D1303 VSS a_2879_57487# 0.01fF
C_D1304 VSS a_4128_64391# 0.01fF
C_D1305 VSS a_41731_49525# 0.01fF
C_D1306 VSS a_12447_16143# 0.01fF
C_D1307 VSS _1154_.A 0.01fF
C_D1308 VSS a_40837_46261# 0.01fF
C_D1309 VSS a_3746_58487# 0.01fF
C_D131 VSS _1154_.A 0.01fF
C_D1310 VSS a_1591_31599# 0.01fF
C_D1311 VSS pmat.en_bit_n[2] 0.01fF
C_D1312 VSS a_41731_49525# 0.01fF
C_D1313 VSS _1187_.A2 0.01fF
C_D1314 VSS a_11067_27239# 0.01fF
C_D1315 VSS a_5363_33551# 0.01fF
C_D1316 VSS a_10239_14183# 0.01fF
C_D1317 VSS a_1858_25615# 0.01fF
C_D1318 VSS a_9963_13967# 0.01fF
C_D1319 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D132 VSS a_12447_16143# 0.01fF
C_D1320 VSS a_4075_31591# 0.01fF
C_D1321 VSS a_24407_31375# 0.01fF
C_D1322 VSS a_6559_33767# 0.01fF
C_D1323 VSS a_5363_33551# 0.01fF
C_D1324 VSS a_1781_9308# 0.01fF
C_D1325 VSS clk_ena 0.01fF
C_D1326 VSS a_1899_35051# 0.01fF
C_D1327 VSS a_9135_60967# 0.01fF
C_D1328 VSS a_10515_15055# 0.01fF
C_D1329 VSS a_17842_27497# 0.01fF
C_D133 VSS pmat.rowon_n[7] 0.01fF
C_D1330 VSS config_1_in[6] 0.01fF
C_D1331 VSS a_17139_30503# 0.01fF
C_D1332 VSS a_11067_64015# 0.01fF
C_D1333 VSS a_1674_57711# 0.01fF
C_D1334 VSS a_17139_30503# 0.01fF
C_D1335 VSS a_38851_28327# 0.01fF
C_D1336 VSS pmat.rowon_n[3] 0.01fF
C_D1337 VSS a_6467_29415# 0.01fF
C_D1338 VSS pmat.row_n[0] 0.01fF
C_D1339 VSS a_3746_58487# 0.01fF
C_D134 VSS a_2791_57703# 0.01fF
C_D1340 VSS a_40837_46261# 0.01fF
C_D1341 VSS a_24591_28327# 0.01fF
C_D1342 VSS a_8583_29199# 0.01fF
C_D1343 VSS a_2419_53351# 0.01fF
C_D1344 VSS a_2835_13077# 0.01fF
C_D1345 VSS a_15667_27239# 0.01fF
C_D1346 VSS a_2419_69455# 0.01fF
C_D1347 VSS a_6283_31591# 0.01fF
C_D1348 VSS a_26891_28327# 0.01fF
C_D1349 VSS a_30663_50087# 0.01fF
C_D135 VSS a_1586_63927# 0.01fF
C_D1350 VSS a_12116_40871# 0.01fF
C_D1351 VSS cgen.dlycontrol2_in[0] 0.01fF
C_D1352 VSS a_2791_57703# 0.01fF
C_D1353 VSS _1179_.X 0.01fF
C_D1354 VSS a_5651_66975# 0.01fF
C_D1355 VSS a_13641_23439# 0.01fF
C_D1356 VSS a_32687_46607# 0.01fF
C_D1357 VSS a_1923_31743# 0.01fF
C_D1358 VSS _1519_.A 0.01fF
C_D1359 VSS nmat.sw 0.01fF
C_D136 VSS a_5351_19913# 0.01fF
C_D1360 VSS a_13091_28327# 0.01fF
C_D1361 VSS config_1_in[4] 0.01fF
C_D1362 VSS a_4075_50087# 0.01fF
C_D1363 VSS a_13641_23439# 0.01fF
C_D1364 VSS _1154_.A 0.01fF
C_D1365 VSS pmat.rowon_n[7] 0.01fF
C_D1366 VSS a_7109_29423# 0.01fF
C_D1367 VSS pmat.row_n[9] 0.01fF
C_D1368 VSS a_2791_57703# 0.01fF
C_D1369 VSS a_2419_69455# 0.01fF
C_D137 VSS nmat.rowon_n[7] 0.01fF
C_D138 VSS a_2419_53351# 0.01fF
C_D139 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D14 VSS a_30663_50087# 0.01fF
C_D140 VSS pmat.row_n[12] 0.01fF
C_D141 VSS a_12447_16143# 0.01fF
C_D142 VSS config_2_in[2] 0.01fF
C_D143 VSS _1192_.B1 0.01fF
C_D144 VSS a_38851_28327# 0.01fF
C_D145 VSS a_33423_47695# 0.01fF
C_D146 VSS a_8443_20719# 0.01fF
C_D147 VSS a_1923_61759# 0.01fF
C_D148 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D149 VSS inp_analog 0.01fF
C_D15 VSS a_4351_55527# 0.01fF
C_D150 VSS a_5351_19913# 0.01fF
C_D151 VSS _1187_.A2 0.01fF
C_D152 VSS a_1923_61759# 0.01fF
C_D153 VSS a_5081_53135# 0.01fF
C_D154 VSS a_9963_13967# 0.01fF
C_D155 VSS a_2419_69455# 0.01fF
C_D156 VSS a_2046_30184# 0.01fF
C_D157 VSS a_1923_61759# 0.01fF
C_D158 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D159 VSS a_7415_29397# 0.01fF
C_D16 VSS _1184_.A2 0.01fF
C_D160 VSS a_1957_43567# 0.01fF
C_D161 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D162 VSS _1192_.B1 0.01fF
C_D163 VSS a_30111_47911# 0.01fF
C_D164 VSS ANTENNA__1190__A2.DIODE 0.01fF
C_D165 VSS a_10055_31591# 0.01fF
C_D166 VSS _1183_.A2 0.01fF
C_D167 VSS _1194_.A2 0.01fF
C_D168 VSS a_13459_28111# 0.01fF
C_D169 VSS a_11948_49783# 0.01fF
C_D17 VSS _1154_.X 0.01fF
C_D170 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D171 VSS a_5363_33551# 0.01fF
C_D172 VSS a_10515_61839# 0.01fF
C_D173 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D174 VSS _1154_.A 0.01fF
C_D175 VSS a_25879_31591# 0.01fF
C_D176 VSS a_6927_30503# 0.01fF
C_D177 VSS a_9135_60967# 0.01fF
C_D178 VSS a_10515_61839# 0.01fF
C_D179 VSS a_21371_50087# 0.01fF
C_D18 VSS a_1769_13103# 0.01fF
C_D180 VSS a_1586_50247# 0.01fF
C_D181 VSS a_2215_47375# 0.01fF
C_D182 VSS _1179_.X 0.01fF
C_D183 VSS cgen.dlycontrol4_in[4] 0.01fF
C_D184 VSS cgen.dlycontrol4_in[0] 0.01fF
C_D185 VSS a_1739_47893# 0.01fF
C_D186 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D187 VSS a_1923_61759# 0.01fF
C_D188 VSS a_11067_30287# 0.01fF
C_D189 VSS config_1_in[15] 0.01fF
C_D19 VSS a_11435_58791# 0.01fF
C_D190 VSS a_8583_29199# 0.01fF
C_D191 VSS a_41731_49525# 0.01fF
C_D192 VSS a_7717_14735# 0.01fF
C_D193 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D194 VSS a_2149_45717# 0.01fF
C_D195 VSS a_11948_49783# 0.01fF
C_D196 VSS a_4351_55527# 0.01fF
C_D197 VSS _1183_.A2 0.01fF
C_D198 VSS a_35244_32411# 0.01fF
C_D199 VSS a_1769_47919# 0.01fF
C_D2 VSS a_10781_42364# 0.01fF
C_D20 VSS a_2419_53351# 0.01fF
C_D200 VSS a_16311_28327# 0.01fF
C_D201 VSS _1192_.A2 0.01fF
C_D202 VSS a_9963_13967# 0.01fF
C_D203 VSS cgen.enable_dlycontrol_in 0.01fF
C_D204 VSS nmat.en_bit_n[0] 0.01fF
C_D205 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D206 VSS a_12263_50959# 0.01fF
C_D207 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D208 VSS a_10515_13967# 0.01fF
C_D209 VSS a_2407_49289# 0.01fF
C_D21 VSS a_29937_31055# 0.01fF
C_D210 VSS a_24867_53135# 0.01fF
C_D211 VSS a_2835_13077# 0.01fF
C_D212 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D213 VSS a_31675_47695# 0.01fF
C_D214 VSS pmat.sw 0.01fF
C_D215 VSS nmat.sw 0.01fF
C_D216 VSS a_6451_67655# 0.01fF
C_D217 VSS _1196_.B1 0.01fF
C_D218 VSS a_6283_31591# 0.01fF
C_D219 VSS _1194_.B1 0.01fF
C_D22 VSS config_2_in[8] 0.01fF
C_D220 VSS ANTENNA__1190__A2.DIODE 0.01fF
C_D221 VSS cgen.enable_dlycontrol_in 0.01fF
C_D222 VSS _1196_.B1 0.01fF
C_D223 VSS a_10515_61839# 0.01fF
C_D224 VSS _1183_.A2 0.01fF
C_D225 VSS a_28915_50959# 0.01fF
C_D226 VSS a_37820_30485# 0.01fF
C_D227 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D228 VSS a_4985_51433# 0.01fF
C_D229 VSS a_11067_49871# 0.01fF
C_D23 VSS a_2007_25597# 0.01fF
C_D230 VSS _1194_.A2 0.01fF
C_D231 VSS a_33423_47695# 0.01fF
C_D232 VSS a_2407_49289# 0.01fF
C_D233 VSS pmat.row_n[2] 0.01fF
C_D234 VSS _1154_.X 0.01fF
C_D235 VSS a_38851_28327# 0.01fF
C_D236 VSS a_2215_47375# 0.01fF
C_D237 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D238 VSS pmat.sw 0.01fF
C_D239 VSS a_3339_59879# 0.01fF
C_D24 VSS a_3339_70759# 0.01fF
C_D240 VSS a_4075_68583# 0.01fF
C_D241 VSS a_2419_53351# 0.01fF
C_D242 VSS a_11041_39860# 0.01fF
C_D243 VSS pmat.rowoff_n[12] 0.01fF
C_D244 VSS clk_vcm 0.01fF
C_D245 VSS a_21279_48999# 0.01fF
C_D246 VSS _1194_.A2 0.01fF
C_D247 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D248 VSS a_4075_50087# 0.01fF
C_D249 VSS a_41731_49525# 0.01fF
C_D25 VSS a_6283_31591# 0.01fF
C_D250 VSS a_24591_28327# 0.01fF
C_D251 VSS a_13641_23439# 0.01fF
C_D252 VSS a_11067_27239# 0.01fF
C_D253 VSS _1183_.A2 0.01fF
C_D254 VSS a_14379_6567# 0.01fF
C_D255 VSS a_30663_50087# 0.01fF
C_D256 VSS pmat.row_n[3] 0.01fF
C_D257 VSS nmat.sw 0.01fF
C_D258 VSS a_35312_31599# 0.01fF
C_D259 VSS a_18563_27791# 0.01fF
C_D26 VSS _1192_.A2 0.01fF
C_D260 VSS a_3746_58487# 0.01fF
C_D261 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D262 VSS a_1781_9308# 0.01fF
C_D263 VSS a_2007_25597# 0.01fF
C_D264 VSS a_11435_58791# 0.01fF
C_D265 VSS a_5081_53135# 0.01fF
C_D266 VSS pmat.row_n[14] 0.01fF
C_D267 VSS a_5363_70543# 0.01fF
C_D268 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D269 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D27 VSS a_13275_48783# 0.01fF
C_D270 VSS clk_ena 0.01fF
C_D271 VSS a_29937_31055# 0.01fF
C_D272 VSS a_3339_59879# 0.01fF
C_D273 VSS a_12309_38659# 0.01fF
C_D274 VSS a_11149_36924# 0.01fF
C_D275 VSS a_13091_18535# 0.01fF
C_D276 VSS a_8583_29199# 0.01fF
C_D277 VSS a_16311_28327# 0.01fF
C_D278 VSS _1194_.B1 0.01fF
C_D279 VSS config_1_in[2] 0.01fF
C_D28 VSS a_3339_59879# 0.01fF
C_D280 VSS a_26891_28327# 0.01fF
C_D281 VSS a_4075_50087# 0.01fF
C_D282 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D283 VSS a_4075_50087# 0.01fF
C_D284 VSS pmat.en_bit_n[2] 0.01fF
C_D285 VSS a_25879_31591# 0.01fF
C_D286 VSS a_2263_43719# 0.01fF
C_D287 VSS a_17139_30503# 0.01fF
C_D288 VSS nmat.rowon_n[7] 0.01fF
C_D289 VSS pmat.row_n[15] 0.01fF
C_D29 VSS a_7109_29423# 0.01fF
C_D290 VSS a_6467_29415# 0.01fF
C_D291 VSS a_6451_67655# 0.01fF
C_D292 VSS a_6467_29415# 0.01fF
C_D293 VSS a_30571_50959# 0.01fF
C_D294 VSS a_2411_43301# 0.01fF
C_D295 VSS a_25879_31591# 0.01fF
C_D296 VSS a_1586_63927# 0.01fF
C_D297 VSS a_10873_39605# 0.01fF
C_D298 VSS config_2_in[6] 0.01fF
C_D299 VSS a_1923_31743# 0.01fF
C_D3 VSS a_14287_69455# 0.01fF
C_D30 VSS clk_ena 0.01fF
C_D300 VSS a_4259_73807# 0.01fF
C_D301 VSS a_12447_16143# 0.01fF
C_D302 VSS a_17139_30503# 0.01fF
C_D303 VSS pmat.rowon_n[3] 0.01fF
C_D304 VSS a_1586_50247# 0.01fF
C_D305 VSS a_33423_47695# 0.01fF
C_D306 VSS _1196_.B1 0.01fF
C_D307 VSS a_12263_50959# 0.01fF
C_D308 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D309 VSS a_6559_33767# 0.01fF
C_D31 VSS a_10515_15055# 0.01fF
C_D310 VSS a_25879_31591# 0.01fF
C_D311 VSS a_2046_30184# 0.01fF
C_D312 VSS _1224_.X 0.01fF
C_D313 VSS a_6007_33767# 0.01fF
C_D314 VSS a_10515_61839# 0.01fF
C_D315 VSS a_4383_7093# 0.01fF
C_D316 VSS a_1781_9308# 0.01fF
C_D317 VSS a_3339_70759# 0.01fF
C_D318 VSS a_21371_50087# 0.01fF
C_D319 VSS config_2_in[7] 0.01fF
C_D32 VSS _1183_.A2 0.01fF
C_D320 VSS a_2879_57487# 0.01fF
C_D321 VSS pmat.row_n[5] 0.01fF
C_D322 VSS a_10781_42869# 0.01fF
C_D323 VSS a_30571_50959# 0.01fF
C_D324 VSS _1183_.A2 0.01fF
C_D325 VSS nmat.col_n[13] 0.01fF
C_D326 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D327 VSS _1179_.X 0.01fF
C_D328 VSS _1192_.B1 0.01fF
C_D329 VSS a_5363_33551# 0.01fF
C_D33 VSS cgen.dlycontrol4_in[4] 0.01fF
C_D330 VSS a_1586_18231# 0.01fF
C_D331 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D332 VSS _1184_.A2 0.01fF
C_D333 VSS a_4075_31591# 0.01fF
C_D334 VSS a_9135_60967# 0.01fF
C_D335 VSS a_17139_30503# 0.01fF
C_D336 VSS a_1586_18231# 0.01fF
C_D337 VSS a_13275_48783# 0.01fF
C_D338 VSS a_2419_53351# 0.01fF
C_D339 VSS a_13091_28327# 0.01fF
C_D34 VSS a_10239_14183# 0.01fF
C_D340 VSS a_7109_29423# 0.01fF
C_D341 VSS _1184_.A2 0.01fF
C_D342 VSS a_18243_28327# 0.01fF
C_D343 VSS a_1957_43567# 0.01fF
C_D344 VSS a_10441_21263# 0.01fF
C_D345 VSS a_6559_33767# 0.01fF
C_D346 VSS a_11067_64015# 0.01fF
C_D347 VSS a_6787_47607# 0.01fF
C_D348 VSS comp_latch 0.01fF
C_D349 VSS a_26891_28327# 0.01fF
C_D35 VSS a_1586_18231# 0.01fF
C_D350 VSS a_7415_29397# 0.01fF
C_D351 VSS a_41731_49525# 0.01fF
C_D352 VSS a_35244_32411# 0.01fF
C_D353 VSS a_11435_58791# 0.01fF
C_D354 VSS a_10515_13967# 0.01fF
C_D355 VSS a_3339_70759# 0.01fF
C_D356 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D357 VSS a_10239_14183# 0.01fF
C_D358 VSS comp_latch 0.01fF
C_D359 VSS pmat.rowon_n[0] 0.01fF
C_D36 VSS ANTENNA__1183__B1.DIODE 0.01fF
C_D360 VSS _1154_.A 0.01fF
C_D361 VSS a_11067_30287# 0.01fF
C_D362 VSS a_35244_32411# 0.01fF
C_D363 VSS a_1957_43567# 0.01fF
C_D364 VSS a_10873_38517# 0.01fF
C_D365 VSS pmat.rowon_n[7] 0.01fF
C_D366 VSS a_30111_47911# 0.01fF
C_D367 VSS a_2046_30184# 0.01fF
C_D368 VSS a_6467_29415# 0.01fF
C_D369 VSS cgen.dlycontrol4_in[1] 0.01fF
C_D37 VSS nmat.col[19] 0.01fF
C_D370 VSS a_2021_26677# 0.01fF
C_D371 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D372 VSS a_10883_3303# 0.01fF
C_D373 VSS a_12447_16143# 0.01fF
C_D374 VSS nmat.en_bit_n[1] 0.01fF
C_D375 VSS a_9963_13967# 0.01fF
C_D376 VSS nmat.sw 0.01fF
C_D377 VSS a_24747_29967# 0.01fF
C_D378 VSS a_24591_28327# 0.01fF
C_D379 VSS a_4991_69831# 0.01fF
C_D38 VSS a_15667_27239# 0.01fF
C_D380 VSS ANTENNA_fanout52_A.DIODE 0.01fF
C_D381 VSS a_10515_15055# 0.01fF
C_D382 VSS a_2149_45717# 0.01fF
C_D383 VSS a_25695_28111# 0.01fF
C_D384 VSS a_3339_70759# 0.01fF
C_D385 VSS a_28915_50959# 0.01fF
C_D386 VSS a_24867_53135# 0.01fF
C_D387 VSS a_9785_28879# 0.01fF
C_D388 VSS a_8491_47911# 0.01fF
C_D389 VSS a_40837_46261# 0.01fF
C_D39 VSS a_2263_43719# 0.01fF
C_D390 VSS a_14887_46377# 0.01fF
C_D391 VSS a_2791_57703# 0.01fF
C_D392 VSS a_7717_14735# 0.01fF
C_D393 VSS a_13091_28327# 0.01fF
C_D394 VSS a_4075_50087# 0.01fF
C_D395 VSS a_25695_28111# 0.01fF
C_D396 VSS clk_ena 0.01fF
C_D397 VSS pmat.row_n[13] 0.01fF
C_D398 VSS a_1674_57711# 0.01fF
C_D399 VSS a_10239_14183# 0.01fF
C_D4 VSS nmat.col_n[24] 0.01fF
C_D40 VSS a_1769_14735# 0.01fF
C_D400 VSS a_6787_47607# 0.01fF
C_D401 VSS nmat.col_n[1] 0.01fF
C_D402 VSS pmat.row_n[1] 0.01fF
C_D403 VSS _1187_.A2 0.01fF
C_D404 VSS a_18243_28327# 0.01fF
C_D405 VSS a_10239_14183# 0.01fF
C_D406 VSS a_4383_7093# 0.01fF
C_D407 VSS a_10515_61839# 0.01fF
C_D408 VSS _1154_.X 0.01fF
C_D409 VSS nmat.rowon_n[12] 0.01fF
C_D41 VSS nmat.col_n[31] 0.01fF
C_D410 VSS a_2263_43719# 0.01fF
C_D411 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D412 VSS nmat.col[12] 0.01fF
C_D413 VSS a_2215_47375# 0.01fF
C_D414 VSS a_8583_29199# 0.01fF
C_D415 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D416 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D417 VSS pmat.row_n[6] 0.01fF
C_D418 VSS a_2407_49289# 0.01fF
C_D419 VSS a_10239_14183# 0.01fF
C_D42 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D420 VSS _1192_.A2 0.01fF
C_D421 VSS a_24867_53135# 0.01fF
C_D422 VSS pmat.row_n[15] 0.01fF
C_D423 VSS config_2_in[15] 0.01fF
C_D424 VSS a_38851_28327# 0.01fF
C_D425 VSS start_conversion_in 0.01fF
C_D426 VSS cgen.dlycontrol4_in[0] 0.01fF
C_D427 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D428 VSS a_3746_58487# 0.01fF
C_D429 VSS a_2215_47375# 0.01fF
C_D43 VSS a_7939_31591# 0.01fF
C_D430 VSS a_1674_57711# 0.01fF
C_D431 VSS a_28915_50959# 0.01fF
C_D432 VSS a_1739_47893# 0.01fF
C_D433 VSS a_21371_50087# 0.01fF
C_D434 VSS a_10515_15055# 0.01fF
C_D435 VSS pmat.row_n[1] 0.01fF
C_D436 VSS a_9963_13967# 0.01fF
C_D437 VSS cgen.enable_dlycontrol_in 0.01fF
C_D438 VSS a_11067_27239# 0.01fF
C_D439 VSS a_13459_28111# 0.01fF
C_D44 VSS a_35244_32411# 0.01fF
C_D440 VSS a_10781_42869# 0.01fF
C_D441 VSS config_2_in[1] 0.01fF
C_D442 VSS a_13091_52047# 0.01fF
C_D443 VSS a_8491_47911# 0.01fF
C_D444 VSS a_2046_30184# 0.01fF
C_D445 VSS _1154_.X 0.01fF
C_D446 VSS a_4075_50087# 0.01fF
C_D447 VSS a_1769_13103# 0.01fF
C_D448 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D449 VSS pmat.row_n[7] 0.01fF
C_D45 VSS a_6283_31591# 0.01fF
C_D450 VSS a_38851_28327# 0.01fF
C_D451 VSS a_1858_25615# 0.01fF
C_D452 VSS a_3339_70759# 0.01fF
C_D453 VSS nmat.sw 0.01fF
C_D454 VSS a_13643_29415# 0.01fF
C_D455 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D456 VSS a_11067_27239# 0.01fF
C_D457 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D458 VSS cgen.dlycontrol1_in[1] 0.01fF
C_D459 VSS _1154_.X 0.01fF
C_D46 VSS a_10515_13967# 0.01fF
C_D460 VSS a_10055_31591# 0.01fF
C_D461 VSS a_37820_30485# 0.01fF
C_D462 VSS a_10873_36341# 0.01fF
C_D463 VSS a_1586_18231# 0.01fF
C_D464 VSS a_10239_14183# 0.01fF
C_D465 VSS a_8491_47911# 0.01fF
C_D466 VSS a_9411_2215# 0.01fF
C_D467 VSS a_40837_46261# 0.01fF
C_D468 VSS a_21371_50087# 0.01fF
C_D469 VSS a_30111_47911# 0.01fF
C_D47 VSS a_7415_29397# 0.01fF
C_D470 VSS a_9411_2215# 0.01fF
C_D471 VSS a_29937_31055# 0.01fF
C_D472 VSS a_4075_31591# 0.01fF
C_D473 VSS a_38851_28327# 0.01fF
C_D474 VSS a_9411_2215# 0.01fF
C_D475 VSS a_33423_47695# 0.01fF
C_D476 VSS a_4259_31375# 0.01fF
C_D477 VSS pmat.rowon_n[7] 0.01fF
C_D478 VSS a_25695_28111# 0.01fF
C_D479 VSS a_10515_15055# 0.01fF
C_D48 VSS pmat.row_n[13] 0.01fF
C_D480 VSS pmat.rowon_n[11] 0.01fF
C_D481 VSS a_37820_30485# 0.01fF
C_D482 VSS a_12069_38517# 0.01fF
C_D483 VSS a_22199_30287# 0.01fF
C_D484 VSS nmat.col[3] 0.01fF
C_D485 VSS clk_ena 0.01fF
C_D486 VSS a_11435_58791# 0.01fF
C_D487 VSS a_11067_49871# 0.01fF
C_D488 VSS pmat.rowon_n[0] 0.01fF
C_D489 VSS a_1957_43567# 0.01fF
C_D49 VSS a_4128_64391# 0.01fF
C_D490 VSS a_11067_30287# 0.01fF
C_D491 VSS pmat.row_n[0] 0.01fF
C_D492 VSS a_4383_7093# 0.01fF
C_D493 VSS a_2835_13077# 0.01fF
C_D494 VSS a_7109_29423# 0.01fF
C_D495 VSS a_4075_68583# 0.01fF
C_D496 VSS a_13091_52047# 0.01fF
C_D497 VSS a_37820_30485# 0.01fF
C_D498 VSS a_30663_50087# 0.01fF
C_D499 VSS a_11067_64015# 0.01fF
C_D5 VSS _1179_.X 0.01fF
C_D50 VSS a_21739_29415# 0.01fF
C_D500 VSS a_11067_64015# 0.01fF
C_D501 VSS a_13275_48783# 0.01fF
C_D502 VSS a_35244_32411# 0.01fF
C_D503 VSS pmat.row_n[12] 0.01fF
C_D504 VSS a_7109_29423# 0.01fF
C_D505 VSS a_2263_43719# 0.01fF
C_D506 VSS a_11067_16359# 0.01fF
C_D507 VSS a_2046_30184# 0.01fF
C_D508 VSS config_1_in[5] 0.01fF
C_D509 VSS a_1769_47919# 0.01fF
C_D51 VSS a_2648_29397# 0.01fF
C_D510 VSS ANTENNA__1195__A1.DIODE 0.01fF
C_D511 VSS a_4259_73807# 0.01fF
C_D512 VSS cgen.dlycontrol1_in[4] 0.01fF
C_D513 VSS a_40837_46261# 0.01fF
C_D514 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D515 VSS a_1586_63927# 0.01fF
C_D516 VSS a_4075_31591# 0.01fF
C_D517 VSS a_2411_43301# 0.01fF
C_D518 VSS a_4985_51433# 0.01fF
C_D519 VSS a_1586_50247# 0.01fF
C_D52 VSS a_16311_28327# 0.01fF
C_D520 VSS a_1586_50247# 0.01fF
C_D521 VSS _1194_.B1 0.01fF
C_D522 VSS a_26891_28327# 0.01fF
C_D523 VSS a_2149_45717# 0.01fF
C_D524 VSS a_3615_71631# 0.01fF
C_D525 VSS nmat.col[28] 0.01fF
C_D526 VSS a_11067_27239# 0.01fF
C_D527 VSS a_10515_61839# 0.01fF
C_D528 VSS a_9135_60967# 0.01fF
C_D529 VSS a_6787_47607# 0.01fF
C_D53 VSS a_10883_3303# 0.01fF
C_D530 VSS a_5651_66975# 0.01fF
C_D531 VSS a_4075_50087# 0.01fF
C_D532 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D533 VSS a_4991_69831# 0.01fF
C_D534 VSS config_2_in[12] 0.01fF
C_D535 VSS cgen.dlycontrol2_in[1] 0.01fF
C_D536 VSS a_4383_7093# 0.01fF
C_D537 VSS a_10441_21263# 0.01fF
C_D538 VSS a_11149_40188# 0.01fF
C_D539 VSS a_5351_19913# 0.01fF
C_D54 VSS a_10515_13967# 0.01fF
C_D540 VSS a_2791_57703# 0.01fF
C_D541 VSS a_10055_31591# 0.01fF
C_D542 VSS a_2879_57487# 0.01fF
C_D543 VSS a_1781_9308# 0.01fF
C_D544 VSS a_15667_27239# 0.01fF
C_D545 VSS nmat.col_n[26] 0.01fF
C_D546 VSS pmat.row_n[7] 0.01fF
C_D547 VSS _1187_.A2 0.01fF
C_D548 VSS pmat.row_n[3] 0.01fF
C_D549 VSS a_24407_31375# 0.01fF
C_D55 VSS a_3615_71631# 0.01fF
C_D550 VSS a_24867_53135# 0.01fF
C_D551 VSS pmat.row_n[10] 0.01fF
C_D552 VSS a_10883_3303# 0.01fF
C_D553 VSS cgen.dlycontrol1_in[3] 0.01fF
C_D554 VSS a_4075_50087# 0.01fF
C_D555 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D556 VSS a_10055_31591# 0.01fF
C_D557 VSS a_5363_70543# 0.01fF
C_D558 VSS a_33423_47695# 0.01fF
C_D559 VSS a_4128_64391# 0.01fF
C_D56 VSS a_11067_16359# 0.01fF
C_D560 VSS a_1899_35051# 0.01fF
C_D561 VSS a_4259_31375# 0.01fF
C_D562 VSS a_9963_13967# 0.01fF
C_D563 VSS a_23395_53135# 0.01fF
C_D564 VSS a_10781_42364# 0.01fF
C_D565 VSS cgen.dlycontrol1_in[0] 0.01fF
C_D566 VSS nmat.col_n[7] 0.01fF
C_D567 VSS a_5363_70543# 0.01fF
C_D568 VSS a_4985_51433# 0.01fF
C_D569 VSS a_10515_15055# 0.01fF
C_D57 VSS a_2407_49289# 0.01fF
C_D570 VSS pmat.row_n[9] 0.01fF
C_D571 VSS a_18243_28327# 0.01fF
C_D572 VSS a_15667_27239# 0.01fF
C_D573 VSS config_1_in[10] 0.01fF
C_D574 VSS _1192_.A2 0.01fF
C_D575 VSS a_5363_33551# 0.01fF
C_D576 VSS a_4128_64391# 0.01fF
C_D577 VSS nmat.en_bit_n[1] 0.01fF
C_D578 VSS a_3615_71631# 0.01fF
C_D579 VSS a_5651_66975# 0.01fF
C_D58 VSS a_1899_35051# 0.01fF
C_D580 VSS a_35244_32411# 0.01fF
C_D581 VSS a_13459_28111# 0.01fF
C_D582 VSS a_1586_63927# 0.01fF
C_D583 VSS nmat.sample_n 0.01fF
C_D584 VSS a_32687_46607# 0.01fF
C_D585 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D586 VSS a_26891_28327# 0.01fF
C_D587 VSS config_1_in[14] 0.01fF
C_D588 VSS nmat.rowon_n[7] 0.01fF
C_D589 VSS a_11067_27239# 0.01fF
C_D59 VSS a_5081_53135# 0.01fF
C_D590 VSS a_6927_30503# 0.01fF
C_D591 VSS a_10055_31591# 0.01fF
C_D592 VSS a_9963_13967# 0.01fF
C_D593 VSS _1224_.X 0.01fF
C_D594 VSS _1183_.A2 0.01fF
C_D595 VSS a_1858_25615# 0.01fF
C_D596 VSS a_6467_29415# 0.01fF
C_D597 VSS a_25695_28111# 0.01fF
C_D598 VSS a_10239_14183# 0.01fF
C_D599 VSS nmat.col[30] 0.01fF
C_D6 VSS a_10515_15055# 0.01fF
C_D60 VSS a_11435_58791# 0.01fF
C_D600 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D601 VSS a_1923_61759# 0.01fF
C_D602 VSS _1224_.X 0.01fF
C_D603 VSS a_18563_27791# 0.01fF
C_D604 VSS a_6664_26159# 0.01fF
C_D605 VSS a_12447_16143# 0.01fF
C_D606 VSS a_32405_32463# 0.01fF
C_D607 VSS nmat.col[21] 0.01fF
C_D608 VSS a_10055_31591# 0.01fF
C_D609 VSS a_2835_13077# 0.01fF
C_D61 VSS _1194_.A2 0.01fF
C_D610 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D611 VSS a_6787_47607# 0.01fF
C_D612 VSS nmat.sw 0.01fF
C_D613 VSS a_15667_27239# 0.01fF
C_D614 VSS a_9411_2215# 0.01fF
C_D615 VSS a_13091_28327# 0.01fF
C_D616 VSS a_1923_31743# 0.01fF
C_D617 VSS a_2046_30184# 0.01fF
C_D618 VSS a_11317_36924# 0.01fF
C_D619 VSS a_18243_28327# 0.01fF
C_D62 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D620 VSS a_13091_28327# 0.01fF
C_D621 VSS nmat.sw 0.01fF
C_D622 VSS a_2149_45717# 0.01fF
C_D623 VSS a_4991_69831# 0.01fF
C_D624 VSS a_2007_25597# 0.01fF
C_D625 VSS a_1899_35051# 0.01fF
C_D626 VSS a_2648_29397# 0.01fF
C_D627 VSS a_13091_28327# 0.01fF
C_D628 VSS a_8491_47911# 0.01fF
C_D629 VSS a_2149_45717# 0.01fF
C_D63 VSS a_2879_57487# 0.01fF
C_D630 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D631 VSS a_2021_26677# 0.01fF
C_D632 VSS ANTENNA__1190__A2.DIODE 0.01fF
C_D633 VSS a_9411_2215# 0.01fF
C_D634 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D635 VSS a_1957_43567# 0.01fF
C_D636 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D637 VSS a_12069_38517# 0.01fF
C_D638 VSS a_6451_67655# 0.01fF
C_D639 VSS a_6787_47607# 0.01fF
C_D64 VSS a_2648_29397# 0.01fF
C_D640 VSS cgen.dlycontrol2_in[2] 0.01fF
C_D641 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D642 VSS a_13459_28111# 0.01fF
C_D643 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D644 VSS a_2407_49289# 0.01fF
C_D645 VSS a_11067_16359# 0.01fF
C_D646 VSS a_4719_30287# 0.01fF
C_D647 VSS a_13091_52047# 0.01fF
C_D648 VSS a_4985_51433# 0.01fF
C_D649 VSS nmat.col_n[28] 0.01fF
C_D65 VSS a_15667_27239# 0.01fF
C_D650 VSS clk_dig 0.01fF
C_D651 VSS a_3615_71631# 0.01fF
C_D652 VSS nmat.col[7] 0.01fF
C_D653 VSS pmat.rowon_n[7] 0.01fF
C_D654 VSS _1194_.B1 0.01fF
C_D655 VSS a_11067_30287# 0.01fF
C_D656 VSS a_3339_59879# 0.01fF
C_D657 VSS a_35244_32411# 0.01fF
C_D658 VSS a_28915_50959# 0.01fF
C_D659 VSS clk_ena 0.01fF
C_D66 VSS a_13091_52047# 0.01fF
C_D660 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D661 VSS a_5081_53135# 0.01fF
C_D662 VSS a_2149_45717# 0.01fF
C_D663 VSS ndecision_finish 0.01fF
C_D664 VSS a_11435_58791# 0.01fF
C_D665 VSS _1187_.A2 0.01fF
C_D666 VSS a_2791_57703# 0.01fF
C_D667 VSS a_30571_50959# 0.01fF
C_D668 VSS _1154_.X 0.01fF
C_D669 VSS a_1586_63927# 0.01fF
C_D67 VSS a_2149_45717# 0.01fF
C_D670 VSS a_11067_64015# 0.01fF
C_D671 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D672 VSS config_2_in[9] 0.01fF
C_D673 VSS a_7415_29397# 0.01fF
C_D674 VSS a_30663_50087# 0.01fF
C_D675 VSS _1192_.A2 0.01fF
C_D676 VSS a_10873_40693# 0.01fF
C_D677 VSS a_26891_28327# 0.01fF
C_D678 VSS a_11041_39860# 0.01fF
C_D679 VSS a_10515_61839# 0.01fF
C_D68 VSS a_2411_43301# 0.01fF
C_D680 VSS a_24407_31375# 0.01fF
C_D681 VSS a_3339_70759# 0.01fF
C_D682 VSS a_1781_9308# 0.01fF
C_D683 VSS nmat.rowon_n[7] 0.01fF
C_D684 VSS a_30571_50959# 0.01fF
C_D685 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D686 VSS a_2835_13077# 0.01fF
C_D687 VSS nmat.rowon_n[7] 0.01fF
C_D688 VSS _1194_.A2 0.01fF
C_D689 VSS a_3746_58487# 0.01fF
C_D69 VSS a_2648_29397# 0.01fF
C_D690 VSS config_1_in[13] 0.01fF
C_D691 VSS a_22199_30287# 0.01fF
C_D692 VSS a_24407_31375# 0.01fF
C_D693 VSS ANTENNA_fanout52_A.DIODE 0.01fF
C_D694 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D695 VSS a_10515_15055# 0.01fF
C_D696 VSS a_1858_25615# 0.01fF
C_D697 VSS pmat.rowoff_n[12] 0.01fF
C_D698 VSS a_12263_50959# 0.01fF
C_D699 VSS a_2648_29397# 0.01fF
C_D7 VSS a_26891_28327# 0.01fF
C_D70 VSS a_2411_43301# 0.01fF
C_D700 VSS a_24407_31375# 0.01fF
C_D701 VSS _1192_.B1 0.01fF
C_D702 VSS a_2149_45717# 0.01fF
C_D703 VSS a_10055_31591# 0.01fF
C_D704 VSS a_11067_64015# 0.01fF
C_D705 VSS pmat.rowon_n[7] 0.01fF
C_D706 VSS _1179_.X 0.01fF
C_D707 VSS a_38851_28327# 0.01fF
C_D708 VSS _1194_.A2 0.01fF
C_D709 VSS a_10515_13967# 0.01fF
C_D71 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D710 VSS ANTENNA__1183__B1.DIODE 0.01fF
C_D711 VSS a_32687_46607# 0.01fF
C_D712 VSS _1184_.A2 0.01fF
C_D713 VSS a_1781_9308# 0.01fF
C_D714 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D715 VSS a_1586_63927# 0.01fF
C_D716 VSS a_5651_66975# 0.01fF
C_D717 VSS a_4259_73807# 0.01fF
C_D718 VSS a_4259_31375# 0.01fF
C_D719 VSS cgen.dlycontrol4_in[2] 0.01fF
C_D72 VSS a_4351_55527# 0.01fF
C_D720 VSS a_18243_28327# 0.01fF
C_D721 VSS a_2648_29397# 0.01fF
C_D722 VSS ANTENNA__1190__A2.DIODE 0.01fF
C_D723 VSS a_24591_28327# 0.01fF
C_D724 VSS a_2419_69455# 0.01fF
C_D725 VSS a_2419_53351# 0.01fF
C_D726 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D727 VSS a_4991_69831# 0.01fF
C_D728 VSS cgen.dlycontrol3_in[2] 0.01fF
C_D729 VSS a_7717_14735# 0.01fF
C_D73 VSS a_9411_2215# 0.01fF
C_D730 VSS a_2046_30184# 0.01fF
C_D731 VSS a_1586_50247# 0.01fF
C_D732 VSS a_12079_9615# 0.01fF
C_D733 VSS a_1586_63927# 0.01fF
C_D734 VSS a_11067_64015# 0.01fF
C_D735 VSS a_1858_25615# 0.01fF
C_D736 VSS a_11113_39747# 0.01fF
C_D737 VSS a_3615_71631# 0.01fF
C_D738 VSS a_1957_43567# 0.01fF
C_D739 VSS a_4719_30287# 0.01fF
C_D74 VSS a_1781_9308# 0.01fF
C_D740 VSS a_11067_30287# 0.01fF
C_D741 VSS a_31675_47695# 0.01fF
C_D742 VSS a_2407_49289# 0.01fF
C_D743 VSS a_6283_31591# 0.01fF
C_D744 VSS ANTENNA_fanout52_A.DIODE 0.01fF
C_D745 VSS a_25695_28111# 0.01fF
C_D746 VSS a_5179_31591# 0.01fF
C_D747 VSS _1184_.A2 0.01fF
C_D748 VSS a_10883_3303# 0.01fF
C_D749 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D75 VSS a_6451_67655# 0.01fF
C_D750 VSS a_5363_70543# 0.01fF
C_D751 VSS a_11067_16359# 0.01fF
C_D752 VSS _1194_.B1 0.01fF
C_D753 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D754 VSS a_1769_47919# 0.01fF
C_D755 VSS a_30111_47911# 0.01fF
C_D756 VSS a_17139_30503# 0.01fF
C_D757 VSS a_14887_46377# 0.01fF
C_D758 VSS a_6927_30503# 0.01fF
C_D759 VSS a_18597_31599# 0.01fF
C_D76 VSS a_30663_50087# 0.01fF
C_D760 VSS a_1769_47919# 0.01fF
C_D761 VSS clk_ena 0.01fF
C_D762 VSS a_3615_71631# 0.01fF
C_D763 VSS a_5351_19913# 0.01fF
C_D764 VSS a_11067_30287# 0.01fF
C_D765 VSS a_5363_33551# 0.01fF
C_D766 VSS a_13641_23439# 0.01fF
C_D767 VSS a_2879_57487# 0.01fF
C_D768 VSS a_11435_58791# 0.01fF
C_D769 VSS a_3339_70759# 0.01fF
C_D77 VSS a_1899_35051# 0.01fF
C_D770 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D771 VSS a_10873_36341# 0.01fF
C_D772 VSS a_6451_67655# 0.01fF
C_D773 VSS a_12263_50959# 0.01fF
C_D774 VSS a_10883_3303# 0.01fF
C_D775 VSS comp_latch 0.01fF
C_D776 VSS _1192_.A2 0.01fF
C_D777 VSS a_5363_33551# 0.01fF
C_D778 VSS a_1586_18231# 0.01fF
C_D779 VSS a_41731_49525# 0.01fF
C_D78 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D780 VSS ANTENNA__1183__B1.DIODE 0.01fF
C_D781 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D782 VSS a_3339_59879# 0.01fF
C_D783 VSS a_1586_63927# 0.01fF
C_D784 VSS a_1923_31743# 0.01fF
C_D785 VSS a_11149_36924# 0.01fF
C_D786 VSS a_24867_53135# 0.01fF
C_D787 VSS a_1923_31743# 0.01fF
C_D788 VSS a_1923_31743# 0.01fF
C_D789 VSS nmat.col_n[18] 0.01fF
C_D79 VSS a_11297_36091# 0.01fF
C_D790 VSS a_9411_2215# 0.01fF
C_D791 VSS a_16311_28327# 0.01fF
C_D792 VSS a_4351_55527# 0.01fF
C_D793 VSS a_28915_50959# 0.01fF
C_D794 VSS a_4128_64391# 0.01fF
C_D795 VSS a_11067_64015# 0.01fF
C_D796 VSS a_1923_31743# 0.01fF
C_D797 VSS a_21371_50087# 0.01fF
C_D798 VSS a_1586_18231# 0.01fF
C_D799 VSS ANTENNA__1197__A.DIODE 0.01fF
C_D8 VSS a_10147_29415# 0.01fF
C_D80 VSS a_6787_47607# 0.01fF
C_D800 VSS clk_dig 0.01fF
C_D801 VSS a_5179_31591# 0.01fF
C_D802 VSS a_18563_27791# 0.01fF
C_D803 VSS a_26891_28327# 0.01fF
C_D804 VSS a_2419_53351# 0.01fF
C_D805 VSS a_21739_29415# 0.01fF
C_D806 VSS a_6559_33767# 0.01fF
C_D807 VSS a_41731_49525# 0.01fF
C_D808 VSS pmat.rowon_n[7] 0.01fF
C_D809 VSS a_29937_31055# 0.01fF
C_D81 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D810 VSS pmat.rowon_n[11] 0.01fF
C_D811 VSS a_10515_15055# 0.01fF
C_D812 VSS config_1_in[0] 0.01fF
C_D813 VSS a_28915_50959# 0.01fF
C_D814 VSS a_19541_28879# 0.01fF
C_D815 VSS a_12447_16143# 0.01fF
C_D816 VSS a_4259_31375# 0.01fF
C_D817 VSS nmat.rowon_n[7] 0.01fF
C_D818 VSS _1154_.X 0.01fF
C_D819 VSS a_11113_40835# 0.01fF
C_D82 VSS a_11435_58791# 0.01fF
C_D820 VSS a_23395_53135# 0.01fF
C_D821 VSS a_2648_29397# 0.01fF
C_D822 VSS nmat.en_bit_n[0] 0.01fF
C_D823 VSS a_1739_47893# 0.01fF
C_D824 VSS a_5363_33551# 0.01fF
C_D825 VSS a_3339_59879# 0.01fF
C_D826 VSS a_21739_29415# 0.01fF
C_D827 VSS a_10515_61839# 0.01fF
C_D828 VSS a_1923_61759# 0.01fF
C_D829 VSS a_5081_53135# 0.01fF
C_D83 VSS a_14887_46377# 0.01fF
C_D830 VSS a_5363_70543# 0.01fF
C_D831 VSS a_24747_29967# 0.01fF
C_D832 VSS a_10055_31591# 0.01fF
C_D833 VSS a_11067_16359# 0.01fF
C_D834 VSS a_13091_52047# 0.01fF
C_D835 VSS a_7415_29397# 0.01fF
C_D836 VSS a_5351_19913# 0.01fF
C_D837 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D838 VSS ANTENNA__1197__B.DIODE 0.01fF
C_D839 VSS a_2879_57487# 0.01fF
C_D84 VSS a_18243_28327# 0.01fF
C_D840 VSS a_1674_57711# 0.01fF
C_D841 VSS rst_n 0.01fF
C_D842 VSS a_33423_47695# 0.01fF
C_D843 VSS _1179_.X 0.01fF
C_D844 VSS ANTENNA__1395__B1.DIODE 0.01fF
C_D845 VSS a_10883_3303# 0.01fF
C_D846 VSS a_4351_55527# 0.01fF
C_D847 VSS cgen.dlycontrol4_in[1] 0.01fF
C_D848 VSS a_22199_30287# 0.01fF
C_D849 VSS cgen.enable_dlycontrol_in 0.01fF
C_D85 VSS _1179_.X 0.01fF
C_D850 VSS ANTENNA__1190__A1.DIODE 0.01fF
C_D851 VSS pmat.sample_n 0.01fF
C_D852 VSS a_12263_50959# 0.01fF
C_D853 VSS _1192_.B1 0.01fF
C_D854 VSS a_10873_39605# 0.01fF
C_D855 VSS a_21739_29415# 0.01fF
C_D856 VSS a_11067_30287# 0.01fF
C_D857 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D858 VSS a_21739_29415# 0.01fF
C_D859 VSS a_40837_46261# 0.01fF
C_D86 VSS pmat.rowoff_n[15] 0.01fF
C_D860 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D861 VSS a_18243_28327# 0.01fF
C_D862 VSS a_7717_14735# 0.01fF
C_D863 VSS pmat.rowoff_n[4] 0.01fF
C_D864 VSS a_26891_28327# 0.01fF
C_D865 VSS a_24747_29967# 0.01fF
C_D866 VSS pmat.en_bit_n[0] 0.01fF
C_D867 VSS ANTENNA__1196__A2.DIODE 0.01fF
C_D868 VSS a_22199_30287# 0.01fF
C_D869 VSS config_2_in[11] 0.01fF
C_D87 VSS a_9963_28111# 0.01fF
C_D870 VSS a_1586_63927# 0.01fF
C_D871 VSS a_1923_31743# 0.01fF
C_D872 VSS a_11435_58791# 0.01fF
C_D873 VSS a_2215_47375# 0.01fF
C_D874 VSS a_30111_47911# 0.01fF
C_D875 VSS ANTENNA__1184__B1.DIODE 0.01fF
C_D876 VSS a_1674_57711# 0.01fF
C_D877 VSS config_2_in[10] 0.01fF
C_D878 VSS a_11067_16359# 0.01fF
C_D879 VSS a_2835_13077# 0.01fF
C_D88 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D880 VSS a_2879_57487# 0.01fF
C_D881 VSS a_1957_43567# 0.01fF
C_D882 VSS pmat.rowoff_n[7] 0.01fF
C_D883 VSS a_12447_16143# 0.01fF
C_D884 VSS a_1586_63927# 0.01fF
C_D885 VSS a_7415_29397# 0.01fF
C_D886 VSS a_12263_50959# 0.01fF
C_D887 VSS a_6927_30503# 0.01fF
C_D888 VSS a_6927_30503# 0.01fF
C_D889 VSS a_6467_29415# 0.01fF
C_D89 VSS a_1769_14735# 0.01fF
C_D890 VSS config_2_in[4] 0.01fF
C_D891 VSS a_32405_32463# 0.01fF
C_D892 VSS a_22199_30287# 0.01fF
C_D893 VSS a_16311_28327# 0.01fF
C_D894 VSS pmat.rowon_n[8] 0.01fF
C_D895 VSS a_10883_3303# 0.01fF
C_D896 VSS cgen.enable_dlycontrol_in 0.01fF
C_D897 VSS a_5081_53135# 0.01fF
C_D898 VSS config_2_in[14] 0.01fF
C_D899 VSS config_1_in[7] 0.01fF
C_D9 VSS ANTENNA__1395__A1.DIODE 0.01fF
C_D90 VSS a_23395_53135# 0.01fF
C_D900 VSS a_10147_29415# 0.01fF
C_D901 VSS a_11497_40719# 0.01fF
C_D902 VSS a_2879_57487# 0.01fF
C_D903 VSS pmat.sw 0.01fF
C_D904 VSS a_6283_31591# 0.01fF
C_D905 VSS pmat.row_n[11] 0.01fF
C_D906 VSS _1154_.A 0.01fF
C_D907 VSS a_16311_28327# 0.01fF
C_D908 VSS a_11711_50959# 0.01fF
C_D909 VSS _1196_.B1 0.01fF
C_D91 VSS a_11711_50959# 0.01fF
C_D910 VSS a_40837_46261# 0.01fF
C_D911 VSS ANTENNA__1187__B1.DIODE 0.01fF
C_D912 VSS _1192_.B1 0.01fF
C_D913 VSS a_24867_53135# 0.01fF
C_D914 VSS a_3339_70759# 0.01fF
C_D915 VSS a_6787_47607# 0.01fF
C_D916 VSS a_10873_40693# 0.01fF
C_D917 VSS pmat.rowoff_n[4] 0.01fF
C_D918 VSS a_9411_2215# 0.01fF
C_D919 VSS a_1858_25615# 0.01fF
C_D92 VSS a_7717_14735# 0.01fF
C_D920 VSS a_30571_50959# 0.01fF
C_D921 VSS a_18563_27791# 0.01fF
C_D922 VSS a_13459_28111# 0.01fF
C_D923 VSS a_13091_28327# 0.01fF
C_D924 VSS a_11067_27239# 0.01fF
C_D925 VSS a_41731_49525# 0.01fF
C_D926 VSS a_12263_50959# 0.01fF
C_D927 VSS a_1586_18231# 0.01fF
C_D928 VSS a_24591_28327# 0.01fF
C_D929 VSS a_4351_55527# 0.01fF
C_D93 VSS a_13091_52047# 0.01fF
C_D930 VSS _1187_.A2 0.01fF
C_D931 VSS nmat.col[1] 0.01fF
C_D932 VSS a_10515_15055# 0.01fF
C_D933 VSS a_24867_53135# 0.01fF
C_D934 VSS a_28915_50959# 0.01fF
C_D935 VSS a_41731_49525# 0.01fF
C_D936 VSS a_4075_31591# 0.01fF
C_D937 VSS comp_latch 0.01fF
C_D938 VSS _1187_.A2 0.01fF
C_D939 VSS a_22199_30287# 0.01fF
C_D94 VSS a_2149_45717# 0.01fF
C_D940 VSS pmat.row_n[11] 0.01fF
C_D941 VSS cgen.dlycontrol3_in[4] 0.01fF
C_D942 VSS a_33423_47695# 0.01fF
C_D943 VSS a_6664_26159# 0.01fF
C_D944 VSS a_24591_28327# 0.01fF
C_D945 VSS _1224_.X 0.01fF
C_D946 VSS a_35244_32411# 0.01fF
C_D947 VSS a_1591_31599# 0.01fF
C_D948 VSS cgen.dlycontrol3_in[3] 0.01fF
C_D949 VSS a_9135_60967# 0.01fF
C_D95 VSS a_23395_53135# 0.01fF
C_D950 VSS a_2419_69455# 0.01fF
C_D951 VSS _1192_.A2 0.01fF
C_D952 VSS a_17842_27497# 0.01fF
C_D953 VSS nmat.col_n[21] 0.01fF
C_D954 VSS a_18243_28327# 0.01fF
C_D955 VSS a_24867_53135# 0.01fF
C_D956 VSS _1154_.X 0.01fF
C_D957 VSS a_13459_28111# 0.01fF
C_D958 VSS a_1674_57711# 0.01fF
C_D959 VSS a_2407_49289# 0.01fF
C_D96 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D960 VSS cgen.dlycontrol4_in[3] 0.01fF
C_D961 VSS a_30571_50959# 0.01fF
C_D962 VSS a_9135_60967# 0.01fF
C_D963 VSS ANTENNA__1395__A2.DIODE 0.01fF
C_D964 VSS a_5351_19913# 0.01fF
C_D965 VSS a_26891_28327# 0.01fF
C_D966 VSS nmat.col_n[29] 0.01fF
C_D967 VSS a_24591_28327# 0.01fF
C_D968 VSS a_1781_9308# 0.01fF
C_D969 VSS a_25879_31591# 0.01fF
C_D97 VSS a_31675_47695# 0.01fF
C_D970 VSS nmat.sw 0.01fF
C_D971 VSS a_5351_19913# 0.01fF
C_D972 VSS a_17842_27497# 0.01fF
C_D973 VSS a_4351_55527# 0.01fF
C_D974 VSS a_2835_13077# 0.01fF
C_D975 VSS ANTENNA__1190__B1.DIODE 0.01fF
C_D976 VSS config_1_in[3] 0.01fF
C_D977 VSS config_2_in[0] 0.01fF
C_D978 VSS a_2419_53351# 0.01fF
C_D979 VSS a_24867_53135# 0.01fF
C_D98 VSS a_35244_32411# 0.01fF
C_D980 VSS a_35244_32411# 0.01fF
C_D981 VSS nmat.col[10] 0.01fF
C_D982 VSS a_7717_14735# 0.01fF
C_D983 VSS a_4259_73807# 0.01fF
C_D984 VSS config_1_in[12] 0.01fF
C_D985 VSS inn_analog 0.01fF
C_D986 VSS a_7415_29397# 0.01fF
C_D987 VSS nmat.col_n[3] 0.01fF
C_D988 VSS a_12447_16143# 0.01fF
C_D989 VSS clk_ena 0.01fF
C_D99 VSS a_3339_70759# 0.01fF
C_D990 VSS a_38851_28327# 0.01fF
C_D991 VSS a_6007_33767# 0.01fF
C_D992 VSS config_2_in[3] 0.01fF
C_D993 VSS nmat.col[13] 0.01fF
C_D994 VSS a_21279_48999# 0.01fF
C_D995 VSS a_2149_45717# 0.01fF
C_D996 VSS pmat.row_n[4] 0.01fF
C_D997 VSS a_1781_9308# 0.01fF
C_D998 VSS a_28915_50959# 0.01fF
C_D999 VSS a_7415_29397# 0.01fF
R0 dummypin[11] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 adc_top_84.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R10 VDD adc_top_92.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R11 dummypin[6] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R12 VSS a_14833_72049# sky130_fd_pr__res_generic_po w=480000u l=45000u
R13 VDD adc_top_81.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R14 VDD adc_top_86.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R15 VDD adc_top_93.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R16 VSS dummypin[15] sky130_fd_pr__res_generic_po w=480000u l=45000u
R17 VDD adc_top_87.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R18 VDD pmat.rowoff_n[0] sky130_fd_pr__res_generic_po w=480000u l=45000u
R19 dummypin[7] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R2 pmat.en_C0_n VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R20 VSS dummypin[13] sky130_fd_pr__res_generic_po w=480000u l=45000u
R21 VSS dummypin[1] sky130_fd_pr__res_generic_po w=480000u l=45000u
R22 VSS dummypin[8] sky130_fd_pr__res_generic_po w=480000u l=45000u
R23 VDD adc_top_88.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R24 adc_top_96.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R25 VSS a_20583_28529# sky130_fd_pr__res_generic_po w=480000u l=45000u
R26 dummypin[9] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R27 adc_top_94.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R28 adc_top_82.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R29 adc_top_89.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R3 VSS a_14833_23089# sky130_fd_pr__res_generic_po w=480000u l=45000u
R30 VDD a_20583_53080# sky130_fd_pr__res_generic_po w=480000u l=45000u
R31 nmat.rowoff_n[0] VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R32 dummypin[10] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R33 VDD adc_top_90.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R34 VSS dummypin[14] sky130_fd_pr__res_generic_po w=480000u l=45000u
R35 dummypin[4] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R36 pmat.rowon_n[15] VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R37 VDD adc_top_91.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R38 a_14833_56053# VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R39 adc_top_95.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R4 VSS a_14833_8945# sky130_fd_pr__res_generic_po w=480000u l=45000u
R40 VDD adc_top_85.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
R41 VSS dummypin[3] sky130_fd_pr__res_generic_po w=480000u l=45000u
R42 nmat.en_C0_n VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R43 VSS dummypin[2] sky130_fd_pr__res_generic_po w=480000u l=45000u
R5 dummypin[0] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R6 dummypin[5] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
R7 adc_top_83.HI VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R8 nmat.rowon_n[15] VDD sky130_fd_pr__res_generic_po w=480000u l=45000u
R9 dummypin[12] VSS sky130_fd_pr__res_generic_po w=480000u l=45000u
X0 a_1644_72917# a_1591_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=4.7895e+15p ps=3.06454e+10u w=420000u l=150000u
X1 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u M=530
X10 a_34134_20942# a_18162_20536# a_34226_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X100 vcm a_18162_23548# a_48282_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1000 a_44570_9858# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10000 VDD a_6664_26159# a_8206_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10001 a_22178_57134# a_18546_57176# a_22086_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10002 VDD pmat.rowoff_n[12] a_49194_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10003 a_40250_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10004 a_19074_72194# a_18162_72234# a_19166_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10005 a_23182_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10006 a_49194_61150# a_18162_61190# a_49286_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10007 VSS pmat.row_n[6] a_22482_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10008 a_6244_34863# a_6127_35076# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10009 VDD a_33957_48437# a_36209_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=2
X1001 a_19605_32149# a_19439_32149# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10010 a_43662_9460# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10011 VSS a_45187_38129# a_45133_38155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10012 VDD pmat.rowoff_n[4] a_39154_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10013 VSS a_16837_35515# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X10014 a_16311_28327# a_45915_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=8
X10015 a_41475_31751# a_26479_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10016 VDD a_21239_47349# a_18547_51565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10017 vcm a_18162_68218# a_26194_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10018 a_11113_40835# a_36617_42043# a_37680_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10019 VDD pmat.rowon_n[15] a_26102_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1002 a_47186_15922# pmat.row_n[7] a_47678_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10020 VSS a_14773_37218# a_13837_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X10021 VSS a_5271_23447# a_4516_21531# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X10022 a_26479_32117# a_27443_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X10023 vcm a_18162_18528# a_44266_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10024 VDD a_41297_27221# nmat.col[22] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10025 a_5123_52423# a_4075_50087# a_5185_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10026 a_26194_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10027 VSS a_2835_13077# a_12949_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10028 a_45064_44807# a_33423_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10029 VSS pmat.row_n[10] a_47582_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1003 a_49590_7850# VDD a_49194_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10030 a_2250_65693# a_2163_65469# a_1846_65579# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X10031 a_12323_12937# a_11877_12565# a_12227_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10032 a_51598_64202# pmat.rowon_n[8] a_51202_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10033 VDD nmat.rowon_n[14] a_29114_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10034 a_24094_21946# a_18162_21540# a_24186_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10035 VDD pmat.rowon_n[7] a_34134_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10036 a_21174_18528# a_18546_18526# a_21082_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10037 a_41558_56170# pmat.rowon_n[0] a_41162_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10038 VDD nmat.rowon_n[5] a_38150_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10039 a_34226_17524# a_18546_17522# a_34134_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1004 VSS pmat.row_n[13] a_47582_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10040 VSS pmat.row_n[9] a_20474_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10041 a_49286_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10042 a_14747_63401# a_11067_64015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10043 VSS a_19965_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X10044 a_28116_39655# a_26957_39867# a_28079_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10045 a_13160_31433# a_12245_31061# a_12813_31029# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X10046 a_31518_21906# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10047 VDD a_8397_71285# a_8287_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10048 a_39154_69182# a_18162_69222# a_39246_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10049 a_11054_71311# a_11019_71543# a_10751_71543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 a_5602_11471# a_1717_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X10050 a_34134_57134# pmat.row_n[1] a_34626_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10051 vcm a_18162_14512# a_22178_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10052 a_33413_31599# a_32771_31599# a_33331_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10053 a_43262_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10054 a_45574_55166# VSS a_45178_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10055 vcm a_18162_56170# a_21174_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10056 VDD a_17739_50871# a_17163_50857# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X10057 VDD a_2672_20553# a_2847_20479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10058 VSS a_2683_22089# a_7847_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10059 a_2621_48981# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1006 a_42258_24552# a_18546_24550# a_42166_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10060 a_28506_65206# pmat.rowon_n[9] a_28110_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10061 a_27106_9898# a_18162_9492# a_27198_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10062 vcm a_18162_13508# a_35230_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10063 VSS a_6283_31591# a_7571_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10064 a_21478_13874# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10065 VDD a_15899_47939# a_15711_47899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10066 VDD pmat.rowon_n[12] a_46182_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10067 VDD a_8727_70197# a_7658_71543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10068 a_34530_12870# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10069 a_46578_63198# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1007 a_82863_64213# _1154_.A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u M=3
X10070 a_11159_28585# a_5991_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X10071 a_24638_49159# a_21215_48071# a_24941_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10072 VSS a_18823_50247# a_19439_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X10073 VDD a_8928_56457# a_9103_56383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10074 a_35068_46805# a_35540_46983# a_35306_46831# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X10075 a_6292_69831# a_8539_76181# a_8497_76457# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10076 a_2325_34017# a_2107_33775# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X10077 a_38557_47381# a_38391_47381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X10078 VDD a_28901_48437# a_30189_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X10079 a_6559_6031# a_6337_6825# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1008 a_1899_35051# a_2419_69455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X10080 vcm a_18162_72234# a_47278_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10081 a_1761_7119# a_1591_7119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10082 a_16381_42919# a_16689_43132# a_16355_43123# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10083 a_2672_8585# a_1591_8213# a_2325_8181# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10084 a_51294_70186# a_18546_70228# a_51202_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10085 a_20063_30877# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X10086 a_44174_22950# pmat.row_n[14] a_44666_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10087 nmat.rowoff_n[11] a_9963_13967# a_14287_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10088 a_47278_60146# a_18546_60188# a_47186_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10089 a_47678_64524# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1009 a_41254_66170# a_18546_66212# a_41162_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10090 VSS pmat.row_n[7] a_23486_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10091 a_20474_60186# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10092 a_20474_19898# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10093 VDD pmat.rowon_n[6] a_51202_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10094 a_51202_64162# a_18162_64202# a_51294_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10095 a_12629_68047# a_12789_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10096 a_37542_23914# pmat.rowoff_n[15] a_37146_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10097 VDD a_12407_28853# a_12437_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10098 a_4503_70455# a_3615_71631# a_4677_70561# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10099 a_33526_18894# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X101 a_31614_21508# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1010 a_51694_13476# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10100 a_13252_18377# a_12171_18005# a_12905_17973# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10101 a_10053_15521# a_9835_15279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10102 a_24186_72194# a_18546_72236# a_24094_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10103 a_37638_56492# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10104 a_48682_7452# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10105 a_44570_7850# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10106 a_24937_41479# a_24197_42405# a_25319_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10107 VSS a_10378_7637# a_10319_7663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10108 a_21574_22512# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10109 a_46723_30485# a_43776_30287# a_47005_30511# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X1011 a_5692_55509# a_5784_52423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X10110 a_42258_22544# a_18546_22542# a_42166_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10111 VSS pmat.row_n[1] a_37542_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10112 a_48190_60146# pmat.row_n[4] a_48682_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10113 VSS a_1717_13647# a_8732_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10114 VDD a_35290_44527# a_36111_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10115 VSS a_33719_34191# a_33825_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10116 a_7109_29423# a_4339_27804# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=0p ps=0u w=650000u l=150000u M=4
X10117 a_19405_28853# a_7415_29397# a_19439_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10118 a_9195_60039# a_1769_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10119 a_25098_72194# VDD a_25590_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1012 a_37238_56130# a_18546_56172# a_37146_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10120 a_36538_70226# pmat.rowon_n[14] a_36142_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10121 a_25590_21508# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10122 a_25190_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10123 a_46274_21540# a_18546_21538# a_46182_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10124 a_22086_14918# a_18162_14512# a_22178_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10125 a_35534_9858# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10126 VDD a_7385_51701# a_7275_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10127 VSS nmat.rowon_n[7] nmat.rowoff_n[8] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X10128 a_17440_38567# a_16377_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10129 a_50594_65206# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1013 a_34626_23516# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10130 a_8363_73865# a_7847_73493# a_8268_73853# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X10131 a_31479_31375# a_31339_31787# a_30527_31573# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10132 a_7521_47081# a_6830_44655# a_7165_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.3328e+12p pd=1.271e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X10133 VSS a_8749_57141# a_8507_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X10134 a_19166_23548# a_18546_23546# a_19074_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10135 a_6970_67191# a_2407_49289# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10136 a_2621_48981# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10137 a_28602_12472# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10138 a_13160_31433# a_12079_31061# a_12813_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10139 a_40554_57174# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1014 a_20811_44535# a_19417_43990# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X10140 a_26102_13914# a_18162_13508# a_26194_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10141 VDD nmat.rowon_n[13] a_32126_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10142 a_23486_67214# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10143 a_46182_63158# pmat.row_n[7] a_46674_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10144 a_12461_29673# a_11603_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X10145 a_28573_48463# a_28629_48437# a_21215_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10146 VSS a_20503_48981# pmat.row_n[9] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X10147 a_15439_48071# a_15711_47899# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10148 a_30514_68218# pmat.rowon_n[12] a_30118_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10149 a_50690_61512# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1015 a_34226_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10150 a_9287_77055# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10151 a_44266_69182# a_18546_69224# a_44174_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10152 VSS a_11142_64783# a_11793_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10153 VSS a_2411_43301# a_2461_45565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10154 a_13804_65161# a_12889_64789# a_13457_64757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10155 VDD a_46817_43541# a_46582_46519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10156 a_3484_58229# a_3746_58487# a_3704_58575# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X10157 a_41654_19500# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10158 VDD a_17996_44007# a_17900_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10159 VSS a_25879_31591# a_31535_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1016 a_14005_22589# a_3305_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X10160 VDD a_31263_28309# a_31209_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X10161 a_45915_29941# a_46723_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X10162 a_10845_12559# a_10471_12791# a_10773_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X10163 a_22482_9858# nmat.rowon_n[14] a_22086_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10164 a_44647_36201# a_35244_32411# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X10165 vcm a_18162_61190# a_19166_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10166 a_19719_52521# a_11067_64015# a_19623_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10167 a_23700_36391# a_22541_36603# a_23663_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10168 a_18546_62196# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X10169 a_23582_63520# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1017 VDD pmat.rowon_n[2] a_41162_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10170 a_29391_36395# a_24833_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10171 a_33526_59182# pmat.rowon_n[3] a_33130_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10172 a_3876_58255# a_2957_58255# a_3621_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X10173 a_18162_16520# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X10174 a_27598_18496# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10175 a_5325_9269# a_4611_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10176 a_2867_43541# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10177 a_6737_77295# a_5547_77295# a_6628_77295# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X10178 VDD nmat.rowon_n[7] a_31122_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10179 a_48282_68178# a_18546_68220# a_48190_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1018 a_23663_36649# a_22541_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X10180 vcm a_18162_65206# a_45270_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10181 a_45178_69182# pmat.row_n[13] a_45670_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10182 a_35499_28023# a_26891_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X10183 a_12488_38543# a_12237_38772# a_12267_38870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X10184 VSS a_12038_55687# a_11835_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10185 a_4909_54447# a_4843_54826# a_4837_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10186 a_32126_67174# a_18162_67214# a_32218_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10187 a_25681_46831# a_25090_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10188 VDD a_11202_55687# a_11877_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10189 VSS pmat.en_bit_n[1] a_34530_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1019 a_19623_52521# a_19584_52423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10190 VSS a_13837_36893# a_13529_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10191 a_11521_64239# a_10049_60663# a_11533_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X10192 VDD a_10878_58487# a_10190_60663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10193 a_31122_7890# a_18162_7484# a_31214_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10194 a_22178_65166# a_18546_65208# a_22086_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10195 a_38841_31055# a_31339_31787# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10196 a_22578_69544# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10197 a_46274_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10198 a_45923_28111# ANTENNA__1195__A1.DIODE nmat.col_n[25] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X10199 a_5725_76207# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X102 a_31214_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1020 VSS a_4075_50087# a_5123_52423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X10200 VDD a_12437_28879# a_16966_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X10201 a_19399_48437# a_19283_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10202 a_22086_59142# a_18162_59182# a_22178_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10203 a_4308_24135# a_4339_27804# a_4450_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10204 a_42562_17890# nmat.rowon_n[6] a_42166_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10205 a_3429_76725# a_3211_77129# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X10206 a_13699_72777# a_13183_72405# a_13604_72765# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X10207 a_1828_25589# a_2007_25597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X10208 a_40158_55126# VDD a_40650_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10209 a_7565_15279# a_6375_15279# a_7456_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1021 VSS pmat.row_n[5] a_37542_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10210 a_49590_23914# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10211 VDD a_76962_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10212 a_39013_43655# a_39193_43131# a_40315_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10213 a_23090_65166# pmat.row_n[9] a_23582_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10214 result_out[13] a_1644_72917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X10215 a_44266_14512# a_18546_14510# a_44174_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10216 a_54136_39932# comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top comp.adc_comp_circuit_0.adc_comp_buffer_0.in VDD sky130_fd_pr__pfet_01v8 ad=1.32e+12p pd=9.32e+06u as=1.24e+12p ps=9.24e+06u w=2e+06u l=150000u M=2
X10217 a_43262_56130# a_18546_56172# a_43170_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10218 VSS a_10953_34951# a_12255_34473# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X10219 a_51598_72234# VDD a_51202_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1022 a_2012_23805# a_1895_23610# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X10220 a_26102_58138# a_18162_58178# a_26194_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10221 a_35012_39655# a_33949_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10222 a_10141_60431# a_10049_60663# a_10058_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10223 a_39550_15882# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10224 VSS nmat.sample_n a_18162_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X10225 VSS pmat.row_n[5] a_43566_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10226 a_27249_28995# a_22459_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10227 a_40554_10862# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10228 VSS a_11091_26311# a_10791_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10229 a_6741_42721# a_6523_42479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1023 a_41558_11866# nmat.rowon_n[12] a_41162_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10230 VDD a_39472_47753# a_39647_47679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10231 VDD comp.adc_comp_circuit_0.adc_comp_buffer_0.in a_53622_39932# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u M=2
X10232 a_26102_17930# pmat.row_n[9] a_26594_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10233 VSS pmat.row_n[15] a_26498_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10234 VDD pmat.rowon_n[15] a_34134_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10235 a_9459_5461# a_10747_6727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X10236 a_23486_20902# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10237 a_11979_22057# a_11892_21959# a_11897_21813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10238 a_30610_15484# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10239 a_30514_21906# nmat.rowon_n[2] a_30118_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1024 a_31879_34191# a_31702_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10240 a_30463_41271# a_30857_41245# a_30523_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X10241 VDD a_9279_71829# a_9183_72007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10242 VDD pmat.rowon_n[1] a_33130_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10243 a_48586_70226# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10244 a_36253_38567# a_36561_38780# a_36227_38771# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10245 VDD a_3325_43023# a_3983_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10246 VSS a_9963_13967# a_13446_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10247 a_19470_18894# nmat.rowon_n[5] a_19074_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10248 a_20474_13874# nmat.rowon_n[10] a_20078_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10249 vcm a_18162_8488# a_40250_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1025 a_30514_56170# pmat.rowon_n[0] a_30118_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10250 a_38546_62194# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10251 a_33526_12870# pmat.rowoff_n[4] a_33130_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10252 a_40158_72194# a_18162_72234# a_40250_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10253 a_45574_63198# pmat.rowon_n[7] a_45178_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10254 VSS pmat.row_n[4] a_42562_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10255 vcm a_18162_64202# a_21174_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10256 a_31122_11906# pmat.row_n[3] a_31614_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10257 VSS pmat.row_n[11] a_42562_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10258 a_21082_68178# pmat.row_n[12] a_21574_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10259 VSS a_17187_49783# a_17139_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X1026 VDD nmat.rowon_n[5] a_27106_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10260 vcm a_18162_21540# a_35230_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10261 VDD pmat.rowon_n[3] a_24094_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10262 a_26317_40726# a_25393_41317# a_26515_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10263 VSS a_19332_41959# a_19145_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10264 a_39646_24520# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10265 a_26194_8488# a_18546_8486# a_26102_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10266 VDD a_17054_28995# a_17306_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10267 VDD nmat.rowon_n[1] a_43170_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10268 vcm a_18162_58178# a_43262_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10269 a_27345_46831# a_26155_46831# a_27236_46831# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1027 a_24586_15484# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10270 VSS a_28245_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X10271 a_1644_71285# a_1591_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10272 VDD a_5320_57863# a_3770_57399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10273 a_47005_30511# a_43533_30761# a_46921_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10274 VDD cgen.dlycontrol3_in[0] a_10767_39087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10275 a_4535_38377# a_4533_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X10276 a_45546_49257# a_45370_48169# a_45238_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.25e+11p pd=2.65e+06u as=0p ps=0u w=1e+06u l=150000u
X10277 a_18203_48981# a_18359_49140# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10278 a_23663_38825# a_23700_38567# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X10279 a_24719_39605# a_24895_39605# a_24847_39631# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X1028 a_45270_65166# a_18546_65208# a_45178_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10280 VSS a_25061_43132# a_24753_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10281 VSS pmat.row_n[15] a_50594_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10282 VSS a_13688_47893# a_13632_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10283 a_49590_64202# pmat.rowon_n[8] a_49194_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10284 a_47678_72556# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10285 VDD nmat.rowon_n[2] a_47186_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10286 a_42955_31849# a_35244_32411# a_42307_31756# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10287 a_20353_49667# a_10515_13967# a_20257_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10288 VDD pmat.rowon_n[14] a_51202_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10289 vcm a_18162_69222# a_33222_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1029 a_9135_49257# a_4719_30287# a_9217_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X10290 a_44266_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10291 a_44444_32233# a_35312_31599# a_45164_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10292 VDD a_12993_66415# a_14443_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10293 a_47186_62154# a_18162_62194# a_47278_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10294 a_30118_19938# pmat.row_n[11] a_30610_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10295 a_3173_25045# a_2648_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10296 a_51294_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10297 a_39550_56170# pmat.rowon_n[0] a_39154_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10298 a_20170_13508# a_18546_13506# a_20078_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10299 a_46863_28585# a_38851_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X103 VSS a_46947_39215# _1187_.A2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=8
X1030 vcm a_18162_62194# a_42258_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10300 a_34226_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10301 VDD nmat.rowon_n[10] a_37146_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10302 a_2107_20553# a_1591_20181# a_2012_20541# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X10303 VSS a_13091_52047# a_18011_50729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10304 VSS a_25647_39783# a_11339_39319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10305 VDD a_12967_12863# a_12954_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10306 VDD a_14195_7351# a_14195_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X10307 a_33222_12504# a_18546_12502# a_33130_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10308 a_10681_12879# comp_latch VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10309 VSS a_3480_17143# a_2467_16341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1031 a_12723_53609# a_9581_56079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X10310 vcm a_18162_19532# a_42258_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10311 VSS a_27794_28879# a_28626_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.72e+11p ps=4.36e+06u w=650000u l=150000u
X10312 a_18176_41605# a_17113_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10313 a_33845_27765# a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10314 a_48282_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10315 a_24186_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10316 a_41558_18894# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10317 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top vcm.sky130_fd_sc_hd__buf_4_0.X vcm VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=500000u M=2
X10318 VDD a_40099_52245# pmat.col[20] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10319 a_2325_50337# a_2107_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1032 a_45670_69544# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10320 a_12651_29423# a_6830_22895# a_12461_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X10321 a_27605_28995# a_25315_28335# a_27532_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X10322 a_1769_47919# a_1769_13103# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X10323 a_22086_22950# a_18162_22544# a_22178_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10324 a_45270_71190# a_18546_71232# a_45178_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10325 VDD a_10239_77295# a_10383_75637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10326 a_35138_21946# a_18162_21540# a_35230_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10327 VDD pmat.rowon_n[7] a_45178_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10328 a_32218_18528# a_18546_18526# a_32126_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10329 a_7201_62313# a_1823_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 a_42166_66170# pmat.row_n[10] a_42658_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10330 VSS pmat.row_n[1] a_45574_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10331 VSS a_2163_31741# a_2124_31867# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10332 pmat.col_n[19] a_39757_50700# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10333 VDD a_21147_49525# pmat.row_n[13] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10334 VSS pmat.row_n[9] a_31518_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10335 VDD a_17154_43671# a_17159_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10336 VDD a_9405_66627# a_10167_64239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X10337 a_20179_51843# a_18547_51565# a_20083_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10338 VSS pmat.row_n[2] a_39550_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10339 a_4611_9839# a_4338_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1034 a_9983_32385# a_2046_30184# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10340 a_46182_71190# pmat.row_n[15] a_46674_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10341 a_41254_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10342 a_3473_77117# a_3429_76725# a_3307_77129# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10343 a_7313_74005# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10344 VDD a_6787_47607# a_12235_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10345 VDD pmat.rowon_n[6] a_49194_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10346 vcm a_18162_14512# a_33222_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10347 a_6741_42721# a_6523_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10348 vcm a_18162_56170# a_32218_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10349 a_31923_42367# cgen.dlycontrol4_in[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1035 VDD a_8051_46607# a_8453_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10350 a_11071_39631# a_10817_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10351 a_32522_13874# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10352 VDD ANTENNA__1195__A1.DIODE a_22377_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10353 a_33222_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10354 VDD a_35244_32411# a_47499_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10355 a_78448_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_0.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10356 a_23582_71552# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10357 a_44266_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10358 a_19566_61512# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10359 a_5462_58038# a_4351_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1036 a_35138_15922# a_18162_15516# a_35230_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10360 a_27198_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10361 a_13013_27023# a_9217_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10362 VDD a_6976_32375# a_5963_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10363 a_7900_54269# a_5211_57172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10364 a_44570_66210# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10365 a_42166_8894# pmat.row_n[0] a_42658_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10366 a_42166_23954# pmat.row_n[15] a_42658_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10367 VSS a_7999_31359# a_4259_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X10368 a_13279_68841# a_13173_68597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10369 a_42166_19938# a_18162_19532# a_42258_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1037 VDD a_2439_13889# a_2400_13763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10370 VDD a_18568_51959# a_18199_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10371 a_36538_8854# nmat.rowon_n[15] a_36142_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10372 a_6639_23413# pmat.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10373 a_13322_31055# a_12245_31061# a_13160_31433# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10374 a_48282_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10375 a_33239_46287# a_14887_46377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10376 a_45178_55126# a_18162_55166# a_45270_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10377 a_3879_42997# a_2021_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10378 a_35630_18496# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10379 a_35534_24918# nmat.en_bit_n[2] a_35138_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1038 VDD a_20848_41605# a_20752_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X10380 VSS pmat.row_n[7] a_34530_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10381 VDD a_37823_34191# nmat.sample_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X10382 a_24490_69222# pmat.rowon_n[13] a_24094_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10383 VSS pmat.row_n[10] a_21478_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10384 a_24490_8854# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10385 a_28602_8456# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10386 vcm a_18162_17524# a_31214_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10387 a_4073_37039# a_4031_37191# a_2467_35925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X10388 a_10949_43124# a_10979_42390# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10389 a_45178_14918# pmat.row_n[6] a_45670_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1039 a_45238_49007# a_44774_48695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X10390 a_48682_17492# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10391 a_48586_23914# pmat.rowoff_n[15] a_48190_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10392 a_46182_18934# a_18162_18528# a_46274_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10393 a_2847_18303# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10394 a_28110_24958# VDD a_28602_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10395 VSS pmat.row_n[0] a_34530_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10396 a_32618_22512# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10397 a_2203_18377# a_1757_18005# a_2107_18377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10398 a_22178_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10399 VDD a_9581_56079# a_12461_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X104 a_44382_41167# a_44774_40821# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=0p ps=0u w=650000u l=150000u M=4
X1040 a_14465_29575# a_12851_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10400 a_38546_15882# pmat.rowoff_n[7] a_38150_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10401 a_23479_43447# a_22357_43493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10402 VDD a_5323_71829# a_5271_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10403 nmat.col[30] _1154_.X a_84090_3087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X10404 VSS a_18823_50247# a_24270_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10405 a_18272_39429# a_17113_39141# a_18176_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10406 VSS pmat.row_n[9] a_25494_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10407 a_8725_10422# comp_latch a_8511_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X10408 a_1761_9839# a_1591_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10409 a_31203_28111# _1154_.X nmat.col_n[9] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X1041 a_8206_26703# a_2683_22089# a_8114_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X10410 VSS a_14113_43132# a_13805_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10411 a_22578_14480# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10412 VDD nmat.rowon_n[6] a_25098_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10413 vcm a_18162_66210# a_39246_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10414 a_49194_13914# pmat.row_n[5] a_49686_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10415 a_29163_29423# a_28626_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X10416 a_20078_15922# a_18162_15516# a_20170_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10417 a_23182_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10418 a_43262_64162# a_18546_64204# a_43170_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10419 vcm a_18162_61190# a_40250_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1042 a_25098_11906# pmat.row_n[3] a_25590_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10420 a_4298_69367# a_4075_68583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10421 a_43662_68540# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10422 VDD a_6741_42721# a_6631_42845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X10423 a_39646_58500# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10424 VDD a_13896_8585# a_14071_8511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10425 a_33130_14918# a_18162_14512# a_33222_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10426 a_1761_6031# a_1591_6031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10427 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10428 VSS pmat.row_n[3] a_39550_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10429 VSS a_24407_31375# a_31388_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1043 VSS config_2_in[2] a_1591_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10430 VDD a_12248_42583# a_12061_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10431 VSS pmat.row_n[0] a_28506_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10432 a_44665_45519# a_44573_45173# a_44447_45431# VSS sky130_fd_pr__nfet_01v8 ad=6.24e+11p pd=5.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10433 a_15048_40517# a_13985_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10434 a_30210_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10435 VDD nmat.rowon_n[7] a_29114_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10436 a_26594_13476# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10437 a_23090_10902# pmat.row_n[2] a_23582_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10438 VSS a_5687_71829# a_11990_73309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10439 VDD nmat.rowon_n[12] a_30118_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1044 VSS a_23807_41959# a_12116_39783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10440 vcm a_18162_60186# a_44266_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10441 a_28356_29199# a_16478_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10442 a_7445_29673# a_7415_29397# a_7027_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10443 VDD pmat.rowon_n[12] a_20078_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10444 a_44174_64162# pmat.row_n[8] a_44666_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10445 a_6611_57399# a_4025_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X10446 vcm a_18162_8488# a_49286_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10447 a_10499_67503# a_10226_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10448 VSS a_38711_37683# a_38651_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X10449 a_9669_28585# a_5351_19913# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1045 a_40127_28111# ANTENNA__1195__A1.DIODE nmat.col_n[20] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10450 nmat.rowon_n[14] a_19474_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10451 a_20811_35831# a_19689_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X10452 vcm a_18162_72234# a_21174_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10453 a_5253_18543# a_5087_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10454 VDD a_14287_69455# a_14839_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X10455 a_21174_60146# a_18546_60188# a_21082_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10456 vcm a_18162_71230# a_34226_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10457 VDD pmat.rowon_n[11] a_24094_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10458 a_21574_64524# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10459 a_38242_15516# a_18546_15514# a_38150_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1046 a_27603_34191# cgen.dlycontrol2_in[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10460 a_25821_34219# a_25755_34343# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10461 a_5278_19958# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10462 a_3052_29967# a_2217_29973# a_3080_30333# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10463 a_33775_29111# a_31339_31787# a_34009_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10464 VSS a_14149_39747# a_20251_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X10465 a_34626_63520# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10466 VSS a_2655_72373# a_1823_74557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10467 VDD a_45112_47607# a_45943_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X10468 a_4683_30511# a_4333_30511# a_4588_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X10469 a_38907_47753# a_38391_47381# a_38812_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X1047 VSS a_5087_19319# a_5087_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10470 VDD a_2983_48071# a_2971_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10471 a_35167_52521# a_34942_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10472 a_24490_22910# nmat.rowon_n[1] a_24094_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10473 a_10955_55687# a_11743_55329# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10474 a_1881_65327# a_1846_65579# a_1643_65301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10475 a_28506_58178# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10476 VSS a_12463_22351# a_13641_23439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X10477 a_13805_36391# a_14113_36604# a_13779_36595# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10478 a_6799_75637# a_6803_77269# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10479 a_22086_60146# pmat.row_n[4] a_22578_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1048 VDD pmat.rowon_n[13] a_22086_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10480 vcm a_18162_11500# a_39246_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10481 a_22620_32509# a_6007_33767# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X10482 a_30118_68178# a_18162_68218# a_30210_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10483 a_49590_72234# VDD a_49194_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10484 a_18546_59184# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X10485 a_36341_39141# a_35108_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X10486 VDD a_11979_47068# a_11910_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X10487 a_44266_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10488 pmat.rowon_n[13] a_14839_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10489 VSS a_4339_27804# a_9135_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1049 a_36234_17524# a_18546_17522# a_36142_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10490 a_10697_75218# a_14071_74879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10491 a_12247_20175# a_11995_20291# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10492 a_28765_36395# a_28431_34735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10493 VSS pmat.row_n[5] a_36538_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10494 a_20170_21540# a_18546_21538# a_20078_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10495 a_8693_11769# a_2021_11043# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10496 a_40554_18894# nmat.rowon_n[5] a_40158_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10497 VSS pmat.row_n[15] a_19470_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10498 a_33130_59142# a_18162_59182# a_33222_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10499 vcm a_18162_22544# a_29206_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X105 a_14371_66665# a_13718_68591# a_14289_66421# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1050 a_46182_65166# pmat.row_n[9] a_46674_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10500 a_5711_18909# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10501 VSS a_1586_50247# a_8583_47381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10502 a_33222_20536# a_18546_20534# a_33130_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10503 a_47582_24918# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10504 a_29206_10496# a_18546_10494# a_29114_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10505 vcm a_18162_69222# a_41254_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10506 a_51202_16926# pmat.row_n[8] a_51694_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10507 a_6242_70767# a_6200_70919# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10508 vcm a_18162_59182# a_37238_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10509 a_41254_57134# a_18546_57176# a_41162_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1051 a_1881_53181# a_1846_52947# a_1643_52789# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10510 a_37542_16886# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10511 a_18546_24550# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X10512 a_24719_38517# a_12513_39100# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10513 VSS pmat.row_n[6] a_41558_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10514 a_37638_9460# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10515 a_2931_40277# a_2419_69455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10516 VSS pmat.row_n[3] a_30514_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10517 a_24094_18934# pmat.row_n[10] a_24586_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10518 VSS VDD a_24490_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10519 VSS a_15839_49525# a_10515_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X1052 ANTENNA__1395__B1.DIODE a_45187_38129# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=0p ps=0u w=650000u l=150000u M=8
X10520 a_25287_51157# a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X10521 a_3570_11471# a_2493_11477# a_3408_11849# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10522 VDD pmat.rowon_n[15] a_45178_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10523 a_4437_24643# a_3325_26159# a_4341_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10524 a_45270_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10525 a_35138_9898# pmat.row_n[1] a_35630_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10526 vcm a_18162_9492# a_20170_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10527 VSS a_37129_36130# a_36193_35805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X10528 a_28202_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10529 VSS _1154_.A a_47449_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1053 a_32218_61150# a_18546_61192# a_32126_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10530 VSS pmat.row_n[7] a_27502_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10531 a_31518_55166# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10532 a_31518_13874# nmat.rowon_n[10] a_31122_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10533 a_10045_19677# a_3688_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10534 a_22083_46831# pmat.rowon_n[7] a_21987_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X10535 VDD pmat.rowon_n[14] a_49194_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10536 a_7364_63303# a_7796_62723# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10537 a_39154_11906# a_18162_11500# a_39246_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10538 a_40250_18528# a_18546_18526# a_40158_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10539 a_20267_27497# a_10223_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X1054 a_8013_56085# a_7847_56085# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10540 a_4517_35727# a_4257_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10541 vcm a_18162_64202# a_32218_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10542 VDD a_20316_47607# a_20267_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10543 a_32126_68178# pmat.row_n[12] a_32618_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10544 a_43566_66210# pmat.rowon_n[10] a_43170_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10545 VDD a_1923_61759# a_8175_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10546 a_28110_58138# pmat.row_n[2] a_28602_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10547 a_46848_35951# a_43533_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10548 VDD pmat.rowoff_n[15] a_41162_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10549 VSS a_11339_39319# a_12289_40214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1055 a_4450_23983# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10550 VDD a_47731_36103# a_47592_35643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10551 a_28506_11866# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10552 a_11980_71671# a_11793_71311# a_11893_71427# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X10553 VDD a_40837_46261# a_45966_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10554 a_20170_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10555 a_12199_62621# a_12217_66389# a_12079_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10556 vcm a_18162_14512# a_41254_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10557 VDD a_4429_76751# a_5101_76751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10558 a_9033_27907# a_7140_27805# a_8951_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10559 a_8951_27907# a_7140_27805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1056 a_14336_46983# a_14486_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10560 VDD nmat.rowon_n[14] a_22086_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10561 a_47582_65206# pmat.rowon_n[9] a_47186_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10562 a_5065_69679# a_4991_69831# a_4719_69929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X10563 a_38150_21946# pmat.row_n[13] a_38642_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10564 a_38150_17930# a_18162_17524# a_38242_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10565 a_42258_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10566 VSS a_20315_29098# nmat.col[0] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10567 a_45178_63158# a_18162_63198# a_45270_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10568 a_5865_32687# a_5821_32929# a_5699_32687# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X10569 a_4910_15862# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1057 a_27106_8894# pmat.row_n[0] a_27598_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10570 a_35230_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10571 a_37542_57174# pmat.rowon_n[1] a_37146_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10572 a_30610_57496# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10573 VSS a_27566_43805# a_20438_35431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X10574 vcm a_18162_15516# a_27198_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10575 VDD a_25325_29125# a_25327_28992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10576 VSS a_1643_71829# a_1591_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10577 a_31214_13508# a_18546_13506# a_31122_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10578 a_2203_8585# a_1757_8213# a_2107_8585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X10579 a_8859_22467# a_7779_22583# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X1058 a_11235_26159# a_10791_26409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X10580 pmat.rowoff_n[5] a_13814_59663# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10581 VDD nmat.rowon_n[10] a_48190_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10582 VSS a_22541_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X10583 a_7373_49007# a_6895_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10584 a_22178_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10585 a_12907_13647# a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X10586 a_7578_58294# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10587 VSS pmat.row_n[4] a_30514_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10588 VDD a_2122_19087# a_2228_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10589 a_8113_13353# a_7165_13353# a_8031_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1059 a_36142_57134# pmat.row_n[1] a_36634_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10590 a_36459_29673# a_37291_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10591 a_22482_70226# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10592 VSS a_2263_43719# a_3891_60431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X10593 a_5760_54991# a_5955_55223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10594 a_20078_9898# a_18162_9492# a_20170_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10595 a_44570_8854# nmat.rowon_n[15] a_44174_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10596 a_8841_60405# a_8491_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X10597 a_38546_7850# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10598 a_20078_23954# a_18162_23548# a_20170_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10599 a_43262_72194# a_18546_72236# a_43170_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X106 VDD a_46386_33231# _1194_.A2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u M=16
X1060 vcm a_18162_63198# a_19166_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10600 a_12809_16367# a_11619_16367# a_12700_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X10601 a_36142_24958# nmat.en_bit_n[0] a_36634_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10602 a_39246_62154# a_18546_62196# a_39154_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10603 a_40650_22512# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10604 a_39646_66532# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10605 VSS a_4503_6335# a_4437_6409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X10606 a_33130_22950# a_18162_22544# a_33222_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10607 VDD pmat.rowon_n[8] a_43170_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10608 VDD a_13837_39069# a_13443_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10609 a_28621_47381# a_28455_47381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1061 a_40650_55488# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10610 VSS a_19086_34343# a_19091_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10611 a_10525_12879# a_10471_12791# a_10443_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10612 a_39154_56130# a_18162_56170# a_39246_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10613 a_34924_41605# a_33765_41317# a_34887_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10614 a_25494_61190# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10615 a_32522_62194# pmat.rowon_n[6] a_32126_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10616 a_14864_38567# a_13801_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10617 a_2107_41225# a_1757_40853# a_2012_41213# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X10618 a_34009_28879# a_20439_27247# a_33925_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10619 a_44174_72194# VDD a_44666_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1062 VSS a_40099_52245# pmat.col[20] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10620 a_36142_8894# a_18162_8488# a_36234_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10621 a_7037_70521# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10622 a_41162_14918# a_18162_14512# a_41254_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10623 VSS config_2_in[8] a_1591_41935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10624 a_44666_60508# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10625 a_31015_29111# a_31263_28309# a_31165_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X10626 vcm a_18162_57174# a_30210_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10627 a_4399_51157# a_4175_49667# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10628 a_5320_57863# a_5535_57993# a_5462_58038# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X10629 VDD a_7521_19631# a_5351_19913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=6
X1063 VSS a_46135_38127# a_47223_38671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10630 a_46274_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10631 a_36025_30333# a_35646_29967# a_35953_30333# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10632 a_29510_60186# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10633 VSS a_11927_27399# a_21187_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X10634 VDD a_1586_33927# a_1591_43029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10635 a_29510_19898# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10636 a_41654_7452# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10637 a_31122_70186# a_18162_70226# a_31214_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10638 a_9785_28879# a_9323_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X10639 a_12061_74895# a_10697_75218# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1064 a_46578_20902# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10640 a_30514_14878# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10641 a_4249_9615# a_2021_9563# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10642 VDD VSS a_37146_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10643 a_21574_72556# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10644 a_38242_23548# a_18546_23546# a_38150_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10645 VSS a_36288_44527# a_36394_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10646 VDD a_15420_44007# a_15324_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10647 VDD VDD a_51202_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10648 VDD a_23883_40693# a_23707_40693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10649 a_21082_62154# a_18162_62194# a_21174_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1065 a_19074_67174# pmat.row_n[11] a_19566_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10650 VDD pmat.rowon_n[4] a_21082_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10651 a_34626_71552# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10652 a_42562_67214# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10653 VDD a_29711_47679# a_29698_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10654 VDD VDD a_27106_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10655 VSS VDD a_23486_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10656 a_2882_54991# a_2163_55233# a_2319_54965# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X10657 a_34134_61150# a_18162_61190# a_34226_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10658 a_37542_10862# nmat.rowon_n[13] a_37146_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10659 VDD a_27411_46805# a_27398_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1066 vcm a_18162_23548# a_41254_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10660 a_21031_37217# a_21219_36885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10661 VDD a_13091_52047# a_16863_47428# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10662 VDD pmat.rowoff_n[4] a_24094_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10663 a_33526_7850# VDD a_33130_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10664 a_31539_51946# a_31631_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X10665 a_37404_39429# a_36341_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10666 a_7497_11769# a_2021_9563# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10667 a_46674_18496# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10668 VDD a_6179_69831# a_3936_70197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10669 a_43170_15922# pmat.row_n[7] a_43662_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1067 a_33526_8854# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10670 a_46578_24918# VSS a_46182_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10671 VDD nmat.rowon_n[7] a_50198_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10672 a_11697_56775# a_11902_56775# a_11860_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10673 VDD a_1717_13647# a_8725_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10674 a_7935_20719# a_6981_21263# a_7847_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10675 VSS pmat.row_n[10] a_32522_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10676 VDD a_33395_43455# a_33255_43777# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10677 a_5602_11791# a_5746_11703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10678 VDD a_4298_69367# a_4255_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X10679 a_36538_58178# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1068 a_1846_65579# a_2124_65595# a_2080_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10680 a_45201_47919# a_43315_48437# a_45370_48169# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X10681 a_36538_16886# nmat.rowon_n[7] a_36142_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10682 a_1907_9334# a_1725_9334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10683 a_13236_8573# a_12257_8527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10684 a_19470_68218# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10685 VDD a_21981_34191# a_23807_41959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10686 a_49590_57174# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10687 a_6619_41909# a_6369_39465# a_7005_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10688 a_25098_7890# a_18162_7484# a_25190_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10689 VDD nmat.rowon_n[5] a_23090_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1069 a_23582_65528# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10690 a_51202_67174# a_18162_67214# a_51294_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10691 a_30863_46831# a_30833_46805# a_11067_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X10692 a_3339_70759# a_4075_49007# a_4263_49007# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X10693 vcm a_18162_67214# a_37238_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10694 a_45253_27221# a_16311_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10695 a_11977_66665# a_3923_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10696 a_41254_65166# a_18546_65208# a_41162_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10697 a_14209_52093# a_14174_51859# a_13739_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10698 a_46884_45743# a_29937_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X10699 a_41654_69544# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X107 VSS a_14600_37607# a_23239_37217# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1070 a_20078_62154# pmat.row_n[6] a_20570_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10700 a_37238_55126# a_18546_55168# a_37146_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10701 VDD a_11427_73180# a_11358_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X10702 a_37638_59504# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10703 a_21987_46831# clk_ena a_21797_47081# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10704 a_34226_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10705 a_47290_45717# a_47026_45519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10706 a_48282_7484# a_18546_7482# a_48190_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10707 VSS a_36193_35805# a_35885_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10708 a_11561_40214# a_11389_40443# a_11347_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X10709 a_41162_59142# a_18162_59182# a_41254_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1071 a_49194_56130# pmat.row_n[0] a_49686_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10710 a_5085_59343# a_5053_59575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10711 a_10329_30753# a_10111_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X10712 VSS a_7658_71543# a_9135_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10713 VSS a_1923_61759# a_2369_64061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10714 pmat.row_n[11] a_9963_13967# a_14931_53135# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X10715 a_23700_42919# a_22541_43131# a_23604_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10716 VSS a_2263_43719# a_26933_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10717 a_24094_69182# a_18162_69222# a_24186_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10718 VSS pmat.row_n[1] a_26498_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10719 VDD a_36227_38771# a_36253_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1072 vcm a_18162_13508# a_37238_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10720 a_30514_55166# VSS a_30118_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10721 a_35715_29941# a_35520_30083# a_36025_30333# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X10722 a_17138_46403# a_16083_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10723 VDD a_2983_48071# a_4167_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10724 a_42166_65166# pmat.row_n[9] a_42658_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10725 vcm a_18162_9492# a_29206_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10726 a_44084_52271# ANTENNA__1197__A.DIODE a_43781_52245# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10727 a_27198_66170# a_18546_66212# a_27106_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10728 a_13012_57487# a_12613_57141# a_12341_57141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X10729 VDD nmat.rowon_n[4] a_27106_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1073 a_18563_27791# a_17845_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X10730 VSS a_11207_31764# a_10764_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10731 a_5363_73807# a_4259_73807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X10732 VDD pmat.rowon_n[12] a_31122_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10733 VDD a_3325_36495# a_4181_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10734 VSS a_32827_46805# a_30999_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10735 a_31518_63198# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10736 a_11611_50332# a_11455_50237# a_11756_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X10737 VSS a_11149_40188# a_11093_40214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10738 VSS a_41573_51701# pmat.col_n[21] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10739 VSS a_4871_17429# a_4383_7093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X1074 VDD cgen.dlycontrol4_in[0] a_29627_43983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10740 a_42562_20902# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10741 VSS pmat.row_n[15] a_45574_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10742 VSS a_24407_31375# a_33135_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10743 a_45670_9460# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10744 vcm a_18162_72234# a_32218_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10745 VDD a_8891_66964# a_8723_67191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10746 a_36234_16520# a_18546_16518# a_36142_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10747 a_45178_56130# pmat.row_n[0] a_45670_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10748 vcm a_18162_62194# a_28202_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10749 a_28110_66170# pmat.row_n[10] a_28602_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1075 VSS pmat.row_n[15] a_44570_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10750 vcm a_18162_22544# a_50290_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10751 a_32218_60146# a_18546_60188# a_32126_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10752 a_32618_64524# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10753 a_49286_15516# a_18546_15514# a_49194_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10754 VSS pmat.row_n[7] a_35534_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10755 VDD a_6803_77269# a_6790_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10756 VSS a_4523_21276# a_13367_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.68e+11p ps=1.64e+06u w=420000u l=150000u
X10757 a_23810_47375# a_22733_47381# a_23648_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10758 a_1881_58799# a_1846_59051# a_1643_58773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10759 VDD a_8325_10901# a_8355_11254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1076 a_41254_11500# a_18546_11498# a_41162_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10760 a_22482_23914# pmat.rowoff_n[15] a_22086_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10761 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10762 a_19689_35877# a_18272_35077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X10763 a_29645_47753# a_28455_47381# a_29536_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X10764 a_22578_56492# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10765 a_49194_55126# VDD a_49686_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10766 a_45328_49007# a_44870_48437# a_45238_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X10767 VSS pmat.row_n[14] a_44570_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10768 a_36142_58138# pmat.row_n[2] a_36634_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10769 a_27001_30511# a_24861_29673# a_27181_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1077 a_2319_52789# a_2124_52931# a_2629_53181# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X10770 a_22365_32149# a_22199_32149# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X10771 a_33130_60146# pmat.row_n[4] a_33622_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10772 a_36538_11866# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10773 a_42258_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10774 VSS a_13459_28111# a_47120_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10775 a_19470_21906# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10776 a_15667_27239# a_43659_28853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X10777 a_49590_10862# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10778 VDD a_17996_36391# a_17900_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10779 a_26594_55488# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1078 a_46043_43343# a_40105_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=0p ps=0u w=650000u l=150000u M=2
X10780 vcm a_18162_23548# a_27198_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10781 a_25815_43957# a_10873_39605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10782 a_6975_76823# a_9287_77055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10783 VSS pmat.row_n[5] a_47582_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10784 a_21478_70226# pmat.rowon_n[14] a_21082_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10785 a_31214_21540# a_18546_21538# a_31122_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10786 a_35717_28111# a_26891_28327# a_35499_28023# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10787 VDD a_9367_53511# a_7163_53333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X10788 a_51598_18894# nmat.rowon_n[5] a_51202_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10789 a_27198_11500# a_18546_11498# a_27106_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1079 a_33130_61150# pmat.row_n[5] a_33622_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10790 VDD a_7631_15253# a_7618_15645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10791 VDD nmat.en_bit_n[2] a_35138_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10792 a_29114_9898# a_18162_9492# a_29206_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10793 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10794 a_29109_38571# a_23821_35279# a_29023_38571# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X10795 a_29510_13874# nmat.rowon_n[10] a_29114_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10796 VSS pmat.row_n[2] a_26498_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10797 vcm a_18162_59182# a_48282_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10798 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10799 a_5248_30511# a_4167_30511# a_4901_30753# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X108 a_34134_65166# a_18162_65206# a_34226_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1080 a_36538_12870# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10800 VDD a_11339_39319# a_12757_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X10801 a_7631_75895# a_6795_76989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10802 a_49194_72194# a_18162_72234# a_49286_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10803 a_48586_16886# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10804 a_5578_54991# a_4075_68583# a_5329_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5e+11p pd=2.5e+06u as=3.85e+11p ps=2.77e+06u w=1e+06u l=150000u
X10805 a_39246_70186# a_18546_70228# a_39154_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10806 a_31122_63158# pmat.row_n[7] a_31614_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10807 VDD a_9375_72007# a_11014_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10808 nmat.col[18] ANTENNA__1183__B1.DIODE a_82735_2223# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=7.085e+11p ps=7.38e+06u w=650000u l=150000u M=2
X10809 a_36634_20504# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1081 a_42258_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10810 VDD pmat.rowoff_n[15] a_39154_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10811 a_5179_31591# a_1781_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X10812 a_35138_18934# pmat.row_n[10] a_35630_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10813 VDD VDD a_43170_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10814 a_36234_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10815 a_36895_29673# pmat.sw a_10147_29415# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=0p ps=0u w=1e+06u l=150000u
X10816 nmat.col[21] ANTENNA__1187__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10817 a_14103_15936# a_12447_16143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10818 a_39154_64162# a_18162_64202# a_39246_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10819 a_43262_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1082 a_18546_66212# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X10820 a_5275_65327# a_5595_65301# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=150000u
X10821 a_2672_16201# a_1591_15829# a_2325_15797# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10822 a_26194_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10823 a_28506_60186# pmat.rowon_n[4] a_28110_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10824 pmat.col_n[6] ANTENNA__1190__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10825 VDD a_8175_12533# a_5579_12394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10826 a_28506_19898# nmat.rowon_n[4] a_28110_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10827 a_4712_27023# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X10828 VDD a_17625_42902# a_16689_43132# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X10829 VDD a_39359_49172# a_38695_48634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1083 a_50290_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10830 a_13988_55369# a_13073_54997# a_13641_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X10831 VDD a_9411_15831# a_3571_13627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10832 a_41162_22950# a_18162_22544# a_41254_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10833 a_8356_23671# a_4703_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10834 VDD a_30155_36893# a_30181_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X10835 a_12990_13967# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10836 a_37146_12910# a_18162_12504# a_37238_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10837 a_38569_46831# a_11948_49783# a_38581_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10838 a_46578_7850# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10839 a_53622_39932# comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top comp.adc_comp_circuit_0.adc_comp_buffer_1.in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.24e+12p ps=9.24e+06u w=2e+06u l=150000u M=2
X1084 VSS pmat.row_n[2] a_40554_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10840 a_33222_68178# a_18546_68220# a_33130_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10841 VSS pmat.row_n[13] a_37542_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10842 vcm a_18162_65206# a_30210_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10843 a_30118_69182# pmat.row_n[13] a_30610_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10844 a_21977_52245# _1194_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10845 a_29206_58138# a_18546_58180# a_29114_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10846 a_41558_67214# pmat.rowon_n[11] a_41162_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10847 VSS pmat.row_n[1] a_39550_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10848 a_51294_18528# a_18546_18526# a_51202_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10849 VDD a_11261_41245# a_10867_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1085 VDD a_38851_28327# a_43451_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X10850 VDD a_5351_19913# a_14477_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10851 a_5256_42301# a_5134_41909# a_5184_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10852 VSS pmat.row_n[9] a_50594_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10853 vcm a_18162_10496# a_26194_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10854 a_24719_37429# a_11497_38543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10855 a_4768_16055# a_3688_17179# a_4910_15862# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X10856 a_5318_28701# a_4241_28335# a_5156_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10857 a_20879_47893# a_21215_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X10858 a_38546_65206# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10859 a_31214_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1086 VSS a_4989_11079# a_5012_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.3925e+11p ps=9.39e+06u w=650000u l=150000u M=2
X10860 VSS a_18547_51565# a_18660_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10861 a_27198_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10862 VSS a_34942_51701# a_36631_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10863 vcm a_18162_56170# a_51294_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10864 VDD a_13653_40956# a_13259_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10865 a_21478_24918# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10866 a_51598_13874# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10867 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10868 a_2215_34141# a_1591_33775# a_2107_33775# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X10869 a_35534_58178# pmat.rowon_n[2] a_35138_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1087 a_19470_22910# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10870 a_21981_34191# a_21815_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X10871 a_17187_49783# a_17459_49641# a_17417_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10872 a_34530_23914# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10873 a_2858_72531# a_3136_72515# a_3092_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10874 a_38642_61512# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10875 a_14649_16911# a_10515_15055# a_14565_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10876 vcm a_18162_16520# a_25190_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10877 a_28202_19532# a_18546_19530# a_28110_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10878 a_46274_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10879 a_48586_57174# pmat.rowon_n[1] a_48190_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1088 VSS pmat.row_n[12] a_23486_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10880 a_43170_66170# a_18162_66210# a_43262_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10881 a_17996_44007# a_16837_44219# a_17959_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10882 a_13140_50247# a_13290_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10883 a_7118_32509# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10884 a_28613_40229# a_28116_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X10885 a_10321_20291# a_4523_21276# a_10239_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10886 a_24490_15882# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10887 a_2834_38671# a_1757_38677# a_2672_39049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10888 a_12471_39126# a_12289_39126# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10889 a_24490_9858# nmat.rowon_n[14] a_24094_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1089 a_41121_30511# a_28704_29568# a_41049_30511# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10890 a_50594_60186# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10891 a_50594_19898# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10892 VDD a_11435_58791# a_14103_15936# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10893 VSS pmat.row_n[10] a_40554_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10894 a_33526_70226# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10895 a_37238_63158# a_18546_63200# a_37146_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10896 a_36617_36603# a_34924_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X10897 a_37638_67536# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10898 VDD pmat.rowon_n[9] a_41162_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10899 a_35230_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X109 a_37542_14878# nmat.rowon_n[9] a_37146_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1090 a_26594_56492# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10900 a_47186_24958# VDD a_47678_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10901 a_10999_39958# a_10817_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10902 a_11159_28585# a_9741_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10903 a_10219_30877# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10904 a_37146_57134# a_18162_57174# a_37238_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10905 VDD a_17927_48437# pmat.row_n[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10906 a_7645_53909# a_7479_53909# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X10907 a_51694_22512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10908 a_22576_30511# a_22628_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=0p ps=0u w=650000u l=150000u M=4
X10909 a_23486_62194# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1091 a_12595_31433# a_12245_31061# a_12500_31421# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X10910 a_41254_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10911 VDD a_2046_30184# a_4167_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10912 a_30514_63198# pmat.rowon_n[7] a_30118_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10913 VDD pmat.rowon_n[4] a_19074_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10914 a_6464_71855# a_6200_70919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10915 a_13073_54997# a_12907_54997# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X10916 VDD a_10839_11989# a_11207_11079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10917 VSS pmat.row_n[14] a_37542_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10918 a_9953_53903# a_9581_56079# a_9871_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X10919 VDD a_39781_40157# a_39387_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1092 _1154_.A a_37471_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X10920 a_41654_14480# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10921 VDD nmat.rowon_n[6] a_44174_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10922 a_41558_20902# pmat.rowoff_n[12] a_41162_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10923 a_83166_9839# ANTENNA__1190__A1.DIODE a_82788_9991# VSS sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=3.25e+11p ps=2.3e+06u w=650000u l=150000u
X10924 a_24586_24520# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10925 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10926 a_21574_8456# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10927 VSS a_7779_22583# a_9135_22057# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10928 VDD a_20475_49783# a_22265_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10929 a_27198_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1093 VDD a_38972_39655# a_38876_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X10930 a_2871_51701# a_2715_51969# a_3016_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X10931 nmat.col[13] _1183_.A2 a_14747_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10932 a_4535_74031# a_4505_74005# a_4441_74031# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X10933 a_4319_71311# a_2727_58470# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10934 a_36234_24552# a_18546_24550# a_36142_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10935 a_45670_13476# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10936 a_35230_66170# a_18546_66212# a_35138_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10937 a_42166_10902# pmat.row_n[2] a_42658_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10938 vcm a_18162_70226# a_28202_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10939 VDD nmat.rowon_n[15] a_31122_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1094 a_10864_68565# a_10391_69653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10940 VDD VSS a_48190_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10941 a_28602_23516# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10942 a_25098_20942# pmat.row_n[12] a_25590_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10943 a_40554_68218# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10944 a_25098_16926# a_18162_16520# a_25190_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10945 a_28202_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10946 a_49286_23548# a_18546_23546# a_49194_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10947 VSS a_13985_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X10948 a_32618_72556# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10949 a_16764_47081# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1095 a_21478_71230# pmat.rowon_n[15] a_21082_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10950 VDD nmat.rowon_n[2] a_32126_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10951 VDD pmat.rowon_n[2] a_35138_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10952 a_14369_50345# a_11711_50959# a_14287_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10953 a_35534_11866# nmat.rowon_n[12] a_35138_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10954 a_32126_62154# a_18162_62194# a_32218_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10955 VSS a_4259_73807# a_4893_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10956 a_24490_56170# pmat.rowon_n[0] a_24094_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10957 VDD a_6343_18517# a_6330_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10958 VSS start_conversion_in a_1591_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10959 VDD nmat.rowon_n[10] a_22086_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1096 VSS pmat.row_n[14] a_48586_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10960 a_48586_10862# nmat.rowon_n[13] a_48190_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10961 VDD a_23301_47349# a_23191_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10962 vcm a_18162_62194# a_36234_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10963 a_2405_19087# a_2228_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10964 a_36142_66170# pmat.row_n[10] a_36634_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10965 a_40250_60146# a_18546_60188# a_40158_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10966 a_40650_64524# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10967 a_43566_59182# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10968 a_29114_15922# a_18162_15516# a_29206_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10969 a_2325_23413# a_2107_23817# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X1097 a_31214_22544# a_18546_22542# a_31122_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10970 VDD cgen.dlycontrol2_in[4] a_29163_38545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10971 vcm a_18162_61190# a_49286_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10972 a_1761_6031# a_1591_6031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X10973 a_33222_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10974 a_8655_64783# a_8031_64789# a_8547_65161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10975 a_3202_29941# a_3052_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.184e+11p pd=2.2e+06u as=0p ps=0u w=840000u l=150000u
X10976 a_19074_11906# pmat.row_n[3] a_19566_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10977 a_36854_44527# a_36677_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10978 vcm a_18162_8488# a_42258_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10979 a_4885_58255# a_1823_60949# a_4801_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 VSS a_14249_49525# a_12044_49641# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X10980 a_30210_71190# a_18546_71232# a_30118_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10981 a_47582_58178# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10982 a_41791_51727# a_21739_29415# a_41573_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10983 VDD a_11149_40188# a_11561_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10984 a_41162_60146# pmat.row_n[4] a_41654_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10985 a_26194_61150# a_18546_61192# a_26102_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10986 VDD pmat.rowon_n[12] a_29114_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10987 a_34797_27791# a_24591_28327# nmat.col[14] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10988 a_6909_21263# a_3305_17999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10989 VSS a_4737_23957# a_4671_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1099 a_27198_12504# a_18546_12502# a_27106_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10990 VDD pmat.rowon_n[7] a_30118_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10991 a_6742_10499# a_2021_9563# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10992 a_40567_32403# a_40903_32375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10993 a_9129_27907# a_9075_28023# a_9033_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10994 vcm a_18162_67214# a_48282_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10995 VSS a_9075_28023# a_8951_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10996 a_3880_70543# a_3838_70455# a_3577_70197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10997 a_3881_68047# a_2727_58470# a_3069_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10998 VSS a_2511_25615# a_1923_31743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X10999 a_28202_8488# a_18546_8486# a_28110_8894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11 a_45178_69182# a_18162_69222# a_45270_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X110 a_5573_12015# a_5173_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1100 VSS a_12407_28853# a_12437_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X11000 VDD a_22199_30287# a_27903_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11001 a_13347_64783# a_12723_64789# a_13239_65161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11002 a_3987_47375# a_3799_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11003 VSS pmat.row_n[15] a_38546_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11004 VSS pmat.row_n[2] a_24490_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11005 a_35230_11500# a_18546_11498# a_35138_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11006 a_20629_32521# a_19439_32149# a_20520_32521# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X11007 a_31122_71190# pmat.row_n[15] a_31614_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11008 VSS a_2944_52789# a_2882_52815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11009 a_27106_61150# pmat.row_n[5] a_27598_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1101 a_46274_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11010 a_3795_70223# a_3936_70197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11011 a_36234_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11012 a_35138_69182# a_18162_69222# a_35230_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11013 a_48282_10496# a_18546_10494# a_48190_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11014 a_37404_38341# a_36341_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11015 VDD a_7693_22365# a_12051_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11016 a_84028_9615# _1196_.B1 a_83839_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X11017 a_10851_30485# a_10676_30511# a_11030_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11018 a_39246_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11019 VSS a_82787_14709# nmat.col_n[18] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u M=2
X1102 a_43170_20942# a_18162_20536# a_43262_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11020 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11021 VDD a_10764_32117# a_10702_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11022 a_10641_52815# a_10363_53153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X11023 VSS a_1586_18231# a_1591_20181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11024 a_14458_4399# a_9411_2215# a_14372_4399# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X11025 a_25190_22544# a_18546_22542# a_25098_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11026 VDD a_8851_63669# a_8782_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11027 VSS a_26957_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X11028 a_40554_21906# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11029 VSS VDD a_43566_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1103 a_6406_26159# a_6634_26133# a_6664_26159# VSS sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X11030 a_37146_20942# a_18162_20536# a_37238_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11031 a_29825_30557# a_29455_31293# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11032 a_1674_57711# a_1644_57685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X11033 a_42791_32375# a_44082_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11034 a_43170_57134# pmat.row_n[1] a_43662_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11035 VDD a_2215_47375# a_7521_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X11036 VSS a_25802_48169# a_27020_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X11037 VDD a_5248_30511# a_5423_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11038 VSS a_14589_40726# a_13653_40956# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X11039 a_42683_32375# a_42791_32375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1104 VDD a_5579_12394# a_5541_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X11040 a_47278_16520# a_18546_16518# a_47186_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11041 VSS a_39013_43655# a_40315_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11042 a_11987_23983# a_11897_21263# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.85e+11p pd=5.7e+06u as=0p ps=0u w=650000u l=150000u
X11043 a_28336_29967# a_18563_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X11044 VSS a_25639_43957# a_12197_43746# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11045 a_19470_70226# pmat.rowon_n[14] a_19074_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11046 a_7456_15279# a_6541_15279# a_7109_15521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11047 a_42151_50095# a_24867_53135# pmat.col[23] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X11048 a_33222_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11049 a_30118_55126# a_18162_55166# a_30210_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1105 a_3762_11837# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X11050 VDD a_13973_66933# a_14001_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X11051 a_5553_65577# a_5495_65479# a_5138_65479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11052 VSS pmat.row_n[7] a_46578_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11053 a_49590_18894# nmat.rowon_n[5] a_49194_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11054 a_20570_18496# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11055 a_20474_24918# nmat.en_C0_n a_20078_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11056 a_17959_44265# a_16837_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11057 a_43566_12870# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11058 a_22225_46653# a_13275_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11059 a_50594_13874# nmat.rowon_n[10] a_50198_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1106 VSS pmat.row_n[6] a_38546_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11060 VSS nmat.sw a_12191_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11061 a_30409_48463# a_29076_48695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X11062 a_10070_32143# a_9944_32259# a_9666_32275# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11063 VSS a_2199_13887# a_6205_5487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11064 a_30118_14918# pmat.row_n[6] a_30610_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11065 a_33622_17492# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11066 a_33526_23914# pmat.rowoff_n[15] a_33130_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11067 a_31122_18934# a_18162_18528# a_31214_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11068 vcm a_18162_64202# a_51294_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11069 VDD a_5779_71285# a_7044_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1107 a_20474_8854# nmat.rowon_n[15] a_20078_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11070 VSS a_37129_36130# a_37739_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11071 a_51202_68178# pmat.row_n[12] a_51694_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11072 VDD a_28915_50959# a_47591_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11073 a_47186_58138# pmat.row_n[2] a_47678_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11074 VSS pmat.row_n[9] a_19470_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11075 a_2834_20175# a_1757_20181# a_2672_20553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11076 a_13896_74953# a_12815_74581# a_13549_74549# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11077 a_23486_15882# pmat.rowoff_n[7] a_23090_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11078 VSS a_4523_21276# a_10651_24617# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11079 a_7933_31433# a_6743_31061# a_7824_31433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1108 VDD a_24833_40719# a_30155_42583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11080 a_47582_11866# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11081 a_8693_11769# a_2021_11043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11082 a_11071_46805# a_11506_47083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11083 vcm a_18162_24552# a_25190_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11084 a_6343_32661# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11085 a_34134_13914# pmat.row_n[5] a_34626_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11086 a_35230_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11087 vcm a_18162_66210# a_24186_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11088 a_10391_62911# a_10216_62985# a_10570_62973# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11089 a_18546_11498# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X1109 a_40250_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11090 a_16745_44581# a_13779_43123# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11091 VDD a_13563_24527# a_13683_24847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11092 a_24586_58500# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11093 a_27502_14878# nmat.rowon_n[9] a_27106_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11094 VSS pmat.row_n[3] a_24490_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11095 VSS a_26317_40726# a_26515_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11096 a_30219_29967# a_29968_30083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11097 VDD VSS a_46182_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11098 VSS a_7644_16341# a_11995_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11099 a_17842_27497# a_7415_29397# a_16965_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X111 nmat.col[21] _1187_.A2 a_83217_4649# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u M=4
X1110 a_42562_60186# pmat.rowon_n[4] a_42166_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11100 VSS _1184_.A2 a_33412_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X11101 VDD a_20616_27791# a_22979_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X11102 a_2781_16201# a_1591_15829# a_2672_16201# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11103 a_39550_67214# pmat.rowon_n[11] a_39154_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11104 VSS pmat.row_n[8] a_36538_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11105 a_14441_57711# a_12447_16143# a_14369_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11106 vcm a_18162_15516# a_46274_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11107 a_27236_46831# a_26321_46831# a_26889_47073# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11108 a_50290_13508# a_18546_13506# a_50198_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11109 VSS a_11693_70767# a_12052_71671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1111 a_42562_19898# nmat.rowon_n[4] a_42166_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11110 a_4162_64561# a_2419_53351# a_4161_64239# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11111 VSS a_4031_40455# a_3199_40455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11112 a_37146_65166# a_18162_65206# a_37238_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11113 a_44174_8894# pmat.row_n[0] a_44666_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11114 a_33395_32463# a_30278_30511# a_33205_32143# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11115 a_41254_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11116 a_47678_20504# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11117 VSS a_20848_36165# a_20811_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11118 a_47278_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11119 a_38546_8854# nmat.rowon_n[15] a_38150_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1112 a_2858_59475# a_3175_59585# a_3133_59709# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X11120 a_26425_32463# a_11067_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11121 a_41558_70226# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11122 a_50594_8854# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11123 vcm a_18162_17524# a_19166_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11124 a_4921_32441# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11125 a_38515_49035# ANTENNA_fanout52_A.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11126 a_23182_15516# a_18546_15514# a_23090_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11127 vcm a_18162_12504# a_20170_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11128 VSS a_4351_55527# a_4903_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X11129 a_37638_12472# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1113 a_25494_70226# pmat.rowon_n[14] a_25098_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11130 a_1925_26935# a_2021_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11131 VDD nmat.rowon_n[13] a_41162_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11132 a_26498_8854# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11133 a_14708_31599# a_4707_32156# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X11134 a_6877_37039# a_6833_37281# a_6711_37039# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11135 a_48190_12910# a_18162_12504# a_48282_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11136 VSS a_3859_22655# a_3793_22729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X11137 a_27198_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11138 a_44570_61190# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11139 VSS a_12061_26703# a_21365_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1114 a_48586_17890# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11140 VDD a_22933_32117# a_22823_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11141 a_27502_71230# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11142 vcm a_18162_11500# a_24186_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11143 VSS a_16863_52815# pmat.rowon_n[0] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X11144 a_2191_27412# a_2283_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11145 VSS a_6608_60663# a_5053_59575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11146 a_25098_24958# a_18162_24552# a_25190_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11147 VDD pmat.rowon_n[10] a_35138_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11148 a_11292_39631# a_11041_39860# a_11071_39958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11149 a_35230_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1115 a_27794_28879# a_27355_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X11150 a_28110_60146# a_18162_60186# a_28202_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11151 a_31053_47081# a_31105_46805# a_11067_49871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X11152 VSS pmat.row_n[5] a_21478_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11153 cgen.dlycontrol4_in[4] a_2235_23983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11154 VDD a_4351_55527# a_4809_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X11155 a_18162_66210# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11156 vcm a_18162_70226# a_36234_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11157 a_47212_29673# a_41731_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X11158 a_27531_51727# ANTENNA__1395__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11159 a_9103_73791# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1116 a_39246_71190# a_18546_71232# a_39154_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11160 a_32522_24918# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11161 a_40650_72556# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11162 a_7169_15055# a_5266_17143# a_7085_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11163 a_2499_13077# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11164 a_29114_23954# a_18162_23548# a_29206_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11165 a_23707_34165# a_11225_35836# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11166 VDD pmat.rowon_n[9] a_39154_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11167 a_36634_62516# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11168 a_3305_62607# a_3345_62839# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11169 a_46578_58178# pmat.rowon_n[2] a_46182_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1117 a_10049_60663# a_10391_62911# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11170 VDD pmat.rowon_n[4] a_40158_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11171 vcm a_18162_59182# a_22178_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11172 a_25325_29125# a_23933_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11173 a_11433_69679# a_11391_69831# a_8439_69653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X11174 a_34828_39429# a_33765_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11175 VDD a_12449_22895# a_14778_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11176 a_33130_7890# VDD a_33622_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11177 a_49686_61512# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11178 VSS pmat.row_n[4] a_25494_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11179 a_22482_16886# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1118 a_2121_55357# a_1643_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11180 VSS pmat.row_n[11] a_25494_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11181 ANTENNA__1395__A1.DIODE a_47591_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11182 a_8695_63937# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11183 a_32947_38825# a_33341_38780# a_33007_38771# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11184 a_42191_48071# a_35186_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11185 VDD cgen.enable_dlycontrol_in a_23655_35279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11186 a_6060_49007# a_5785_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11187 a_20078_10902# a_18162_10496# a_20170_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11188 a_39550_20902# pmat.rowoff_n[12] a_39154_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11189 a_35534_15882# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1119 VDD VSS a_39154_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11190 a_3202_29941# a_3052_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X11191 a_9217_26409# a_2952_25045# a_9135_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11192 a_14607_26703# a_12449_22895# a_14499_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.4e+11p pd=2.88e+06u as=0p ps=0u w=1e+06u l=150000u
X11193 VSS a_40628_39429# a_39781_40157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X11194 vcm a_18162_58178# a_26194_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11195 VDD pmat.rowon_n[15] a_30118_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11196 VSS a_7730_69109# a_8538_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11197 a_37007_52521# a_34705_51959# a_36789_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11198 VDD pmat.rowon_n[5] a_26102_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11199 a_8569_60405# a_8841_60405# a_9240_60751# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X112 a_32827_46805# a_33467_46261# a_33239_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X1120 nmat.col[23] a_27763_27221# a_41703_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X11200 a_12689_29199# a_6830_22895# a_12605_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11201 a_30210_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11202 a_12021_53609# a_9463_53511# a_11925_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X11203 VSS pmat.row_n[10] a_51598_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11204 VDD a_2129_12559# a_3158_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11205 VSS a_25473_52245# pmat.col[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11206 a_48190_57134# a_18162_57174# a_48282_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11207 VDD VDD a_20078_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11208 a_24094_11906# a_18162_11500# a_24186_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11209 a_4910_16189# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1121 a_43262_58138# a_18546_58180# a_43170_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11210 a_25287_32117# clk_ena a_25718_32463# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X11211 a_45837_27791# a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X11212 a_7037_70521# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11213 VDD nmat.rowon_n[5] a_42166_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11214 nmat.col[24] ANTENNA__1190__B1.DIODE a_82736_4943# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11215 a_6607_10615# a_2021_9563# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11216 VSS a_1828_25589# a_1858_25615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X11217 a_15368_31599# a_14287_31599# a_15021_31841# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X11218 a_50198_15922# a_18162_15516# a_50290_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11219 VSS a_1923_69823# a_1881_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1122 vcm a_18162_55166# a_40250_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11220 a_2007_8916# a_2099_8725# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11221 a_12270_30838# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X11222 VSS pmat.row_n[1] a_45574_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11223 a_39154_16926# pmat.row_n[8] a_39646_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11224 VDD a_40837_46261# a_45475_35520# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11225 a_25893_49551# a_25839_49783# pmat.rowoff_n[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11226 VSS pmat.row_n[11] a_28506_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11227 a_40158_11906# pmat.row_n[3] a_40650_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11228 VSS a_11067_64015# a_17478_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11229 a_25494_64202# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1123 a_40158_59142# pmat.row_n[3] a_40650_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11230 a_32522_65206# pmat.rowon_n[9] a_32126_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11231 nmat.rowon_n[9] a_13446_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11232 a_23090_21946# pmat.row_n[13] a_23582_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11233 a_14439_72703# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11234 a_23090_17930# a_18162_17524# a_23182_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11235 a_47278_24552# a_18546_24550# a_47186_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11236 a_46274_66170# a_18546_66212# a_46182_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11237 a_17845_27791# a_7840_27247# a_17323_28111# VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X11238 VDD pmat.rowon_n[12] a_50198_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11239 a_30118_63158# a_18162_63198# a_30210_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1124 VDD a_21037_43658# a_12228_40693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11240 VSS a_2315_44124# a_4175_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11241 VDD pmat.rowon_n[2] a_46182_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11242 a_20170_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11243 a_22482_57174# pmat.rowon_n[1] a_22086_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11244 a_10999_38870# a_10817_38870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11245 a_2242_44477# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11246 a_39646_9460# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11247 a_46578_11866# nmat.rowon_n[12] a_46182_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11248 a_7497_11769# a_2021_9563# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11249 a_2659_35015# a_5558_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1125 VDD a_15753_28879# a_24131_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X11250 a_6711_37039# a_6265_37039# a_6615_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11251 a_29606_15484# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11252 a_41254_7484# a_18546_7482# a_41162_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11253 vcm a_18162_72234# a_51294_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11254 VDD nmat.rowon_n[10] a_33130_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11255 a_4831_34561# a_1586_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11256 a_17113_35877# a_13503_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X11257 vcm a_18162_62194# a_47278_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11258 a_47186_66170# pmat.row_n[10] a_47678_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11259 a_35077_50345# a_30571_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1126 VDD a_18823_50247# a_19584_52423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11260 a_2122_17455# a_1945_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11261 a_51294_60146# a_18546_60188# a_51202_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11262 a_11241_23145# a_6173_22895# a_11159_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11263 a_76962_40202# a_77058_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11264 a_51694_64524# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11265 a_19470_55166# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11266 VDD a_46135_38127# a_47223_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11267 a_5038_28853# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11268 VDD a_2325_15797# a_2215_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11269 nmat.rowoff_n[5] nmat.rowon_n[7] a_14195_11791# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1127 a_4955_40277# a_7079_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11270 vcm a_18162_9492# a_22178_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11271 a_17033_51183# a_16679_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11272 a_10867_38007# a_11261_37981# a_10927_37981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11273 a_41654_56492# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11274 a_21082_24958# VDD a_21574_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11275 a_24186_62154# a_18546_62196# a_24094_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11276 a_22541_38779# a_22085_38550# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11277 VDD a_40105_47375# a_46233_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X11278 VDD pmat.rowon_n[13] a_27106_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11279 VDD a_38913_31055# a_41475_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1128 a_20063_32143# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11280 a_24586_66532# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11281 a_32218_9492# a_18546_9490# a_32126_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11282 a_42258_12504# a_18546_12502# a_42166_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11283 a_16745_34427# a_15144_35077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11284 a_24094_56130# a_18162_56170# a_24186_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11285 a_2375_63316# a_2467_63125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11286 VSS a_2319_54965# a_2250_54991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X11287 VDD a_13641_54965# a_13531_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X11288 VSS a_3199_53877# a_3111_53333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11289 VSS a_5325_9269# a_4989_11079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1129 a_28506_61190# pmat.rowon_n[5] a_28110_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11290 VSS VDD a_36538_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11291 a_45670_55488# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11292 VDD a_14249_49525# a_12044_49641# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11293 vcm a_18162_23548# a_46274_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11294 VSS a_22499_49783# a_37471_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11295 a_40554_70226# pmat.rowon_n[14] a_40158_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11296 a_28602_65528# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11297 a_25098_62154# pmat.row_n[6] a_25590_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11298 a_50290_21540# a_18546_21538# a_50198_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11299 VDD a_1586_8439# a_1591_8213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X113 VSS a_5081_53135# a_6334_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1130 a_24753_42919# a_25061_43132# a_11389_40443# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X11300 a_20184_46983# a_20267_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11301 VSS a_1923_69823# a_3473_77117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11302 a_18546_19530# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11303 VSS pmat.row_n[15] a_49590_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11304 a_46274_11500# a_18546_11498# a_46182_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11305 a_4863_13077# a_2648_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X11306 VSS a_10699_72943# a_11345_70773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11307 VDD nmat.rowon_n[14] a_24094_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11308 a_28116_38567# a_26957_38779# a_28020_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11309 a_47278_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1131 a_18823_50247# a_25839_49783# a_26242_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X11310 VDD a_9869_69921# a_9759_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11311 VDD a_43781_52245# pmat.col_n[24] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11312 VSS pmat.row_n[2] a_45574_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11313 VSS a_22357_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X11314 VDD a_2319_74268# a_2250_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X11315 VDD a_18272_35077# a_18176_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X11316 VDD VSS a_22086_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11317 a_12092_42895# a_11915_42895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11318 VSS pmat.row_n[12] a_28506_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11319 a_2847_28095# a_2672_28169# a_3026_28157# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1132 a_14287_15529# a_10515_61839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X11320 vcm a_18162_20536# a_20170_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11321 a_23182_23548# a_18546_23546# a_23090_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11322 a_43566_61190# pmat.rowon_n[5] a_43170_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11323 a_19166_13508# a_18546_13506# a_19074_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11324 a_24591_28327# a_40567_32403# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X11325 a_26498_71230# pmat.rowon_n[15] a_26102_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11326 a_25695_28111# a_42307_31756# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11327 a_31925_40955# a_31469_40726# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11328 a_22206_31094# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X11329 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1133 a_43533_30761# a_41227_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.62e+12p pd=1.524e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X11330 a_41877_30761# a_40969_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11331 a_13529_34951# a_13801_34427# a_14864_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11332 a_3295_40277# a_2935_38279# a_3514_40079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X11333 a_4028_65871# a_3814_65871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11334 a_48190_20942# a_18162_20536# a_48282_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11335 a_7847_24233# a_7779_22583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11336 a_22482_10862# nmat.rowon_n[13] a_22086_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11337 a_11203_62037# a_11713_64899# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11338 a_44266_59142# a_18546_59184# a_44174_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11339 VDD a_35039_29941# a_31263_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1134 a_5043_37191# a_2659_35015# a_5277_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11340 a_45270_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11341 a_47582_60186# pmat.rowon_n[4] a_47186_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11342 a_19584_52423# a_18823_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11343 a_47582_19898# nmat.rowon_n[4] a_47186_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11344 VSS pmat.row_n[8] a_44570_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11345 a_22086_9898# a_18162_9492# a_22178_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11346 cgen.dlycontrol3_in[3] a_2235_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11347 a_42258_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11348 a_14753_27247# a_14691_27399# a_14637_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=2.795e+11p ps=2.16e+06u w=650000u l=150000u
X11349 VDD a_30140_43781# a_30044_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1135 a_6747_25731# a_3305_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X11350 a_31614_18496# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11351 a_31518_24918# VSS a_31122_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11352 a_35230_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11353 a_32218_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11354 a_48282_58138# a_18546_58180# a_48190_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11355 vcm a_18162_55166# a_45270_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11356 a_45178_59142# pmat.row_n[3] a_45670_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11357 a_21478_58178# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11358 a_20752_42693# a_19689_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11359 VDD a_2195_51701# a_1823_58237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1136 VSS a_3659_39733# a_3295_40277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X11360 a_21478_16886# nmat.rowon_n[7] a_21082_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11361 a_21032_44007# a_19873_44219# a_20936_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11362 VDD a_19487_49159# a_18359_49140# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X11363 a_34530_57174# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11364 a_36634_70548# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11365 a_46815_37013# a_43776_30287# a_47084_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11366 a_26659_34967# a_24833_34191# a_26833_35073# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11367 vcm a_18162_67214# a_22178_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11368 a_20173_32117# a_19955_32521# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11369 a_4677_70561# a_2419_53351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1137 VDD VDD a_47186_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11370 a_12969_40175# a_12543_40214# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11371 a_6082_46831# a_5455_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11372 a_36142_60146# a_18162_60186# a_36234_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11373 a_12250_4175# _1194_.A2 a_12081_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11374 a_50290_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11375 vcm a_18162_17524# a_40250_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11376 a_22178_55126# a_18546_55168# a_22086_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11377 a_5535_57993# a_9305_58229# a_9335_58575# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u M=2
X11378 VDD a_33845_27765# nmat.col_n[14] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11379 a_19074_70186# a_18162_70226# a_19166_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1138 a_22178_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11380 vcm a_18162_66210# a_35230_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11381 a_22578_59504# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11382 a_46274_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11383 a_19965_39867# a_19509_39638# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X11384 a_45557_35773# a_40837_46261# a_45475_35520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11385 a_47806_47081# ANTENNA__1197__B.DIODE a_47724_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11386 VDD a_13203_70767# a_13605_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11387 a_5461_67753# a_5403_67655# a_5046_67655# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X11388 a_5736_56399# a_5682_56311# a_5245_56053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11389 a_15420_44007# a_14261_44219# a_15383_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1139 a_2107_36873# a_1757_36501# a_2012_36861# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11390 a_48282_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11391 a_43662_7452# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11392 VSS a_44811_36469# a_17139_30503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=8
X11393 VDD nmat.rowon_n[13] a_39154_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11394 VSS a_31323_29967# a_31399_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11395 a_13985_34789# a_13529_34951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X11396 a_37542_68218# pmat.rowon_n[12] a_37146_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11397 vcm a_18162_16520# a_44266_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11398 a_5510_28335# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11399 VSS pmat.row_n[8] a_47582_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 VSS pmat.row_n[0] a_23486_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1140 a_33222_69182# a_18546_69224# a_33130_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11400 VDD VDD a_29114_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11401 VSS VDD a_25494_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11402 a_13795_10687# a_13620_10761# a_13974_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11403 VDD a_10697_75218# a_9831_74183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11404 a_20400_40719# a_14533_39631# a_20179_41046# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11405 a_48190_65166# a_18162_65206# a_48282_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11406 a_9510_9839# a_1717_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11407 VDD a_2419_53351# a_3621_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11408 VSS pmat.row_n[15] a_30514_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11409 a_30514_9858# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1141 vcm a_18162_66210# a_30210_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11410 VDD a_1643_56597# a_1591_56623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11411 VSS pmat.row_n[0] a_37542_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11412 VDD pmat.rowon_n[5] a_34134_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11413 a_21174_16520# a_18546_16518# a_21082_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11414 a_7578_58621# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11415 pmat.rowon_n[2] a_12447_16143# a_14741_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11416 a_30118_56130# pmat.row_n[0] a_30610_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11417 VDD nmat.rowon_n[7] a_38150_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11418 a_47045_33775# a_44763_34293# a_46973_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11419 a_34226_15516# a_18546_15514# a_34134_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1142 a_41254_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11420 VSS pmat.row_n[7] a_20474_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11421 a_50198_23954# a_18162_23548# a_50290_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11422 VSS nmat.sw a_15439_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11423 a_9579_26159# a_9135_26409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X11424 a_3052_29967# a_2051_29973# a_2980_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11425 a_42562_62194# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11426 a_31117_27791# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X11427 a_39154_67174# a_18162_67214# a_39246_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11428 a_11877_58261# a_11711_58261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11429 a_2791_57703# a_5692_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X1143 a_35230_8488# a_18546_8486# a_35138_8894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11430 a_31209_28585# a_13641_23439# a_31103_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11431 a_25494_72234# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11432 a_34134_55126# pmat.en_bit_n[1] a_34626_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11433 a_33519_46831# a_14887_46377# a_33382_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11434 a_2163_61761# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11435 VDD clk_ena a_31235_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11436 a_8441_71677# a_8397_71285# a_8275_71689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11437 a_21082_58138# pmat.row_n[2] a_21574_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11438 a_10509_15279# a_9319_15279# a_10400_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X11439 a_11255_35862# a_11297_36091# a_11255_36189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1144 a_20752_39429# a_20848_39429# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X11440 a_27106_7890# a_18162_7484# a_27198_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11441 vcm a_18162_71230# a_43262_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11442 VSS a_1586_63927# a_12723_64789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11443 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11444 a_21478_11866# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11445 vcm a_18162_11500# a_35230_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11446 a_39939_29967# a_39666_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11447 a_43662_24520# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11448 VSS a_2163_67645# a_2124_67771# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11449 a_7044_61519# a_5081_53135# a_6583_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1145 a_29206_59142# a_18546_59184# a_29114_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11450 VDD pmat.rowon_n[10] a_46182_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11451 a_34530_10862# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11452 a_19509_37479# a_19817_37692# a_13597_37571# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X11453 a_46274_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11454 a_3026_36861# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11455 VSS pmat.row_n[5] a_32522_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11456 a_18597_31599# a_18243_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11457 a_29206_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11458 a_19689_38053# a_19233_38215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11459 vcm a_18162_70226# a_47278_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1146 VSS a_34593_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X11460 nmat.col_n[29] ANTENNA__1395__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11461 VDD nmat.en_C0_n a_20078_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11462 a_44174_20942# pmat.row_n[12] a_44666_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11463 a_51694_72556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11464 a_44174_16926# a_18162_16520# a_44266_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11465 VDD a_2199_13887# a_8175_12533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11466 a_4340_67279# a_4298_67191# a_4037_66933# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X11467 a_19470_63198# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11468 a_22085_42902# a_22449_44219# a_23512_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11469 a_47678_62516# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1147 a_14443_66665# a_13919_65871# a_14371_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11470 VDD pmat.rowon_n[4] a_51202_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11471 vcm a_18162_59182# a_33222_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11472 a_51202_62154# a_18162_62194# a_51294_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11473 VSS a_13091_52047# a_17183_52251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11474 a_16657_42567# a_16745_44581# a_17808_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11475 a_6743_47081# a_4955_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.3505e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X11476 a_34134_72194# a_18162_72234# a_34226_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11477 a_37542_21906# nmat.rowon_n[2] a_37146_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11478 a_15021_31841# a_14803_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X11479 a_33526_16886# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1148 a_30610_19500# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11480 a_18563_27791# a_17845_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11481 a_24186_70186# a_18546_70228# a_24094_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11482 a_6976_32375# a_5179_31591# a_7118_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X11483 a_5093_74575# a_4123_76181# a_4505_74005# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11484 vcm a_18162_22544# a_38242_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11485 a_6681_61839# a_4025_54965# a_6583_61519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X11486 a_21574_20504# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11487 VDD pmat.rowoff_n[15] a_24094_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11488 VDD clk_vcm vcm.sky130_fd_sc_hd__nand2_1_0.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11489 a_21174_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1149 a_4174_46831# a_4128_46983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11490 a_42258_20536# a_18546_20534# a_42166_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11491 a_9405_20291# a_6821_18543# a_9309_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11492 a_24094_64162# a_18162_64202# a_24186_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11493 a_45574_69222# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11494 VSS a_10055_31591# a_17588_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11495 a_19834_34191# a_19657_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11496 a_4737_21561# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11497 a_46884_45743# a_46027_44905# a_46968_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X11498 a_3107_25071# a_2683_22089# a_2744_25223# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11499 a_39647_47679# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X115 a_4487_18365# a_3305_17999# a_4124_18231# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1150 a_5645_12015# a_5579_12394# a_5573_12015# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11500 a_25098_70186# pmat.row_n[14] a_25590_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11501 VDD nmat.rowon_n[9] a_27106_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11502 a_25190_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11503 a_22086_12910# a_18162_12504# a_22178_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11504 VSS a_1642_20871# a_1591_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11505 a_38851_30761# a_17842_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11506 a_18199_31094# nmat.en_bit_n[0] a_17740_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11507 a_45270_61150# a_18546_61192# a_45178_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11508 VSS pmat.row_n[13] a_22482_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11509 a_15181_53135# a_10515_15055# a_14931_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X1151 VDD a_77428_38962# vcm.sky130_fd_sc_hd__buf_4_2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X11510 a_49590_68218# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11511 a_12128_30663# a_10147_29415# a_12270_30838# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X11512 a_16911_52423# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11513 a_3793_22729# a_2603_22357# a_3684_22729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11514 VSS a_2007_25597# a_38249_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11515 a_45663_47081# a_30111_47911# a_45567_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11516 a_3431_57167# a_2419_69455# a_3514_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11517 a_3411_33231# a_2787_33237# a_3303_33609# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11518 a_13443_36919# a_13837_36893# a_13503_36893# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11519 a_35138_11906# a_18162_11500# a_35230_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1152 VSS pmat.row_n[8] a_29510_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11520 a_14071_74879# a_13896_74953# a_14250_74941# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11521 a_9675_10396# a_13795_10687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11522 VDD a_31095_42367# a_30955_42689# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11523 a_22787_42325# a_22963_42657# a_22915_42717# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X11524 a_34828_38341# a_33765_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11525 a_19166_21540# a_18546_21538# a_19074_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11526 a_37238_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11527 a_28602_10464# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11528 VSS pmat.row_n[2] a_43566_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11529 a_40554_55166# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1153 VSS a_19689_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X11530 VDD a_23707_34165# a_14589_35286# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11531 VSS pmat.row_n[12] a_26498_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11532 VSS a_27763_27221# nmat.col[23] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11533 VDD a_20310_28029# a_20164_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=2
X11534 a_42783_31849# a_26479_32117# a_42701_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11535 a_23486_65206# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11536 a_46182_61150# pmat.row_n[5] a_46674_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11537 pmat.col_n[28] a_46934_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11538 a_15737_37479# a_16045_37692# a_14719_37737# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X11539 a_7431_71829# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1154 VDD nmat.rowon_n[13] a_34134_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11540 VDD a_21124_39655# a_21028_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11541 a_9889_10681# a_2021_11043# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11542 a_37923_42359# a_36801_42405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X11543 a_20936_44007# a_19873_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11544 VSS a_6799_75637# a_6649_75983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11545 a_44266_67174# a_18546_67216# a_44174_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11546 a_37146_19938# pmat.row_n[11] a_37638_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11547 a_7164_31421# a_7047_31226# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11548 comp.adc_inverter_1.in clk_comp VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11549 VSS a_2411_33749# a_5865_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1155 a_33526_14878# nmat.rowon_n[9] a_33130_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11550 a_14249_49525# nmat.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11551 a_31412_43439# a_31235_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11552 VDD a_14365_68743# a_12789_68021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X11553 a_20474_58178# pmat.rowon_n[2] a_20078_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11554 a_34530_71230# pmat.rowon_n[15] a_34134_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11555 a_19074_63158# pmat.row_n[7] a_19566_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11556 VDD a_11207_11079# a_11417_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11557 a_18546_60188# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11558 VSS pmat.row_n[3] a_29510_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11559 a_12155_20719# a_11903_20969# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1156 a_27198_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11560 a_23582_61512# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11561 a_14646_37782# a_14600_37607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X11562 a_31214_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11563 a_18162_14512# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11564 a_33526_57174# pmat.rowon_n[1] a_33130_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11565 a_27598_16488# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11566 a_32035_44265# a_30913_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11567 a_21174_8488# a_18546_8486# a_21082_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11568 vcm a_18162_63198# a_45270_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11569 a_45178_67174# pmat.row_n[11] a_45670_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1157 VDD ANTENNA__1183__B1.DIODE a_14747_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X11570 VSS a_5331_28309# a_5265_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11571 a_24214_29967# a_24160_30199# a_24131_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X11572 VDD a_4383_7093# a_8113_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11573 VSS a_45112_47607# a_46383_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X11574 VDD a_4608_41909# a_4518_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.89e+11p ps=1.74e+06u w=420000u l=150000u
X11575 VSS a_41665_46805# a_40949_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11576 VSS a_2839_38101# a_2785_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11577 a_3026_26159# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11578 a_22357_35877# a_21124_36391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11579 a_45574_22910# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1158 a_45805_32661# a_40951_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X11580 a_8287_71311# a_7663_71317# a_8179_71689# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11581 VDD a_5136_19783# a_5087_19319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11582 a_22178_63158# a_18546_63200# a_22086_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11583 VSS a_14647_51701# a_14578_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X11584 VSS a_8031_13353# a_9414_12559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11585 a_22578_67536# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11586 a_39246_18528# a_18546_18526# a_39154_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11587 VSS a_17559_51157# pmat.rowoff_n[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X11588 a_32126_24958# VDD a_32618_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11589 a_22817_41317# a_22361_41479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1159 VSS a_5266_17143# a_5541_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X11590 VSS comp_latch a_10525_12879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11591 a_22086_57134# a_18162_57174# a_22178_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11592 VSS pmat.row_n[9] a_38546_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11593 a_42562_15882# pmat.rowoff_n[7] a_42166_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11594 a_25221_46519# a_14887_46377# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11595 VDD a_3956_72373# a_3894_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11596 a_35138_56130# a_18162_56170# a_35230_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11597 VDD a_4032_26311# a_2191_25045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11598 VSS pmat.row_n[14] a_22482_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11599 a_49590_21906# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X116 vcm a_18162_8488# a_23182_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1160 VSS a_8305_20871# a_11803_20535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11600 a_19166_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11601 a_17021_38053# a_13503_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X11602 vcm a_18162_24552# a_44266_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11603 a_26552_36165# a_25393_35877# a_26515_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X11604 a_2347_45743# a_2093_46070# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11605 VSS a_12263_50959# a_17183_51817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11606 vcm a_18162_56170# a_39246_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11607 VSS VDD a_47582_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11608 VDD a_12789_68021# a_12431_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11609 VSS _1187_.A2 a_82778_4399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1161 VDD config_2_in[8] a_1591_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11610 a_10969_71631# a_10699_72943# a_10751_71543# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11611 a_51598_70226# pmat.rowon_n[14] a_51202_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11612 a_43662_58500# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11613 nmat.rowon_n[4] a_14460_11177# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11614 clk_ena a_82815_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11615 VDD a_2319_67740# a_2250_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X11616 a_39550_13874# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11617 a_10057_19203# a_4976_16091# a_9961_19203# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11618 a_22064_31287# a_20310_28029# a_22206_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X11619 VDD a_11057_35836# a_11469_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X1162 a_8723_67191# a_8491_47911# a_8957_67325# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11620 VSS pmat.row_n[3] a_43566_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11621 a_5179_31591# a_37143_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X11622 a_29536_47753# a_28621_47381# a_29189_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X11623 a_45345_31029# a_45019_38645# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11624 a_6601_34863# a_6557_35105# a_6435_34863# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11625 a_13279_68841# a_12719_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11626 a_29510_24918# VSS a_29114_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11627 a_26102_15922# pmat.row_n[7] a_26594_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11628 VSS pmat.row_n[13] a_26498_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11629 a_21174_24552# a_18546_24550# a_21082_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1163 vcm a_18162_65206# a_34226_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11630 a_41558_62194# pmat.rowon_n[6] a_41162_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11631 a_20170_66170# a_18546_66212# a_20078_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11632 a_30610_13476# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11633 a_29606_57496# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11634 VDD nmat.rowon_n[7] a_14460_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X11635 VSS a_2847_36799# a_2781_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X11636 a_23345_47741# a_23301_47349# a_23179_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11637 VDD VSS a_33130_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11638 a_34924_37253# a_33765_36965# a_34887_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X11639 a_3262_72399# a_3136_72515# a_2858_72531# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1164 a_38546_66210# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11640 a_34226_23548# a_18546_23546# a_34134_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11641 VDD pmat.rowon_n[2] a_20078_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11642 VSS pmat.row_n[1] a_40554_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11643 a_38150_8894# pmat.row_n[0] a_38642_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11644 a_19470_16886# nmat.rowon_n[7] a_19074_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11645 a_46513_39009# a_40837_46261# a_46427_39009# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X11646 VDD a_33567_30199# a_32865_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X11647 a_20474_11866# nmat.rowon_n[12] a_20078_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11648 VSS pmat.row_n[4] a_29510_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11649 a_38546_60186# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1165 a_34134_69182# pmat.row_n[13] a_34626_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11650 a_50594_9858# nmat.rowon_n[14] a_50198_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11651 a_14646_37455# a_14600_37607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11652 a_38546_19898# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11653 pmat.col_n[16] a_26891_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.1125e+11p pd=1.95e+06u as=0p ps=0u w=650000u l=150000u
X11654 a_33526_10862# nmat.rowon_n[13] a_33130_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11655 VDD a_13529_34951# a_14864_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11656 a_40158_70186# a_18162_70226# a_40250_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11657 vcm a_18162_62194# a_21174_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11658 VDD a_23700_39655# a_23604_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11659 a_21082_66170# pmat.row_n[10] a_21574_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1166 a_12969_40175# a_12543_40214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11660 a_26423_40183# a_25301_40229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X11661 a_10209_22351# a_6664_26159# a_10137_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X11662 vcm a_18162_61190# a_34226_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11663 a_8727_70197# a_1674_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X11664 a_39646_22512# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11665 VDD pmat.rowoff_n[12] a_43170_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11666 a_30913_38779# a_29864_39429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11667 a_7275_51727# a_6651_51733# a_7167_52105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11668 a_46274_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11669 a_43170_61150# a_18162_61190# a_43262_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1167 a_45574_67214# pmat.rowon_n[11] a_45178_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11670 VDD a_17478_46805# a_12079_9615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11671 VDD a_2791_57703# a_4135_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X11672 a_12323_58633# a_11877_58261# a_12227_58633# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11673 a_26276_39429# a_25117_39141# a_26180_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11674 a_32522_58178# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11675 a_46578_71230# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11676 a_3993_44431# a_2659_35015# a_3911_44431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11677 a_10054_57961# a_7521_47081# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11678 vcm a_18162_68218# a_20170_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11679 a_44174_24958# a_18162_24552# a_44266_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1168 VSS pmat.row_n[8] a_42562_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11680 a_47678_70548# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11681 a_31220_47919# a_31152_48071# a_30947_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=3.4735e+11p ps=3.68e+06u w=650000u l=150000u
X11682 VSS a_10985_42044# a_10677_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11683 a_44266_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11684 vcm a_18162_67214# a_33222_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11685 VDD a_15021_31841# a_14911_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11686 a_47186_60146# a_18162_60186# a_47278_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11687 VSS pmat.row_n[5] a_40554_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11688 a_22915_42717# a_10949_43124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11689 a_4220_62037# a_4520_60975# a_4349_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X1169 a_4859_31274# a_4951_31029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11690 a_10449_60975# a_10286_60405# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11691 VSS a_14645_28381# a_14751_28341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11692 a_20170_11500# a_18546_11498# a_20078_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11693 a_23582_8456# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11694 VSS pmat.row_n[15] a_23486_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11695 VDD nmat.rowon_n[12] a_37146_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11696 vcm a_18162_12504# a_29206_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11697 a_21174_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11698 VSS a_22541_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X11699 a_33222_10496# a_18546_10494# a_33130_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X117 VDD a_17306_28879# a_17748_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X1170 VSS a_5749_57685# a_5683_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11700 VDD nmat.rowon_n[15] a_33130_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11701 vcm a_18162_59182# a_41254_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11702 VDD a_12447_16143# a_14287_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11703 a_9551_31094# a_4259_31375# a_9092_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11704 a_24186_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11705 a_48586_68218# pmat.rowon_n[12] a_48190_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11706 a_22925_28111# ANTENNA__1395__A2.DIODE nmat.col_n[2] VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11707 a_7197_42479# a_6007_42479# a_7088_42479# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11708 a_41558_16886# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11709 a_28705_39141# a_28116_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1171 VDD a_44849_45717# a_44879_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11710 a_2107_26159# a_1591_26159# a_2012_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X11711 a_22086_20942# a_18162_20536# a_22178_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11712 a_25190_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11713 a_11415_14557# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11714 a_2781_43401# a_1591_43029# a_2672_43401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11715 a_11115_71285# a_11203_62037# a_10975_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X11716 a_10541_8573# a_10378_7637# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11717 VSS a_14887_46377# a_34850_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11718 a_2882_61519# a_2124_61635# a_2319_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11719 a_9092_31287# a_4259_31375# a_9234_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1172 a_12437_28585# a_12155_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11720 VSS a_15667_27239# a_45832_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11721 vcm a_18162_18528# a_28202_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11722 a_14725_26703# a_8861_24527# a_14607_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=3.04e+06u as=0p ps=0u w=1e+06u l=150000u
X11723 VDD pmat.rowon_n[5] a_45178_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11724 a_27049_35515# a_26552_36165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11725 a_32218_16520# a_18546_16518# a_32126_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11726 a_4135_37815# a_3325_36495# a_4309_37921# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11727 VDD a_7111_74575# a_2149_45717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X11728 a_43349_47081# a_35186_47375# a_43267_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11729 a_27502_17890# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1173 a_43170_65166# a_18162_65206# a_43262_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11730 VDD nmat.rowon_n[4] a_36142_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11731 VSS pmat.row_n[7] a_31518_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11732 a_34705_51959# a_30663_50087# a_41422_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X11733 a_40554_63198# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11734 a_2163_55233# a_1586_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11735 a_46723_30485# a_35244_32411# a_46921_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X11736 a_37146_68178# a_18162_68218# a_37238_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11737 vcm a_18162_8488# a_44266_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11738 VSS a_1586_18231# a_5087_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11739 VDD vcm.sky130_fd_sc_hd__buf_4_3.A a_77980_38962# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1174 VDD a_7436_16519# a_7387_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11740 a_12002_49917# a_11948_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11741 VSS a_2847_26133# a_2781_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11742 VDD pmat.rowon_n[4] a_49194_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11743 a_32126_58138# pmat.row_n[2] a_32618_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11744 a_22684_40743# a_21621_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11745 a_23420_36165# a_22357_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11746 a_32522_11866# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11747 a_29114_10902# a_18162_10496# a_29206_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11748 a_45943_47375# a_33467_46261# a_45450_48695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11749 a_19074_71190# pmat.row_n[15] a_19566_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1175 a_21239_47349# a_21215_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X11750 a_2369_16189# a_2325_15797# a_2203_16201# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11751 a_44266_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11752 a_20170_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11753 a_10747_6727# a_10378_7637# a_11145_6575# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11754 a_27198_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11755 a_14734_64015# pmat.rowon_n[7] a_14565_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X11756 a_11112_77661# a_10898_77661# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11757 a_44570_64202# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11758 VDD a_43533_30761# a_47035_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X11759 a_7479_22467# a_6817_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X1176 a_9084_51843# a_8385_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11760 a_42166_21946# pmat.row_n[13] a_42658_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11761 a_42166_17930# a_18162_17524# a_42258_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11762 VSS _1192_.A2 a_46481_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X11763 a_11421_17455# a_10995_17782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11764 VSS comp.adc_nor_latch_0.NOR_1/A comp.adc_nor_latch_0.QN VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11765 VDD VSS a_31122_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11766 a_6643_5724# a_6448_5755# a_6953_5487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X11767 VDD a_20221_40835# a_34828_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11768 a_2275_46070# a_2093_46070# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11769 a_1846_69931# a_2124_69947# a_2080_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1177 VSS a_44774_40821# a_45246_41167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X11770 a_35630_16488# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11771 a_36453_29199# a_31263_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11772 VDD cgen.dlycontrol4_in[1] a_1945_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11773 VDD a_38727_32447# a_38714_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11774 a_24490_67214# pmat.rowon_n[11] a_24094_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11775 VSS pmat.row_n[8] a_21478_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11776 a_6643_5724# a_6487_5629# a_6788_5853# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X11777 vcm a_18162_15516# a_31214_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11778 a_48682_15484# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11779 a_48586_21906# nmat.rowon_n[2] a_48190_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1178 a_35534_59182# pmat.rowon_n[3] a_35138_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11780 a_45178_12910# pmat.row_n[4] a_45670_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11781 a_24847_38543# a_12513_39100# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11782 VDD a_24833_34191# a_27579_34967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11783 a_2215_23439# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11784 a_36946_34191# a_36769_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11785 a_22086_65166# a_18162_65206# a_22178_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11786 a_28110_22950# pmat.row_n[14] a_28602_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11787 VSS a_6087_70919# a_4396_69109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X11788 a_32618_20504# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11789 VDD a_4048_74549# a_3986_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1179 a_4491_53511# a_4243_54991# a_4725_53359# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11790 a_32218_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11791 a_35138_64162# a_18162_64202# a_35230_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11792 a_38546_13874# nmat.rowon_n[10] a_38150_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11793 VDD a_6579_21583# a_6981_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11794 VSS a_20221_40835# a_34887_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11795 cgen.dlycontrol1_in[0] a_1591_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11796 a_43359_29967# a_41227_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11797 vcm a_18162_7484# a_33222_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11798 a_19074_18934# a_18162_18528# a_19166_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11799 VDD pmat.rowoff_n[7] a_25098_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X118 a_20175_49667# a_19283_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X1180 a_18162_12504# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11800 a_22578_12472# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11801 vcm a_18162_64202# a_39246_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11802 a_49194_11906# pmat.row_n[3] a_49686_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11803 a_37813_39867# a_36227_38771# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X11804 a_39154_68178# pmat.row_n[12] a_39646_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11805 a_20078_13914# a_18162_13508# a_20170_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11806 a_43262_62154# a_18546_62196# a_43170_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11807 a_4307_35639# a_2563_34837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11808 a_43662_66532# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11809 a_18176_35077# a_17113_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1181 VDD a_22064_31287# a_20895_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11810 a_40158_63158# pmat.row_n[7] a_40650_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11811 a_30140_43781# a_28981_43493# a_30103_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X11812 a_33130_12910# a_18162_12504# a_33222_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11813 a_82925_25615# _1192_.A2 nmat.col[26] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11814 a_9581_73487# a_9103_73791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11815 a_1644_59861# a_1591_58799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11816 VSS a_30111_47911# a_32507_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X11817 a_30663_50087# a_45107_34863# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11818 a_14839_54599# a_14655_53359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11819 VDD a_13805_43990# a_15048_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X1182 VSS a_19551_34191# a_19657_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11820 a_26102_66170# a_18162_66210# a_26194_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11821 a_26594_11468# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11822 a_6631_42845# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11823 a_9004_47741# a_8453_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11824 a_2250_65693# a_2124_65595# a_1846_65579# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11825 VSS a_13275_48783# a_13688_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11826 VDD pmat.rowon_n[10] a_20078_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11827 a_44174_62154# pmat.row_n[6] a_44666_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11828 a_14885_52093# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11829 a_6179_69831# a_2879_57487# a_6524_69679# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X1183 a_44791_43541# a_31675_47695# a_45222_43567# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X11830 a_30118_9898# pmat.row_n[1] a_30610_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11831 VSS a_36161_37462# a_37463_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11832 a_10597_24233# a_10513_24135# a_10515_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11833 ANTENNA__1195__A1.DIODE a_46487_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11834 a_20170_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11835 a_42258_68178# a_18546_68220# a_42166_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11836 a_14504_37607# a_14719_37737# a_14646_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X11837 vcm a_18162_70226# a_21174_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11838 VDD a_7571_32687# a_5363_33551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11839 a_7589_33749# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1184 a_23007_41807# a_10949_42364# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X11840 a_2242_44150# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X11841 a_48190_19938# pmat.row_n[11] a_48682_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11842 a_5871_32362# a_5963_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11843 VDD pmat.rowon_n[9] a_24094_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11844 a_21574_62516# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11845 a_38242_13508# a_18546_13506# a_38150_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11846 a_31518_58178# pmat.rowon_n[2] a_31122_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11847 VDD a_19439_50095# a_16083_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11848 a_45574_71230# pmat.rowon_n[15] a_45178_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11849 a_12889_64789# a_12723_64789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1185 vcm a_18162_17524# a_25190_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11850 vcm.sky130_fd_sc_hd__buf_4_3.X a_77980_38962# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11851 a_10953_43781# a_11261_43421# a_10927_43421# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X11852 a_34626_61512# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11853 cgen.dlycontrol4_in[4] a_2235_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11854 VSS a_6699_76983# a_5047_76983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11855 a_10586_24643# a_5351_19913# a_10513_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X11856 a_46182_8894# pmat.row_n[0] a_46674_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11857 a_24490_20902# pmat.rowoff_n[12] a_24094_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11858 VDD pmat.rowon_n[0] a_27106_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11859 a_12543_39126# a_12513_39100# a_12471_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X1186 a_2781_20553# a_1591_20181# a_2672_20553# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11860 a_49590_70226# pmat.rowon_n[14] a_49194_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11861 a_43566_23914# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11862 a_18546_57176# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11863 pmat.col[30] a_24867_53135# a_47858_53135# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11864 a_50690_18496# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11865 VSS a_4267_35407# a_4601_35727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11866 a_37238_19532# a_18546_19530# a_37146_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11867 a_44266_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11868 VDD a_41475_31751# a_41427_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11869 VDD a_5579_12394# a_5417_11445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X1187 a_6447_40669# a_5823_40303# a_6339_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X11870 VSS a_7797_63151# a_9414_63695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11871 a_20078_58138# a_18162_58178# a_20170_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11872 a_39550_62194# pmat.rowon_n[6] a_39154_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11873 VSS pmat.row_n[10] a_36538_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11874 a_40554_16886# nmat.rowon_n[7] a_40158_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11875 a_13327_70741# a_14439_72703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11876 vcm a_18162_20536# a_29206_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11877 a_33130_57134# a_18162_57174# a_33222_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11878 a_12038_55687# a_10497_54697# a_12252_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=0p ps=0u w=1e+06u l=150000u
X11879 VSS pmat.row_n[9] a_49590_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1188 a_2375_18708# a_2467_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11880 a_20078_17930# pmat.row_n[9] a_20570_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11881 a_3569_59709# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11882 VDD a_2319_31836# a_2250_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X11883 vcm a_18162_67214# a_41254_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11884 VDD config_1_in[2] a_1591_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11885 VDD a_7079_34837# a_6559_33767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X11886 vcm a_18162_57174# a_37238_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11887 a_2107_18377# a_1757_18005# a_2012_18365# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X11888 a_26141_49871# a_25802_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11889 a_9287_77055# a_9112_77129# a_9466_77117# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1189 VDD pmat.rowoff_n[7] a_46182_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11890 a_41254_55126# a_18546_55168# a_41162_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11891 a_6882_49373# a_5805_49007# a_6720_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11892 a_41654_59504# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11893 a_9655_74216# a_9831_74183# a_10041_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11894 a_37542_14878# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11895 a_18546_22542# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11896 a_25384_46403# a_14887_46377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11897 a_22186_30485# a_22628_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11898 a_9666_32275# a_9983_32385# a_9941_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11899 a_37638_7452# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X119 VDD a_2263_43719# a_3891_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1190 VSS a_28812_29575# a_29455_31293# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X11900 a_26498_59182# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11901 VDD ANTENNA__1395__A1.DIODE a_25691_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X11902 a_12693_38543# a_12267_38870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11903 pmat.rowon_n[10] nmat.rowon_n[7] a_14471_62063# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11904 VDD a_5688_52423# a_4659_53738# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X11905 a_26498_17890# nmat.rowon_n[6] a_26102_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11906 VSS a_28061_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X11907 VSS pmat.row_n[1] a_30514_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11908 VDD a_19487_53034# pmat.rowoff_n[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11909 a_24094_16926# pmat.row_n[8] a_24586_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1191 a_11113_40835# a_36617_42043# a_37739_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X11910 a_2215_50461# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11911 a_44665_45519# a_43720_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11912 VSS a_2319_74268# a_2250_74397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11913 a_12709_54223# a_9581_56079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11914 a_2250_52815# a_2124_52931# a_1846_52947# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11915 a_13278_51549# a_12559_51325# a_12715_51420# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X11916 a_32514_50141# a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11917 a_32218_24552# a_18546_24550# a_32126_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11918 a_31214_66170# a_18546_66212# a_31122_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11919 VSS a_31097_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X1192 a_23821_35279# a_23655_35279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11920 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11921 a_12449_39605# a_12116_39783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11922 a_27198_56130# a_18546_56172# a_27106_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11923 a_4985_51433# a_2983_48071# a_4903_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11924 VDD ANTENNA__1183__B1.DIODE a_14565_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X11925 VSS VDD a_19470_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11926 a_35138_7890# VDD a_35630_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11927 a_2007_8916# a_2099_8725# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11928 VDD pmat.rowon_n[2] a_31122_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11929 VSS a_25301_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X1193 clk_ena a_82815_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11930 VSS pmat.row_n[5] a_27502_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11931 VSS a_6200_70919# a_11530_77661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11932 VDD a_18563_27791# a_41237_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11933 a_31518_11866# nmat.rowon_n[12] a_31122_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11934 a_14641_57167# a_14287_57280# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11935 vcm a_18162_18528# a_36234_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11936 VDD a_45253_27221# nmat.col[25] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11937 a_40250_16520# a_18546_16518# a_40158_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11938 a_11041_40948# a_11071_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11939 a_18162_61190# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X1194 pmat.row_n[10] a_21239_50613# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X11940 vcm a_18162_62194# a_32218_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11941 a_11793_27907# a_9741_28585# a_11711_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11942 VDD cgen.enable_dlycontrol_in a_24667_40719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11943 VSS pmat.row_n[10] a_39550_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11944 a_11711_27907# a_9741_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X11945 a_12253_10927# comp_latch a_11207_11079# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11946 a_41254_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11947 a_32126_66170# pmat.row_n[10] a_32618_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11948 VDD a_12967_58559# a_12954_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11949 vcm a_18162_17524# a_49286_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1195 a_20083_51843# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11950 VDD a_11067_27239# a_26234_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X11951 a_39469_39141# a_38972_39655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X11952 a_3445_66237# a_3410_66003# a_3207_65845# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11953 a_43566_64202# pmat.rowon_n[8] a_43170_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11954 a_19487_53034# a_19579_52789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11955 a_37638_23516# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11956 vcm a_18162_12504# a_50290_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11957 a_37238_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11958 VDD nmat.rowon_n[2] a_41162_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11959 a_29698_47375# a_28621_47381# a_29536_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1196 a_35068_46805# a_35186_47375# a_35390_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11960 a_6631_42845# a_6007_42479# a_6523_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11961 a_44266_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11962 VDD a_9827_8181# a_9766_8207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X11963 a_2672_16201# a_1757_15829# a_2325_15797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X11964 VDD a_8851_12533# a_8782_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11965 a_12267_38870# a_12309_38659# a_12267_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11966 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11967 a_13529_43781# a_13837_43421# a_13503_43421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X11968 a_27398_47197# a_26321_46831# a_27236_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X11969 a_44570_72234# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1197 a_39550_58178# pmat.rowon_n[2] a_39154_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11970 VSS a_12107_62037# a_11883_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X11971 VDD VDD a_22086_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11972 a_26194_17524# a_18546_17522# a_26102_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11973 a_38150_15922# a_18162_15516# a_38242_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11974 a_25393_38053# a_23700_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X11975 a_3883_65845# a_3688_65987# a_4193_66237# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X11976 a_4033_56417# a_3967_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11977 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11978 a_42258_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11979 VDD a_82971_11989# nmat.col_n[28] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u M=2
X1198 VSS pmat.en_bit_n[0] a_36538_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u M=2
X11980 VDD a_3923_68021# a_3881_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11981 a_34924_36165# a_33765_35877# a_34887_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X11982 VSS a_12447_16143# a_14011_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11983 a_7033_51433# a_6979_51157# a_6835_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11984 a_26102_57134# pmat.row_n[1] a_26594_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11985 VDD a_39647_48767# a_39634_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11986 a_35230_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11987 a_37542_55166# VSS a_37146_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11988 VSS VDD a_21478_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11989 a_30610_55488# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1199 a_31539_51946# a_31631_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11990 a_3325_20175# a_2847_20479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11991 vcm a_18162_23548# a_31214_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11992 a_22743_35561# a_21621_35515# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11993 a_7895_60214# a_6175_60039# a_7436_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11994 VSS pmat.row_n[5] a_51598_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11995 vcm a_18162_13508# a_27198_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11996 a_48282_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11997 a_3029_69135# a_3069_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11998 a_4699_13647# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11999 VSS pmat.row_n[15] a_34530_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VSS pmat.row_n[1] a_47582_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X120 a_21574_13476# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1200 a_2129_12559# a_1959_12559# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12000 a_31214_11500# a_18546_11498# a_31122_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12001 VDD nmat.rowon_n[12] a_48190_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12002 VDD a_2007_25597# a_35039_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12003 VDD pmat.rowon_n[12] a_38150_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12004 a_5046_67655# a_5307_67655# a_5260_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X12005 a_26498_12870# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12006 a_32218_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12007 VSS pmat.row_n[2] a_30514_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12008 a_33223_42359# a_33617_42333# a_33283_42333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X12009 VDD a_12531_42583# a_12344_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1201 a_20474_72234# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12010 a_20078_7890# a_18162_7484# a_20170_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12011 a_2781_36873# a_1591_36501# a_2672_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X12012 vcm a_18162_72234# a_39246_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12013 a_43262_70186# a_18546_70228# a_43170_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12014 VSS a_1923_31743# a_2369_23805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12015 a_50198_10902# a_18162_10496# a_50290_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12016 a_36142_22950# pmat.row_n[14] a_36634_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12017 a_40158_71190# pmat.row_n[15] a_40650_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12018 a_39246_60146# a_18546_60188# a_39154_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12019 a_29163_29423# a_28626_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=150000u
X1202 VSS a_30913_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X12020 a_40650_20504# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12021 a_39646_64524# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12022 VDD a_1923_53055# a_2195_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12023 a_20776_51959# a_18547_51565# a_21007_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12024 a_40250_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12025 a_43262_7484# a_18546_7482# a_43170_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12026 a_33130_20942# a_18162_20536# a_33222_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12027 VDD pmat.rowon_n[6] a_43170_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12028 a_9457_51163# a_8385_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12029 a_2629_71855# a_2250_72221# a_2557_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1203 a_23788_40517# a_22725_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X12030 VSS pmat.row_n[6] a_28506_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12031 a_2834_8207# a_1757_8213# a_2672_8585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12032 a_25494_18894# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12033 a_30210_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12034 a_32522_60186# pmat.rowon_n[4] a_32126_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12035 a_32522_19898# nmat.rowon_n[4] a_32126_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12036 a_46817_43541# a_46950_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X12037 a_22297_46653# a_15899_47939# a_22225_46653# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12038 vcm a_18162_9492# a_24186_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12039 a_44174_70186# pmat.row_n[14] a_44666_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1204 VSS a_22357_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X12040 a_29206_71190# a_18546_71232# a_29114_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12041 VDD a_3797_14709# a_3687_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12042 a_41162_12910# a_18162_12504# a_41254_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12043 a_48190_68178# a_18162_68218# a_48282_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12044 a_20170_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12045 VDD VSS a_29114_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12046 VSS pmat.row_n[13] a_41558_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12047 a_11603_28335# a_11159_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X12048 a_33222_58138# a_18546_58180# a_33130_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12049 vcm a_18162_55166# a_30210_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1205 VSS pmat.row_n[9] a_19470_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12050 a_34226_9492# a_18546_9490# a_34134_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12051 a_4441_74031# a_4409_74183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12052 a_30118_59142# pmat.row_n[3] a_30610_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12053 a_43548_30287# a_28704_29568# a_43359_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12054 a_33957_48437# a_30111_47911# a_36178_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12055 a_40650_9460# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12056 VSS a_3325_20175# a_8256_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12057 a_38242_21540# a_18546_21538# a_38150_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12058 a_35186_47375# a_33986_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12059 a_21574_70548# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1206 a_50594_61190# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12060 a_42258_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12061 a_2325_50337# a_2107_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X12062 VDD nmat.rowon_n[14] a_50198_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12063 a_47011_31029# a_47685_30517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12064 a_21082_60146# a_18162_60186# a_21174_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12065 VSS pmat.row_n[12] a_45574_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12066 a_42562_65206# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12067 a_32030_48169# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12068 VDD a_7521_47081# a_9871_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12069 a_42658_17492# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1207 a_3704_58575# a_2419_53351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12070 a_31214_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12071 a_14335_23439# a_14371_25071# a_13977_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12072 a_5411_12167# a_4865_12533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12073 a_40158_18934# a_18162_18528# a_40250_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12074 VDD config_2_in[7] a_1591_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12075 a_2463_44477# a_2315_44124# a_2100_44343# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12076 VDD a_4036_70741# a_3710_70455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12077 VDD a_10190_60663# a_10191_57691# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12078 VSS a_45921_42167# a_44966_43255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12079 a_11041_38772# a_11347_36950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1208 vcm a_18162_16520# a_29206_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12080 VDD nmat.rowon_n[13] a_24094_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12081 VSS a_4503_70455# a_4421_70741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12082 a_10959_23983# a_10515_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X12083 a_36341_38053# a_34924_37253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X12084 a_1644_54421# a_1591_54991# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12085 a_22482_68218# pmat.rowon_n[12] a_22086_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12086 VSS pmat.row_n[3] a_48586_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12087 VSS a_3325_26159# a_3891_25623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12088 a_45574_56170# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12089 a_13317_10749# a_13273_10357# a_13151_10761# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1209 a_4583_68021# a_7674_69135# a_8538_69455# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X12090 VSS a_26497_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X12091 a_50290_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12092 a_36234_69182# a_18546_69224# a_36142_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12093 a_46674_16488# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12094 a_43170_13914# pmat.row_n[5] a_43662_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12095 a_28506_66210# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12096 a_14460_61225# nmat.rowon_n[7] a_14287_60975# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X12097 VSS a_13837_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X12098 VSS pmat.row_n[8] a_32522_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12099 a_23847_38007# a_22725_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X121 VSS pmat.row_n[2] a_47582_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1210 a_47186_66170# a_18162_66210# a_47278_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12100 a_7618_15645# a_6541_15279# a_7456_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12101 a_55914_40254# comp.adc_nor_latch_0.NOR_1/A comp.adc_nor_latch_0.QN VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=4.96e+11p ps=4.44e+06u w=800000u l=150000u
X12102 a_45625_36495# a_35244_32411# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X12103 a_4737_21561# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12104 a_6179_69831# a_5081_53135# a_6346_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X12105 a_14642_23983# a_11337_25071# a_14475_24233# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12106 a_33130_65166# a_18162_65206# a_33222_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12107 a_36538_14878# nmat.rowon_n[9] a_36142_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12108 a_17159_47919# a_10055_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X12109 a_25494_59182# pmat.rowon_n[3] a_25098_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1211 a_9287_65087# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12110 VSS pmat.row_n[0] a_22482_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12111 a_19566_18496# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12112 a_11497_38543# a_11071_38870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12113 a_49590_55166# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12114 a_7206_5853# a_6448_5755# a_6643_5724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12115 a_14737_53359# a_14653_53458# a_14655_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12116 VDD nmat.rowon_n[7] a_23090_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12117 vcm a_18162_65206# a_37238_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12118 a_24094_9898# a_18162_9492# a_24186_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12119 a_37146_69182# pmat.row_n[13] a_37638_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1212 a_33222_14512# a_18546_14510# a_33130_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12120 a_41254_63158# a_18546_63200# a_41162_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12121 VDD a_19615_41959# a_19428_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12122 a_41654_67536# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12123 a_2871_51701# a_2676_51843# a_3181_52093# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X12124 a_4984_41935# a_4149_41941# a_5012_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12125 VSS a_2411_33749# a_6877_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12126 VDD a_6795_76989# a_9183_76359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12127 a_51202_24958# VDD a_51694_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12128 a_18429_51189# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12129 a_34226_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1213 a_33526_71230# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12130 a_13985_44581# a_12292_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12131 a_41162_57134# a_18162_57174# a_41254_57134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X12132 VSS a_12197_43746# a_11261_43421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X12133 VSS a_7899_67477# a_7845_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12134 a_10095_16950# a_9913_16950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12135 a_6817_21583# a_3305_17999# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12136 a_24094_67174# a_18162_67214# a_24186_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12137 a_29510_58178# pmat.rowon_n[2] a_29114_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12138 VSS VDD a_26498_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12139 a_2250_59165# a_2124_59067# a_1846_59051# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1214 vcm a_18162_11500# a_30210_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12140 VSS pmat.row_n[14] a_41558_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12141 VSS a_45019_38645# a_44515_38645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12142 a_38242_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12143 a_9995_52299# a_4259_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12144 a_8749_47381# a_8583_47381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12145 a_1757_40853# a_1591_40853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12146 a_2100_44343# a_2315_44124# a_2242_44150# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X12147 a_30095_36919# a_30489_36893# a_30155_36893# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X12148 a_27198_64162# a_18546_64204# a_27106_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12149 VDD a_76962_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_3.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1215 a_37238_64162# a_18546_64204# a_37146_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12150 a_9889_10681# a_2021_11043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12151 a_27598_68540# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12152 VDD pmat.rowon_n[10] a_31122_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12153 a_34530_17890# nmat.rowon_n[6] a_34134_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12154 a_2217_29973# a_2051_29973# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12155 VSS a_2659_35015# a_6559_44431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12156 a_31214_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12157 VDD a_21239_50613# pmat.row_n[10] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X12158 VSS pmat.row_n[13] a_45574_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12159 VDD a_1925_20871# a_1738_20693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1216 a_47678_11468# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12160 VSS a_5768_9527# a_5738_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.64e+11p ps=3.72e+06u w=650000u l=150000u M=2
X12161 a_45670_7452# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12162 a_41558_7850# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12163 a_40250_24552# a_18546_24550# a_40158_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12164 VDD a_4516_21531# a_6997_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12165 a_21867_34709# a_12513_36924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12166 a_11071_38870# a_11113_38659# a_11071_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12167 a_48682_57496# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12168 ANTENNA__1190__B1.DIODE a_47039_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=8
X12169 vcm a_18162_70226# a_32218_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1217 a_24186_7484# a_18546_7482# a_24094_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12170 a_36234_14512# a_18546_14510# a_36142_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12171 a_35230_56130# a_18546_56172# a_35138_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12172 vcm a_18162_60186# a_28202_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12173 a_43566_72234# VDD a_43170_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12174 a_6835_51183# a_6883_51335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12175 VDD a_13357_37429# a_13301_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X12176 a_28110_64162# pmat.row_n[8] a_28602_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12177 vcm a_18162_20536# a_50290_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12178 a_49286_13508# a_18546_13506# a_49194_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12179 a_32618_62516# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1218 a_37638_68540# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12180 VSS pmat.row_n[5] a_35534_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12181 a_24565_34789# a_23700_36391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12182 a_22206_31421# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12183 VSS pmat.row_n[4] a_48586_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12184 a_22482_21906# nmat.rowon_n[2] a_22086_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12185 a_27785_43131# a_27329_42902# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12186 VDD a_2672_26159# a_2847_26133# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12187 VDD pmat.rowon_n[1] a_25098_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12188 VDD a_35068_46805# a_12263_50959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u M=2
X12189 vcm a_18162_22544# a_23182_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1219 _1184_.A2 a_44888_33205# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12190 VSS a_19459_35279# a_19565_35279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12191 a_32522_9858# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12192 VDD a_1957_43567# a_11807_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12193 a_4222_33597# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12194 VSS a_9643_66389# a_9552_67191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X12195 VSS cgen.enable_dlycontrol_in a_21815_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12196 a_38150_23954# a_18162_23548# a_38242_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12197 a_30514_69222# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12198 a_25494_12870# pmat.rowoff_n[4] a_25098_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12199 a_37542_63198# pmat.rowon_n[7] a_37146_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X122 VDD nmat.rowon_n[7] a_24094_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1220 a_6343_32661# a_6168_32687# a_6522_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12200 a_2375_16532# a_2467_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12201 a_13593_74941# a_13549_74549# a_13427_74953# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12202 vcm a_18162_21540# a_27198_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12203 a_45178_71190# a_18162_71230# a_45270_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12204 a_51598_58178# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12205 VSS pmat.row_n[10] a_47582_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12206 a_12292_44869# a_11133_44581# a_12255_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12207 a_30210_61150# a_18546_61192# a_30118_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12208 a_51598_16886# nmat.rowon_n[7] a_51202_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12209 a_39949_50959# ANTENNA__1190__A1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1221 VDD pmat.rowon_n[10] a_41162_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12210 a_34530_68218# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12211 pmat.rowoff_n[11] a_14460_60137# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X12212 a_6170_5739# a_6487_5629# a_6445_5487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X12213 VDD nmat.rowon_n[1] a_35138_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12214 a_25794_49007# a_25802_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12215 VDD pmat.rowon_n[2] a_29114_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12216 a_29114_7890# a_18162_7484# a_29206_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12217 a_10329_30753# a_10111_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12218 a_2129_10383# a_1959_10383# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12219 a_29510_11866# nmat.rowon_n[12] a_29114_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1222 VSS a_23395_53135# a_26695_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X12220 a_20605_40719# a_20179_41046# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12221 vcm a_18162_57174# a_48282_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12222 a_18568_51959# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12223 a_22178_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12224 a_49194_70186# a_18162_70226# a_49286_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12225 a_48586_14878# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12226 VDD a_17635_39605# a_17441_40482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12227 a_5085_59343# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12228 VDD a_25802_48169# a_25893_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12229 a_10233_7913# a_10047_8751# a_9827_8181# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1223 a_31425_37218# a_30913_36603# a_32035_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X12230 a_39646_72556# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12231 a_31122_61150# pmat.row_n[5] a_31614_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12232 a_40250_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12233 a_8325_10901# a_1717_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12234 nmat.col[1] a_10883_3303# a_13565_3087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12235 VSS a_10873_39605# a_25815_43957# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12236 VDD nmat.rowon_n[2] a_39154_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12237 a_24861_29423# a_8583_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12238 VSS a_37960_42693# a_37923_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12239 VDD pmat.rowon_n[14] a_43170_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1224 a_9651_69679# a_9301_69679# a_9556_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X12240 vcm a_18162_69222# a_25190_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12241 a_35138_16926# pmat.row_n[8] a_35630_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12242 a_36234_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12243 a_5271_14557# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12244 a_39154_62154# a_18162_62194# a_39246_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12245 a_13025_51183# a_12646_51549# a_12953_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12246 a_7160_33927# a_6559_33767# a_7302_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12247 a_22086_19938# pmat.row_n[11] a_22578_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12248 VSS a_2046_30184# a_6743_31061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12249 a_43262_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1225 a_46449_46261# a_46582_46519# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X12250 VSS a_30913_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X12251 a_28981_43493# a_28525_43655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12252 a_10789_6575# a_10747_6727# a_9459_5461# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X12253 VDD a_37820_30485# a_45212_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12254 a_26194_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12255 a_7799_58621# a_4843_54826# a_7436_58487# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12256 ANTENNA__1197__A.DIODE a_47407_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X12257 a_9098_71677# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12258 a_25190_12504# a_18546_12502# a_25098_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12259 a_9135_22057# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1226 a_18277_37620# ndecision_finish VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12260 VSS a_13357_37429# a_13301_37782# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12261 a_41162_20942# a_18162_20536# a_41254_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12262 vcm a_18162_68218# a_29206_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12263 a_11113_36483# a_19689_34789# a_20811_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12264 a_11285_39958# a_11113_39747# a_11071_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X12265 VSS pmat.row_n[11] a_37542_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12266 vcm a_18162_63198# a_30210_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12267 vcm a_18162_18528# a_47278_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12268 a_30118_67174# pmat.row_n[11] a_30610_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12269 a_41558_65206# pmat.rowon_n[9] a_41162_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1227 a_21215_48071# a_28629_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.8675e+11p pd=3.79e+06u as=0p ps=0u w=650000u l=150000u M=2
X12270 a_51294_16520# a_18546_16518# a_51202_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12271 VDD ANTENNA__1190__A1.DIODE a_44183_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X12272 a_29206_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12273 a_46578_17890# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12274 VSS pmat.row_n[7] a_50594_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12275 VSS a_11057_35836# a_11476_36189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12276 vcm a_18162_8488# a_38242_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12277 a_38205_32117# a_37987_32521# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12278 a_30514_22910# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12279 a_27106_21946# a_18162_21540# a_27198_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1228 a_41254_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12280 VDD a_6927_30503# a_12453_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X12281 VDD pmat.rowon_n[7] a_37146_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12282 a_24186_18528# a_18546_18526# a_24094_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12283 a_12294_22467# a_5899_21807# a_12212_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12284 a_16745_34427# a_15144_35077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12285 a_17007_50613# a_17163_50857# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X12286 a_4461_26133# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12287 a_7986_31055# a_6909_31061# a_7824_31433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X12288 VDD a_11565_39061# a_11507_39087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X12289 VDD a_4508_65845# a_4446_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1229 a_2080_56989# a_1643_56597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12290 a_51202_58138# pmat.row_n[2] a_51694_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12291 a_9405_66627# a_9287_65087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12292 VSS pmat.row_n[9] a_23486_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12293 a_51598_11866# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12294 a_34530_21906# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12295 a_26321_46831# a_26155_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12296 a_46274_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12297 vcm a_18162_14512# a_25190_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12298 a_48586_55166# VSS a_48190_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12299 a_22628_30485# a_22871_29967# a_22979_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X123 a_14458_14191# a_9963_13967# a_14289_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1230 VDD a_45866_38279# a_46427_39009# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12300 a_11427_71017# a_11019_71543# a_11345_70773# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12301 vcm a_18162_56170# a_24186_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12302 a_6337_6825# a_5654_9527# a_6265_6825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12303 VSS VDD a_32522_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12304 a_28020_39655# a_26957_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X12305 VDD pmat.rowon_n[13] a_36142_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12306 a_24490_13874# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12307 VDD a_10943_8903# a_10378_7637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X12308 a_25190_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12309 a_36234_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1231 VDD pmat.rowon_n[5] a_19074_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12310 VDD a_7109_15521# a_6999_15645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12311 a_49590_63198# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12312 a_19166_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12313 a_22307_27791# a_22056_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X12314 VSS a_37820_30485# a_44371_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12315 a_13973_66933# a_13979_65087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12316 a_31925_40955# a_31469_40726# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12317 a_3325_43023# a_2847_43327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12318 a_36538_66210# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12319 VSS pmat.row_n[8] a_40554_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1232 VDD a_33467_46261# a_33905_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X12320 a_5132_34319# a_4918_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X12321 a_41949_30761# a_41321_30511# a_41877_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X12322 a_8491_47911# a_6787_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X12323 a_15048_44869# a_13985_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12324 a_37638_65528# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12325 a_23182_8488# a_18546_8486# a_23090_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12326 a_6292_69831# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12327 a_41162_65166# a_18162_65206# a_41254_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12328 a_14497_16367# a_12447_16143# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12329 a_47186_22950# pmat.row_n[14] a_47678_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1233 a_24186_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12330 a_1642_26935# a_1738_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12331 a_37146_55126# a_18162_55166# a_37238_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12332 a_51694_20504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12333 a_51294_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12334 VSS pmat.row_n[7] a_26498_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12335 a_23486_60186# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12336 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12337 VDD a_40951_31599# a_44741_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12338 a_23486_19898# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12339 a_37146_14918# pmat.row_n[6] a_37638_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1234 VSS a_13979_65087# a_13913_65161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X12340 VSS pmat.row_n[12] a_37542_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12341 VDD pmat.rowoff_n[7] a_44174_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12342 a_41654_12472# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12343 a_27198_72194# a_18546_72236# a_27106_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12344 a_31978_43439# a_31801_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12345 a_2847_28095# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12346 a_24586_22512# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12347 VSS a_4043_33535# a_3977_33609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X12348 VDD a_10651_42035# a_10677_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12349 VDD a_3305_17999# a_6651_22895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1235 a_14558_24233# a_14287_24349# a_14475_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12350 a_31214_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12351 VSS a_18169_31353# a_18103_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12352 VDD a_37731_44527# pmat.sample_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X12353 a_5651_66975# a_10703_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12354 a_11903_20969# a_11711_20725# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12355 a_16965_27247# a_7026_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12356 pmat.row_n[14] a_22343_50613# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X12357 VSS a_10959_23983# a_11987_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12358 VDD a_1586_33927# a_1591_36501# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12359 VDD a_10927_43421# a_10953_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1236 vcm a_18162_70226# a_42258_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12360 a_9427_50095# a_9176_50345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X12361 a_31518_71230# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12362 a_7435_68021# a_7803_67655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12363 a_4461_26133# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12364 a_35230_64162# a_18546_64204# a_35138_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12365 a_45670_11468# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12366 a_8853_48783# a_3746_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12367 a_35630_68540# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12368 a_9195_47753# a_8749_47381# a_9099_47753# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X12369 a_28110_72194# VDD a_28602_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1237 a_2865_34863# a_2659_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X12370 VDD a_22459_28879# a_27340_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X12371 a_10090_58093# a_10878_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12372 a_28602_21508# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12373 a_45966_38377# a_45866_38279# a_45884_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12374 a_28202_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12375 a_32618_70548# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12376 a_25098_14918# a_18162_14512# a_25190_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12377 a_49286_21540# a_18546_21538# a_49194_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12378 a_1881_69679# a_1846_69931# a_1643_69653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12379 VDD a_28915_50959# a_47806_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1238 a_5363_33551# a_7571_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12380 VDD a_4985_51433# a_5461_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12381 a_32126_60146# a_18162_60186# a_32218_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12382 a_2012_20541# a_1895_20346# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12383 a_2369_43389# a_2325_42997# a_2203_43401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X12384 VDD a_12128_30663# a_10287_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12385 a_5713_77295# a_5547_77295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12386 VDD nmat.rowon_n[12] a_22086_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12387 vcm a_18162_60186# a_36234_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12388 a_1846_52947# a_2124_52931# a_2080_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12389 a_31154_30083# a_30603_29575# a_31072_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1239 a_33765_40229# a_33084_40743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X12390 a_79368_39738# vcm.sky130_fd_sc_hd__nand2_1_1.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12391 a_10287_61127# a_10049_60663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12392 VDD a_6283_31591# a_7571_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12393 a_36142_64162# pmat.row_n[8] a_36634_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12394 a_3684_22729# a_2769_22357# a_3337_22325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12395 a_43566_57174# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12396 a_40650_62516# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12397 a_29114_13914# a_18162_13508# a_29206_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12398 a_8114_26703# a_7779_22583# a_8031_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12399 a_50594_58178# pmat.rowon_n[2] a_50198_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X124 VDD a_2791_57703# a_3399_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X1240 vcm a_18162_60186# a_38242_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12400 a_49194_63158# pmat.row_n[7] a_49686_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12401 a_5402_56079# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12402 a_3859_22655# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12403 a_33526_68218# pmat.rowon_n[12] a_33130_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12404 a_47278_69182# a_18546_69224# a_47186_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12405 a_44666_19500# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12406 a_20016_43781# a_18953_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12407 vcm a_18162_71230# a_26194_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12408 VDD pmat.rowon_n[10] a_29114_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12409 a_26594_63520# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1241 a_37237_29423# a_37291_29397# a_10147_29415# VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=1.105e+12p ps=1.12e+07u w=650000u l=150000u M=4
X12410 a_29367_44535# a_28245_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12411 VSS a_38711_37683# a_39505_38780# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X12412 VDD pmat.rowon_n[5] a_30118_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12413 a_12481_38870# a_12309_38659# a_12267_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X12414 vcm a_18162_65206# a_48282_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12415 a_48190_69182# pmat.row_n[13] a_48682_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12416 VDD nmat.rowon_n[4] a_21082_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12417 a_5871_32362# a_5963_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12418 VDD a_10883_3303# a_12999_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12419 a_2568_45743# a_1769_14735# a_2347_46070# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1242 a_38150_64162# pmat.row_n[8] a_38642_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12420 a_22086_68178# a_18162_68218# a_22178_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12421 a_30679_40513# a_24833_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12422 a_82815_54965# ANTENNA_fanout52_A.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12423 a_36234_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12424 a_35138_67174# a_18162_67214# a_35230_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X12425 a_1881_61885# a_1846_61651# a_1643_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12426 a_12500_31421# a_5535_29980# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12427 a_13151_10761# a_12705_10389# a_13055_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12428 VSS a_20616_27791# a_27155_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12429 a_49286_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1243 a_23700_38567# a_22541_38779# a_23604_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X12430 VSS a_7037_60729# a_6971_60797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12431 a_7829_71317# a_7663_71317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12432 VSS a_5351_60663# a_4317_62215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12433 a_11521_64239# a_5651_66975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12434 a_25098_59142# a_18162_59182# a_25190_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12435 a_20164_27791# a_19611_27247# a_19746_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12436 a_82787_26133# _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X12437 a_25190_20536# a_18546_20534# a_25098_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12438 a_39550_24918# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12439 a_45574_17890# nmat.rowon_n[6] a_45178_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1244 a_35138_23954# a_18162_23548# a_35230_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X12440 VSS a_7467_63303# a_7413_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12441 a_21478_8854# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12442 a_25590_8456# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12443 a_25292_31849# a_24861_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12444 a_43170_55126# VDD a_43662_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12445 a_2319_61493# a_2124_61635# a_2629_61885# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X12446 a_51294_24552# a_18546_24550# a_51202_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12447 a_50290_66170# a_18546_66212# a_50198_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12448 a_47278_14512# a_18546_14510# a_47186_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12449 VSS pmat.row_n[0] a_31518_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1245 VDD pmat.rowon_n[9] a_45178_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12450 a_14867_37455# a_14719_37737# a_14504_37607# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12451 VSS a_31923_42367# a_31869_42689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12452 a_11204_71855# a_11115_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=0p ps=0u w=650000u l=150000u
X12453 VDD ANTENNA_fanout52_A.DIODE a_31419_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12454 cgen.dlycontrol3_in[2] a_1591_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12455 a_46274_56130# a_18546_56172# a_46182_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12456 VSS a_26552_36165# a_26515_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12457 a_29114_58138# a_18162_58178# a_29206_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12458 a_39125_48437# a_38907_48841# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12459 nmat.col[15] a_26891_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1246 a_2843_11849# a_2493_11477# a_2748_11837# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X12460 a_1586_50247# a_1683_46295# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12461 a_23835_34191# a_11225_35836# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12462 a_6800_44629# a_6651_44661# a_7179_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12463 VDD pmat.rowon_n[2] a_50198_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12464 a_2021_9563# a_2847_8511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12465 a_49590_16886# nmat.rowon_n[7] a_49194_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12466 VSS pmat.row_n[5] a_46578_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12467 a_43566_10862# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12468 a_20570_16488# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12469 a_50594_11866# nmat.rowon_n[12] a_50198_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1247 a_41227_29423# a_40954_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12470 VDD a_30278_30511# a_33331_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12471 a_29114_17930# pmat.row_n[9] a_29606_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12472 VDD pmat.rowon_n[15] a_37146_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12473 VDD a_5331_13951# a_5318_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12474 VSS pmat.row_n[15] a_29510_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12475 VDD a_2149_45717# a_5093_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12476 VDD a_29404_36165# a_29308_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X12477 a_4853_14013# a_4809_13621# a_4687_14025# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12478 a_9367_53511# a_9639_53339# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12479 a_33622_15484# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1248 a_42658_62516# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12480 a_33526_21906# nmat.rowon_n[2] a_33130_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12481 a_30118_12910# pmat.row_n[4] a_30610_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12482 VDD a_6487_5629# a_6448_5755# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12483 VDD a_4124_18231# a_2467_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12484 a_4700_44655# a_2983_48071# a_4597_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X12485 vcm a_18162_62194# a_51294_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12486 a_9477_20291# a_9441_20189# a_9405_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12487 a_51202_66170# pmat.row_n[10] a_51694_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12488 VSS pmat.row_n[7] a_19470_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12489 a_23486_13874# nmat.rowon_n[10] a_23090_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1249 a_8727_70197# a_1674_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12490 VDD a_35715_29941# a_35646_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12491 a_25209_36965# a_22059_37683# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X12492 a_43170_72194# a_18162_72234# a_43262_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12493 a_48586_63198# pmat.rowon_n[7] a_48190_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12494 a_4951_32182# a_3746_58487# a_4492_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12495 vcm a_18162_64202# a_24186_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12496 a_34134_11906# pmat.row_n[3] a_34626_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12497 a_33130_8894# a_18162_8488# a_33222_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12498 a_45003_43343# a_44966_43255# a_44573_45173# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X12499 VSS a_9552_67191# a_8819_67197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X125 a_4703_24527# a_4259_24643# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1250 a_13979_65087# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12500 a_24094_68178# pmat.row_n[12] a_24586_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12501 a_35534_66210# pmat.rowon_n[10] a_35138_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12502 vcm a_18162_8488# a_46274_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12503 a_45270_17524# a_18546_17522# a_45178_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12504 a_36936_49257# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12505 VDD pmat.rowon_n[3] a_27106_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12506 a_45432_46983# a_43315_48437# a_45663_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12507 VDD a_4068_25615# a_7970_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12508 VSS a_14504_37607# a_12513_36924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12509 a_14458_58799# a_9963_13967# a_14289_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1251 a_16083_50069# a_19439_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X12510 vcm a_18162_68218# a_50290_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12511 VDD a_2944_69928# a_2882_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X12512 VDD nmat.rowon_n[1] a_46182_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12513 VSS a_24407_31375# a_40127_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12514 VDD a_2871_51701# a_2802_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12515 a_6777_62607# a_3866_57399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X12516 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12517 VSS VDD a_40554_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12518 a_39550_65206# pmat.rowon_n[9] a_39154_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12519 a_5696_60751# a_5497_62839# a_5506_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1252 a_27502_62194# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12520 VSS a_14653_53458# a_19441_47491# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12521 a_13329_47893# a_13462_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12522 vcm a_18162_13508# a_46274_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12523 VDD nmat.rowon_n[9] a_36142_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12524 a_4135_19391# a_3960_19465# a_4314_19453# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12525 a_4338_9839# a_3609_9295# a_4252_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12526 a_50290_11500# a_18546_11498# a_50198_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12527 a_11759_10615# comp_latch a_11993_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12528 a_25671_40719# cgen.dlycontrol3_in[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12529 a_37146_63158# a_18162_63198# a_37238_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1253 a_6772_61839# a_5081_53135# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X12530 a_51294_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12531 a_12445_12533# a_12227_12937# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X12532 a_47278_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12533 VDD a_10873_39605# a_11285_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12534 a_33130_19938# pmat.row_n[11] a_33622_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12535 a_12557_32441# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12536 a_5537_47081# a_4979_38127# a_5455_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12537 vcm a_18162_15516# a_19166_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12538 VDD a_22963_34165# a_22787_34165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X12539 VSS a_9521_31353# a_9455_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1254 a_45270_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12540 a_23182_13508# a_18546_13506# a_23090_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12541 VSS a_2659_35015# a_6651_44661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12542 vcm a_18162_10496# a_20170_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12543 a_37638_10464# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12544 a_30514_71230# pmat.rowon_n[15] a_30118_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12545 a_24946_51727# ANTENNA__1395__B1.DIODE a_24643_51959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12546 a_37238_7484# a_18546_7482# a_37146_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12547 VDD a_4037_66933# a_2944_67752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12548 vcm a_18162_19532# a_45270_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12549 a_13479_26935# a_13335_31359# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X1255 VSS a_5138_65479# a_4508_65845# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12550 a_5497_73719# a_6607_75895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12551 a_4801_69929# a_1823_74557# a_4719_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X12552 a_27198_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12553 VDD _1179_.X a_83090_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X12554 a_13456_68841# a_11837_68591# a_13361_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X12555 a_13423_55369# a_12907_54997# a_13328_55357# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X12556 a_44570_18894# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12557 a_11793_56079# a_10595_53361# a_11877_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12558 a_11987_23983# a_12245_21807# a_12147_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12559 a_35230_72194# a_18546_72236# a_35138_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1256 a_21574_9460# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12560 a_14369_61225# a_10515_61839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12561 a_6621_16885# a_3688_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X12562 a_5541_12559# a_5173_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12563 vcm a_18162_7484# a_35230_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12564 a_25098_22950# a_18162_22544# a_25190_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12565 VSS a_2315_44124# a_3241_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X12566 a_48282_71190# a_18546_71232# a_48190_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12567 VDD pmat.rowon_n[8] a_35138_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12568 a_22178_19532# a_18546_19530# a_22086_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12569 a_7088_42479# a_6173_42479# a_6741_42721# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1257 VSS pmat.row_n[4] a_31518_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12570 pmat.rowon_n[11] nmat.rowon_n[7] a_14399_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X12571 VDD pmat.rowon_n[7] a_48190_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12572 a_2557_55357# a_1923_53055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12573 VSS a_4831_34561# a_4792_34435# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12574 a_24490_62194# pmat.rowon_n[6] a_24094_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12575 VDD a_4976_16091# a_9155_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12576 VSS pmat.row_n[10] a_21478_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12577 a_22357_35877# a_21124_36391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12578 a_2748_11837# a_2129_10383# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12579 a_2672_43401# a_1757_43029# a_2325_42997# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X1258 VSS a_8481_10396# a_10047_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12580 a_8809_77117# a_8765_76725# a_8643_77129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12581 a_22449_44219# a_21124_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12582 a_36142_72194# VDD a_36634_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12583 VSS a_7079_34837# a_7013_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12584 VSS pmat.row_n[9] a_34530_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12585 a_40650_70548# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12586 a_39019_41001# a_39413_40956# a_39079_40947# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X12587 a_19413_40229# a_17996_40743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X12588 a_36634_60508# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12589 a_12174_50461# a_11455_50237# a_11611_50332# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1259 VSS pmat.row_n[11] a_31518_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12590 a_49194_71190# pmat.row_n[15] a_49686_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12591 a_44266_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12592 vcm a_18162_57174# a_22178_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12593 a_7040_8725# a_6956_8965# a_7444_8751# VSS sky130_fd_pr__nfet_01v8 ad=1.44e+11p pd=1.52e+06u as=1.341e+11p ps=1.5e+06u w=360000u l=150000u
X12594 a_50290_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12595 a_46233_43023# a_7109_29423# a_44774_40821# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12596 a_22482_14878# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12597 a_32126_9898# pmat.row_n[1] a_32618_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12598 vcm a_18162_56170# a_35230_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12599 a_11285_38870# a_11113_38659# a_11071_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X126 a_34626_12472# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1260 VDD pmat.rowon_n[1] a_35138_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12600 VDD a_24638_49159# a_23971_49140# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12601 a_8928_56457# a_7847_56085# a_8581_56053# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12602 VSS a_2411_33749# a_6601_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12603 a_35534_13874# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12604 a_6982_77295# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12605 a_14947_26159# a_14696_26409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X12606 a_26594_71552# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12607 a_47278_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12608 a_26102_61150# a_18162_61190# a_26194_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12609 a_47582_66210# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1261 a_5857_74031# a_4351_55527# a_4601_74005# VSS sky130_fd_pr__nfet_01v8 ad=5.72e+11p pd=4.36e+06u as=2.21e+11p ps=1.98e+06u w=650000u l=150000u
X12610 VSS pmat.row_n[8] a_51598_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12611 a_45178_23954# pmat.row_n[15] a_45670_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12612 a_45178_19938# a_18162_19532# a_45270_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12613 VDD a_38531_51348# pmat.col[19] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12614 VDD a_5043_57399# a_4720_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12615 VSS a_32957_30287# a_33491_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X12616 a_29676_40517# a_29772_40517# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X12617 VSS a_13479_26935# a_15395_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X12618 a_48190_55126# a_18162_55166# a_48282_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12619 vcm a_18162_18528# a_21174_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1262 nmat.rowon_n[14] a_19474_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12620 a_11965_42583# a_12061_42325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12621 a_44570_59182# pmat.rowon_n[3] a_44174_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12622 VSS pmat.row_n[0] a_41558_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12623 a_38642_18496# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12624 a_38546_24918# VSS a_38150_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12625 VDD nmat.sample_n a_18162_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X12626 VDD nmat.rowon_n[7] a_42166_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12627 a_27502_69222# pmat.rowon_n[13] a_27106_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12628 VSS pmat.row_n[10] a_24490_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12629 VDD a_13575_68743# a_13529_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1263 a_7067_53511# a_6559_33767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X12630 vcm a_18162_17524# a_34226_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12631 a_48190_14918# pmat.row_n[6] a_48682_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12632 a_22578_23516# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12633 a_22178_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12634 a_49194_18934# a_18162_18528# a_49286_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12635 a_10045_51727# a_9335_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12636 a_7810_15279# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12637 VSS a_27405_52245# pmat.col_n[7] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12638 a_10226_67503# a_9405_66627# a_10057_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X12639 a_50198_13914# a_18162_13508# a_50290_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1264 a_45670_14480# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12640 result_out[10] a_1644_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X12641 a_6607_10615# a_6879_10473# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12642 VDD a_28812_29575# a_30050_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12643 a_2325_36469# a_2107_36873# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X12644 VDD a_18243_28327# a_41335_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12645 VSS a_21124_36391# a_21087_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12646 VSS VDD a_45574_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12647 a_3801_54991# a_1823_58237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12648 a_21883_48981# a_21923_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12649 VSS pmat.row_n[9] a_28506_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1265 a_45574_20902# pmat.rowoff_n[12] a_45178_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12650 VDD nmat.rowon_n[6] a_28110_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12651 VDD a_13275_48783# a_25398_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12652 a_26194_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12653 a_3508_69135# a_3029_69135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12654 a_23090_15922# a_18162_15516# a_23182_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12655 a_46274_64162# a_18546_64204# a_46182_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12656 a_30687_48071# a_29076_48695# a_31220_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X12657 vcm a_18162_61190# a_43262_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12658 VDD a_3325_20175# a_4811_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12659 a_46674_68540# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1266 a_9217_47919# a_8907_48437# a_8079_46519# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12660 VDD pmat.rowon_n[10] a_50198_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12661 a_24405_49667# a_22499_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12662 a_20170_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12663 a_22482_55166# VSS a_22086_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12664 a_50290_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12665 a_39646_7452# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12666 a_1757_20181# a_1591_20181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12667 a_21063_48723# a_21279_48999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X12668 a_6612_15797# a_3571_13627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12669 a_2672_43401# a_1591_43029# a_2325_42997# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1267 vcm a_18162_71230# a_28202_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12670 VSS a_40349_40726# a_40591_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12671 _1519_.A a_46804_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12672 vcm.sky130_fd_sc_hd__buf_4_0.X a_77428_40594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12673 a_33222_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12674 VSS a_16689_43132# a_16381_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12675 a_19166_66170# a_18546_66212# a_19074_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12676 a_29606_13476# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12677 vcm a_18162_70226# a_51294_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12678 VDD nmat.rowon_n[12] a_33130_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12679 VDD nmat.rowon_n[4] a_19074_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1268 VDD nmat.rowon_n[14] a_31122_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12680 VDD a_24861_29673# a_24955_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X12681 vcm a_18162_60186# a_47278_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12682 VDD pmat.rowon_n[12] a_23090_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12683 a_47186_64162# pmat.row_n[8] a_47678_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12684 a_29159_37607# cgen.dlycontrol2_in[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12685 VDD a_78448_39738# a_78261_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12686 a_51694_62516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12687 VDD ANTENNA__1196__A2.DIODE a_13283_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12688 a_36466_47158# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X12689 a_12500_68021# a_11837_68591# a_12629_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X1269 a_12335_12559# a_11711_12565# a_12227_12937# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X12690 a_1846_65579# a_2163_65469# a_2121_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12691 VDD a_12069_38517# a_12481_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12692 vcm a_18162_72234# a_24186_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12693 a_37146_56130# pmat.row_n[0] a_37638_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12694 VDD cgen.dlycontrol1_in[3] a_28247_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X12695 a_25821_37483# a_24015_36911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12696 VDD pmat.rowon_n[1] a_44174_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12697 a_21082_22950# pmat.row_n[14] a_21574_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12698 a_24186_60146# a_18546_60188# a_24094_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12699 vcm a_18162_22544# a_42258_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X127 VDD a_3866_57399# a_6521_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1270 pmat.en_bit_n[0] a_17702_29967# a_18566_30287# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X12700 a_10016_30511# a_9899_30724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X12701 VDD a_12020_40871# a_10949_42364# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12702 a_27590_46831# a_2263_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12703 VDD pmat.rowon_n[11] a_27106_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12704 a_24586_64524# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12705 vcm a_18162_12504# a_38242_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12706 VSS a_10985_35516# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X12707 a_42258_10496# a_18546_10494# a_42166_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12708 VSS a_31085_27221# nmat.col[11] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12709 VSS a_19928_37253# a_19891_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X1271 VDD pmat.rowon_n[0] a_48190_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12710 a_43262_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12711 a_7631_55687# a_6559_33767# a_7805_55563# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12712 a_6087_70919# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12713 a_22745_27247# a_11067_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12714 a_44570_12870# pmat.rowoff_n[4] a_44174_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12715 a_31761_52521# ANTENNA__1197__B.DIODE pmat.col[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12716 a_8477_57141# a_8749_57141# a_9148_57487# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X12717 VDD a_17842_27497# a_39127_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12718 a_10699_75119# a_9581_73487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12719 VDD a_2727_58470# a_4165_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X1272 VSS a_13091_7655# a_13551_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12720 a_27502_22910# nmat.rowon_n[1] a_27106_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12721 VSS pmat.row_n[14] a_36538_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12722 VDD a_6700_57863# a_5528_57685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12723 a_50198_58138# a_18162_58178# a_50290_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12724 vcm a_18162_21540# a_46274_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12725 VSS a_2411_43301# a_7429_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12726 VSS a_2727_58470# a_4341_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12727 a_24895_43957# a_11149_40188# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12728 a_25098_60146# pmat.row_n[4] a_25590_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12729 a_33130_68178# a_18162_68218# a_33222_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1273 a_28602_24520# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12730 a_13531_54991# a_1957_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12731 a_18546_17522# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X12732 a_24937_41479# a_24197_42405# a_25260_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12733 VDD VDD a_24094_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12734 VSS VDD a_20474_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12735 a_50198_17930# pmat.row_n[9] a_50690_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12736 a_47278_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12737 a_26891_28327# a_44515_38645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X12738 VDD a_7730_69109# a_7674_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X12739 a_11932_59887# a_11007_58229# a_11842_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X1274 a_9161_64061# a_8782_63695# a_9089_64061# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12740 a_10969_26409# a_9075_28023# a_10873_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12741 vcm a_18162_23548# a_19166_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12742 a_6063_77295# a_5547_77295# a_5968_77295# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X12743 VSS pmat.row_n[5] a_39550_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12744 a_30514_7850# VDD a_30118_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12745 a_11145_17999# a_10975_17999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12746 a_23182_21540# a_18546_21538# a_23090_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12747 a_41254_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12748 a_43566_18894# nmat.rowon_n[5] a_43170_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12749 a_3521_33205# a_3303_33609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X1275 a_40554_69222# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12750 a_19166_11500# a_18546_11498# a_19074_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12751 a_9740_15279# a_8937_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12752 VDD a_6607_10615# a_5768_9527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X12753 VSS pmat.row_n[12] a_30514_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12754 VSS a_78802_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_1.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12755 vcm a_18162_69222# a_44266_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12756 VSS a_3746_58487# a_8133_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X12757 a_41162_19938# pmat.row_n[11] a_41654_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12758 VDD a_45645_45895# a_44635_46025# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X12759 a_6681_61839# a_5535_57993# a_6772_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1276 a_18162_57174# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X12760 a_44266_57134# a_18546_57176# a_44174_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12761 VDD a_10443_12879# a_10845_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12762 a_45861_29967# a_45019_38645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=8
X12763 VDD a_1674_68047# a_8031_76757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12764 a_2347_46070# a_1769_14735# a_2275_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X12765 a_45270_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12766 VSS pmat.row_n[6] a_44570_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12767 a_38150_10902# a_18162_10496# a_38242_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12768 a_37637_32149# a_37471_32149# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12769 VSS pmat.row_n[3] a_33526_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1277 VDD nmat.rowon_n[1] a_32126_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12770 a_22086_7890# a_18162_7484# a_22178_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12771 VDD VDD a_35138_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12772 a_30514_56170# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12773 a_27106_18934# pmat.row_n[10] a_27598_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12774 VSS VDD a_27502_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12775 VSS a_15899_47939# a_25466_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12776 VSS a_6803_77269# a_6737_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12777 a_21174_69182# a_18546_69224# a_21082_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12778 a_31614_16488# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12779 a_35230_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1278 vcm a_18162_58178# a_32218_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12780 VDD pmat.rowon_n[15] a_48190_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12781 a_32218_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12782 a_18162_72234# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X12783 a_45270_7484# a_18546_7482# a_45178_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12784 VSS a_12069_38517# a_12488_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12785 VDD a_4061_63303# a_2467_63125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X12786 a_48282_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12787 a_20475_49783# a_33685_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12788 a_35077_50345# a_10883_3303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12789 VDD vcm.sky130_fd_sc_hd__buf_4_2.A a_77428_38962# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1279 a_9963_28111# a_14471_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12790 a_21478_14878# nmat.rowon_n[9] a_21082_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12791 vcm a_18162_9492# a_50290_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12792 VDD a_11067_64015# a_17503_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X12793 a_1846_52947# a_2163_53057# a_2121_53181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X12794 a_19965_43131# a_16355_43123# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X12795 a_25190_68178# a_18546_68220# a_25098_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12796 vcm a_18162_65206# a_22178_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12797 a_22086_69182# pmat.row_n[13] a_22578_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12798 a_46182_21946# a_18162_21540# a_46274_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12799 vcm a_18162_9492# a_26194_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X128 a_32126_13914# a_18162_13508# a_32218_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1280 a_18272_35077# a_17113_34789# a_18235_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X12800 a_19176_35279# a_18999_35279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12801 VDD a_1586_33927# a_3983_41941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12802 vcm a_18162_15516# a_40250_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12803 a_43262_18528# a_18546_18526# a_43170_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12804 vcm a_18162_64202# a_35230_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12805 a_7865_59861# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12806 a_35138_68178# pmat.row_n[12] a_35630_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12807 VDD _1224_.X a_82925_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12808 a_46578_66210# pmat.rowon_n[10] a_46182_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12809 VSS a_33765_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X1281 VDD a_3571_13627# a_10791_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12810 VSS a_25667_35253# clk_dig VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X12811 a_13795_72777# a_13349_72405# a_13699_72777# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X12812 VSS a_7631_15253# a_7565_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12813 a_21395_50857# a_22199_49667# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12814 a_23182_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12815 a_19166_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12816 a_4003_7663# a_3663_9269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X12817 VSS a_4339_27804# a_11337_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X12818 a_37092_52271# ANTENNA__1395__A1.DIODE a_36789_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X12819 vcm a_18162_14512# a_44266_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1282 a_35534_12870# pmat.rowoff_n[4] a_35138_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12820 a_22988_47741# a_22276_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X12821 a_14957_52093# a_14578_51727# a_14885_52093# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X12822 a_6842_58038# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X12823 VSS VDD a_51598_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12824 a_9319_51433# a_7521_47081# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12825 VDD a_19948_51959# a_19831_51316# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X12826 a_26498_23914# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12827 a_48190_63158# a_18162_63198# a_48282_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12828 a_11506_47083# a_11784_47099# a_11740_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12829 VSS pmat.row_n[13] a_30514_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1283 a_40645_46519# a_11067_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12830 VSS ANTENNA__1196__A2.DIODE a_22463_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12831 a_6835_14735# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12832 VDD a_30857_41245# a_30463_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12833 VSS a_10049_60663# a_11969_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X12834 a_38242_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12835 a_30558_49551# ANTENNA__1184__B1.DIODE a_30255_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X12836 a_33622_57496# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12837 a_21174_14512# a_18546_14510# a_21082_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12838 a_12993_66415# a_3923_68021# a_13005_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X12839 a_20170_56130# a_18546_56172# a_20078_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1284 a_35084_31599# a_34243_32143# a_34978_31599# VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X12840 a_34226_13508# a_18546_13506# a_34134_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12841 a_2882_72221# a_2124_72123# a_2319_72092# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12842 VSS pmat.row_n[5] a_20474_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12843 a_36637_28111# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12844 VSS pmat.row_n[4] a_33526_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12845 VSS pmat.row_n[7] a_45574_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12846 a_42562_60186# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12847 a_42562_19898# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12848 a_1644_65845# a_1591_65327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12849 a_12463_22351# a_12212_22467# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1285 VSS a_82787_13077# nmat.col_n[21] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u M=2
X12850 a_25494_70226# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12851 a_13531_54991# a_12907_54997# a_13423_55369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12852 a_50198_9898# a_18162_9492# a_50290_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12853 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12854 VDD a_9367_50871# a_9319_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12855 a_11417_11177# a_9675_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12856 a_1761_2767# a_1591_2767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12857 a_23090_23954# a_18162_23548# a_23182_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12858 a_6155_49007# a_5639_49007# a_6060_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X12859 a_46274_72194# a_18546_72236# a_46182_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1286 a_41515_27497# a_21739_29415# a_41297_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12860 a_13290_50345# a_11067_49871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12861 a_14001_65871# a_13432_62581# a_13919_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12862 a_39154_24958# VDD a_39646_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12863 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top vcm.sky130_fd_sc_hd__buf_4_1.X vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X12864 a_28940_41831# a_27877_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X12865 a_26102_9898# a_18162_9492# a_26194_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12866 a_43662_22512# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12867 VDD a_38851_28327# a_47035_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12868 VSS a_27411_46805# a_27345_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12869 a_77245_40202# a_77341_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1287 VSS a_20616_27791# a_25040_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12870 a_22063_46519# clk_ena VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12871 VDD pmat.rowon_n[8] a_46182_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12872 a_2672_36873# a_1757_36501# a_2325_36469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12873 a_22482_63198# pmat.rowon_n[7] a_22086_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12874 VSS a_3325_40847# a_4535_38377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12875 a_50290_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12876 a_28506_61190# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12877 a_9759_70045# a_9135_69679# a_9651_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12878 a_30118_71190# a_18162_71230# a_30210_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12879 VSS pmat.row_n[10] a_32522_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1288 VDD a_2655_72373# a_1823_74557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12880 VDD a_10873_38517# a_11285_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12881 VDD pmat.rowon_n[0] a_36142_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12882 a_25466_47919# a_19541_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12883 ANTENNA__1190__A2.DIODE a_46863_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X12884 a_9135_23983# a_7415_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12885 a_47186_72194# VDD a_47678_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12886 VDD nmat.rowon_n[1] a_20078_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12887 vcm a_18162_58178# a_20170_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12888 a_11921_50095# a_11542_50461# a_11849_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12889 a_51694_70548# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1289 a_84028_9615# ANTENNA__1190__A1.DIODE a_83922_9615# VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X12890 a_44174_14918# a_18162_14512# a_44266_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12891 a_47678_60508# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12892 a_19166_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12893 a_25221_46519# a_11067_30287# a_25384_46403# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12894 a_51202_60146# a_18162_60186# a_51294_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12895 vcm a_18162_57174# a_33222_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12896 a_11823_46973# a_5363_33551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12897 a_34134_70186# a_18162_70226# a_34226_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X12898 a_2203_20553# a_1757_20181# a_2107_20553# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12899 a_33526_14878# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X129 a_44266_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1290 a_4865_8181# a_4503_6335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12900 a_9511_28879# a_4068_25615# a_9405_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
X12901 VSS a_2939_45503# a_2873_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X12902 a_24586_72556# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12903 vcm a_18162_20536# a_38242_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12904 VDD nmat.rowon_n[2] a_24094_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12905 a_17625_42902# a_17113_41317# a_18176_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12906 VSS a_3923_68021# a_12067_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12907 VSS a_13503_39069# a_13443_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12908 a_21174_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12909 a_24094_62154# a_18162_62194# a_24186_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1291 a_2325_27765# a_2107_28169# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X12910 VDD a_1923_61759# a_2464_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12911 a_45574_67214# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12912 VSS pmat.row_n[1] a_36538_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12913 VDD a_42240_29423# a_42701_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X12914 a_34245_48169# _1154_.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12915 a_2215_34141# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12916 a_8459_56457# a_8013_56085# a_8363_56457# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X12917 a_11892_21959# a_12311_19783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12918 a_16837_42043# a_15420_41831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X12919 a_7217_53609# a_7163_53333# a_5211_57172# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1292 VDD nmat.rowon_n[9] a_22086_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12920 a_47026_45519# a_40105_47375# a_46857_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X12921 a_46578_9858# nmat.rowon_n[14] a_46182_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12922 _0467_ a_9528_20407# a_14925_24847# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12923 a_4496_28335# a_4379_28548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X12924 VDD pmat.rowoff_n[4] a_27106_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12925 a_25190_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12926 a_32035_38825# a_30913_38779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12927 VDD a_4705_39759# a_5671_40097# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12928 VSS pmat.row_n[11] a_22482_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12929 a_45670_63520# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1293 vcm a_18162_21540# a_37238_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12930 a_34530_9858# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12931 vcm a_18162_18528# a_32218_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12932 a_13917_72373# a_13699_72777# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X12933 a_49686_18496# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12934 a_2847_38975# a_2672_39049# a_3026_39037# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12935 a_46135_38127# a_45884_38377# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12936 a_31518_17890# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12937 VDD nmat.rowon_n[4] a_40158_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12938 VSS a_5415_71543# a_4409_74183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12939 a_39550_58178# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1294 VSS a_17054_28995# a_17306_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12940 a_41162_68178# a_18162_68218# a_41254_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12941 VDD a_2683_22089# a_9291_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12942 VDD a_14641_57167# a_14839_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12943 VDD pmat.rowon_n[7] a_22086_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12944 VSS a_9919_51959# a_9827_53379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12945 VDD nmat.rowon_n[5] a_26102_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12946 a_13439_74575# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X12947 a_11895_66959# a_11797_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12948 a_30278_30511# a_29931_30517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X12949 a_44266_65166# a_18546_65208# a_44174_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1295 a_13805_42919# a_14113_43132# a_13779_43123# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X12950 a_44666_69544# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12951 a_6925_51183# a_6883_51335# a_6835_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X12952 a_29308_36165# a_28245_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12953 VSS a_10873_38517# a_11292_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12954 a_1941_47375# a_1769_14735# a_1857_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12955 a_38557_48469# a_38391_48469# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12956 a_2672_36873# a_1591_36501# a_2325_36469# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12957 a_44174_59142# a_18162_59182# a_44266_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12958 VDD a_1586_63927# a_1591_63701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12959 a_19074_61150# pmat.row_n[5] a_19566_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1296 a_20078_70186# pmat.row_n[14] a_20570_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12960 a_19566_8456# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12961 VDD a_18563_27791# a_39496_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12962 a_14287_57280# a_10515_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X12963 a_27106_69182# a_18162_69222# a_27198_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12964 VDD a_7865_59861# a_7895_60214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12965 VSS pmat.row_n[1] a_29510_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12966 a_36324_46983# a_36539_47113# a_36466_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X12967 a_31214_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12968 a_33526_55166# VSS a_33130_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12969 a_17012_47349# a_16863_47428# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1297 a_2319_59036# a_2124_59067# a_2629_58799# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X12970 a_20503_48981# a_20659_49140# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12971 VDD pmat.rowon_n[13] a_21082_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12972 a_22427_31421# a_20310_28029# a_22064_31287# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12973 a_45178_65166# pmat.row_n[9] a_45670_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12974 VSS a_78802_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_0.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12975 VDD a_40352_41831# a_39781_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X12976 a_1846_59051# a_2163_58941# a_2121_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12977 a_5408_56399# a_5211_57172# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X12978 pmat.rowoff_n[14] a_14839_70223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12979 a_21174_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1298 a_46182_10902# pmat.row_n[2] a_46674_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12980 a_2107_8585# a_1757_8213# a_2012_8573# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X12981 VSS nmat.en_bit_n[2] a_35534_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12982 a_34530_63198# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12983 VDD a_7040_8725# a_7094_9117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12984 a_21478_66210# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12985 a_45574_20902# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12986 VSS pmat.row_n[15] a_48586_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12987 VDD a_33341_37692# a_32947_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12988 a_14107_39958# a_12969_40175# a_14035_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12989 vcm a_18162_23548# a_40250_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1299 VSS a_46386_33231# _1194_.A2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u M=16
X12990 a_31339_31787# a_18563_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X12991 vcm a_18162_72234# a_35230_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12992 a_39246_16520# a_18546_16518# a_39154_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12993 a_22578_65528# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12994 a_48190_56130# pmat.row_n[0] a_48682_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12995 a_32126_22950# pmat.row_n[14] a_32618_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12996 a_25190_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12997 a_22086_55126# a_18162_55166# a_22178_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12998 VSS pmat.row_n[7] a_38546_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12999 a_22361_41479# a_22357_43493# a_23479_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13 a_28079_38825# a_26957_38779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X130 a_41663_47893# a_42191_48071# a_42138_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=150000u
X1300 result_out[5] a_1644_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X13000 a_42562_13874# nmat.rowon_n[10] a_42166_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13001 VDD a_10055_31591# a_15757_52535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13002 pmat.col[10] a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X13003 VDD a_30663_50087# a_34425_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13004 a_22086_14918# pmat.row_n[6] a_22578_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13005 a_25590_17492# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13006 VSS pmat.row_n[12] a_22482_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13007 a_25494_23914# pmat.rowoff_n[15] a_25098_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13008 a_22063_46519# clk_ena a_22297_46653# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13009 a_47043_29423# a_41731_49525# a_47212_29673# VSS sky130_fd_pr__nfet_01v8 ad=7.605e+11p pd=7.54e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X1301 a_20170_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13010 a_21239_47349# a_21215_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X13011 VSS pmat.row_n[14] a_47582_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13012 a_78448_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_0.X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13013 a_39154_58138# pmat.row_n[2] a_39646_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13014 VSS a_3859_56311# a_3225_55509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13015 a_46817_27221# a_17139_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X13016 a_39550_11866# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13017 a_7067_60470# a_6816_60699# a_6608_60663# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13018 VDD a_1643_67477# a_1591_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13019 a_11877_12565# a_11711_12565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1302 a_40250_61150# a_18546_61192# a_40158_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13020 a_24833_40719# a_24667_40719# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X13021 a_4309_37921# a_4127_37013# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13022 a_15093_39638# a_13985_40229# a_15048_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13023 VSS pmat.row_n[6] a_37542_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13024 a_26102_13914# pmat.row_n[5] a_26594_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13025 VDD a_29711_47679# a_29076_48695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X13026 a_4337_22351# a_3859_22655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13027 VDD a_1923_53055# a_1643_58773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13028 a_20170_64162# a_18546_64204# a_20078_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13029 a_41558_60186# pmat.rowon_n[4] a_41162_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1303 a_11743_55329# a_4128_64391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13030 a_30610_11468# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13031 a_41558_19898# nmat.rowon_n[4] a_41162_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13032 a_29606_55488# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13033 a_20570_68540# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13034 a_2319_56860# a_2163_56765# a_2464_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X13035 VDD a_2676_29941# a_2586_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13036 VSS a_7589_33749# a_7523_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13037 VDD a_31412_43439# a_31518_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13038 VSS a_13739_51701# a_13432_62581# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X13039 a_34226_21540# a_18546_21538# a_34134_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1304 VSS a_2411_43301# a_8257_54269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13040 VSS a_26479_32117# a_40678_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X13041 VDD a_23455_32447# a_23442_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13042 a_5597_44807# a_2389_45859# a_5747_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13043 a_13349_72405# a_13183_72405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13044 VSS a_2163_53057# a_2124_52931# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13045 a_19470_14878# nmat.rowon_n[9] a_19074_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13046 VDD a_31701_37462# a_30765_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X13047 VDD VSS a_38150_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13048 a_9103_56383# a_8928_56457# a_9282_56445# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13049 a_42258_58138# a_18546_58180# a_42166_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1305 a_10851_30485# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13050 VSS pmat.row_n[2] a_29510_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13051 a_2325_34017# a_2107_33775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X13052 ANTENNA__1187__B1.DIODE a_46636_36469# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u M=4
X13053 VDD ANTENNA__1197__A.DIODE a_35802_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X13054 VDD a_8581_56053# a_8471_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X13055 a_14058_8207# a_12981_8213# a_13896_8585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13056 vcm a_18162_60186# a_21174_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13057 a_21082_64162# pmat.row_n[8] a_21574_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13058 VSS a_2835_13077# a_13317_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13059 VDD config_1_in[15] a_1591_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1306 a_29114_20942# pmat.row_n[12] a_29606_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13060 a_82788_10357# ANTENNA__1190__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=0p ps=0u w=650000u l=150000u
X13061 a_34134_63158# pmat.row_n[7] a_34626_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13062 a_39646_20504# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13063 a_22541_39867# a_21124_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X13064 a_11910_47197# a_11784_47099# a_11506_47083# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13065 VDD VDD a_46182_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13066 a_39246_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13067 a_39003_47753# a_38557_47381# a_38907_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13068 a_2957_58255# a_2603_58368# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13069 a_32218_69182# a_18546_69224# a_32126_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1307 a_44570_68218# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13070 a_25190_8488# a_18546_8486# a_25098_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13071 a_46274_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13072 VDD a_24374_29941# a_24131_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13073 a_5687_38279# a_5671_40097# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X13074 a_29206_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13075 a_46023_32937# a_40951_31599# a_45805_32661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13076 a_5508_18543# a_5257_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X13077 a_2191_27412# a_2283_27221# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X13078 VDD a_1687_13621# a_1717_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X13079 a_44174_22950# a_18162_22544# a_44266_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1308 VDD a_9643_66389# a_9601_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13080 a_11409_34789# a_10953_34951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13081 a_41254_19532# a_18546_19530# a_41162_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13082 a_19166_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13083 a_10325_62985# a_9135_62613# a_10216_62985# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13084 a_35517_30333# a_35039_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13085 vcm a_18162_65206# a_33222_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13086 a_36538_61190# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13087 a_33130_69182# pmat.row_n[13] a_33622_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13088 VSS a_77528_39738# a_77341_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13089 VSS pmat.row_n[10] a_40554_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1309 a_29114_16926# a_18162_16520# a_29206_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13090 a_19470_71230# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13091 a_6700_57863# a_6835_51183# a_6842_58038# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X13092 VDD a_4719_30287# a_5383_48783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13093 a_18162_69222# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13094 a_46947_39215# a_46705_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u M=3
X13095 VDD a_2944_52789# a_2882_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X13096 VSS a_14071_8511# a_14005_8585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X13097 a_10167_16950# a_8305_20871# a_10095_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X13098 a_44791_43541# a_31675_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X13099 VSS a_6830_44655# a_6747_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X131 a_77245_39738# a_77341_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1310 VDD pmat.rowon_n[2] a_39154_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13100 vcm a_18162_10496# a_29206_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13101 a_21174_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13102 a_14911_31965# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13103 a_14829_29423# a_14466_28879# a_14745_29423# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=2.43e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13104 vcm a_18162_57174# a_41254_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13105 a_34226_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13106 a_13145_26935# a_13683_24847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13107 a_41558_14878# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13108 a_7165_13353# a_6763_13103# a_7001_13103# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X13109 a_24490_24918# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1311 a_33222_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13110 a_9521_31353# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13111 a_30514_17890# nmat.rowon_n[6] a_30118_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13112 VSS a_44763_34293# a_45107_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13113 a_11271_73085# a_7658_71543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13114 VDD a_35108_39655# a_35012_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13115 VDD a_2325_42997# a_2215_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13116 VSS a_7109_29423# a_44733_44431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13117 a_38546_58178# pmat.rowon_n[2] a_38150_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13118 a_2012_16189# a_1895_15994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X13119 a_26331_42089# a_25209_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1312 a_30118_11906# a_18162_11500# a_30210_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13120 a_45670_71552# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13121 VDD a_22393_37692# a_21999_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13122 a_2882_65693# a_2124_65595# a_2319_65564# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13123 a_2244_26935# rst_n VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13124 vcm a_18162_16520# a_28202_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13125 a_49286_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13126 VDD a_10873_36341# a_10817_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13127 a_26609_51433# a_23395_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13128 a_32218_14512# a_18546_14510# a_32126_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13129 a_31214_56130# a_18546_56172# a_31122_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1313 a_2398_51859# a_2715_51969# a_2673_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X13130 a_27443_32463# a_24374_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13131 VDD a_2839_38101# a_2743_38279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X13132 VDD a_4339_27804# a_10029_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13133 VSS a_4339_27804# a_9779_26819# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13134 VSS a_3123_27399# a_2743_28853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13135 a_27502_15882# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13136 VSS a_2419_69455# a_1899_35051# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X13137 VSS pmat.row_n[5] a_31518_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13138 VSS a_14347_69831# a_12719_69367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13139 a_23389_32521# a_22199_32149# a_23280_32521# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X1314 VSS pmat.row_n[0] a_43566_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13140 VDD pmat.rowon_n[15] a_22086_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13141 VDD a_8695_12801# a_8656_12675# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13142 VSS a_3571_13627# a_12815_8213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13143 a_48586_8854# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13144 VSS pmat.row_n[10] a_43566_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13145 a_44571_32143# a_44320_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X13146 VSS a_12235_39913# a_13259_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13147 a_41654_23516# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13148 a_41254_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13149 VSS a_27313_51701# pmat.col_n[1] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1315 VDD nmat.rowon_n[15] a_47186_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13150 a_44266_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13151 VSS a_3339_59879# a_13593_74941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13152 VDD nmat.rowon_n[5] a_34134_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13153 a_33526_63198# pmat.rowon_n[7] a_33130_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13154 a_13273_10357# a_13055_10761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X13155 a_34816_34191# a_34639_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13156 VDD a_2939_45503# a_2926_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13157 a_20474_66210# pmat.rowon_n[10] a_20078_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13158 VDD a_39321_42333# a_38927_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13159 a_30210_17524# a_18546_17522# a_30118_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1316 a_8568_26703# a_8031_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X13160 VDD a_14933_37429# a_14963_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13161 VDD nmat.rowon_n[6] a_47186_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13162 a_44666_14480# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13163 a_45270_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13164 a_42166_15922# a_18162_15516# a_42258_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13165 a_41162_8894# pmat.row_n[0] a_41654_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13166 a_18162_22544# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13167 a_27598_24520# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13168 a_11464_48285# a_10795_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13169 a_27355_28995# a_25315_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1317 a_36288_44527# a_36111_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13170 VDD nmat.rowon_n[1] a_31122_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13171 VDD a_43776_30287# a_44741_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13172 VDD a_3305_27791# a_5070_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X13173 VDD a_8735_54207# a_8722_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13174 VDD a_18243_28327# a_27535_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13175 a_35534_8854# nmat.rowon_n[15] a_35138_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13176 a_5779_13255# a_5173_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X13177 a_51694_8456# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13178 a_24490_65206# pmat.rowon_n[9] a_24094_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13179 vcm a_18162_13508# a_31214_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1318 a_6369_39465# a_4533_38279# a_6369_39215# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13180 VDD nmat.rowon_n[9] a_21082_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13181 a_39246_24552# a_18546_24550# a_39154_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13182 VSS a_16171_40157# a_16111_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13183 a_38242_66170# a_18546_66212# a_38150_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13184 a_48682_13476# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13185 a_45178_10902# pmat.row_n[2] a_45670_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13186 nmat.col[24] _1154_.X a_83170_5263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X13187 a_31095_42367# cgen.dlycontrol4_in[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X13188 a_2834_26525# a_1757_26159# a_2672_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13189 a_5989_38377# a_4533_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1319 a_39550_11866# nmat.rowon_n[12] a_39154_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13190 VDD pmat.rowon_n[12] a_42166_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13191 a_22086_63158# a_18162_63198# a_22178_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13192 a_28110_20942# pmat.row_n[12] a_28602_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13193 a_10153_60137# a_10058_60431# a_8841_60405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13194 a_43566_68218# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13195 a_28110_16926# a_18162_16520# a_28202_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13196 VDD pmat.rowon_n[2] a_38150_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13197 a_32218_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13198 VSS a_25802_48169# a_25785_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X13199 VSS pmat.row_n[0] a_33526_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X132 a_4529_68367# a_4075_68583# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1320 a_33382_46983# a_14887_46377# a_33596_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X13200 a_38546_11866# nmat.rowon_n[12] a_38150_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13201 a_4933_45199# a_4313_44111# a_4745_45519# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X13202 a_35138_62154# a_18162_62194# a_35230_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13203 VSS a_12309_38659# a_39387_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13204 a_27502_56170# pmat.rowon_n[0] a_27106_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13205 VSS a_12875_16341# a_12809_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13206 VDD nmat.rowon_n[10] a_25098_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13207 VSS _1192_.B1 a_25224_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13208 VSS a_10873_36341# a_10817_36694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13209 a_22578_10464# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1321 VDD a_2163_56765# a_2124_56891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13210 a_14471_62063# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13211 vcm a_18162_62194# a_39246_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13212 a_39154_66170# pmat.row_n[10] a_39646_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13213 a_43262_60146# a_18546_60188# a_43170_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13214 a_43662_64524# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13215 a_40158_61150# pmat.row_n[5] a_40650_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13216 a_37238_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13217 a_14458_5487# _1187_.A2 a_14289_5737# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13218 vcm a_18162_19532# a_30210_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13219 VDD a_2511_34319# a_2411_33749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X1322 a_3399_62607# a_2215_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13220 a_13884_71311# a_3615_71631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X13221 a_5746_11703# a_2021_9563# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13222 a_6646_24527# a_5991_23983# a_6564_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13223 a_32162_34191# a_31985_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13224 a_46973_33775# a_30571_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13225 a_11113_38659# a_13801_38779# a_14864_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13226 a_25879_31591# a_44763_34293# a_44371_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X13227 VSS a_13459_28111# a_47947_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13228 a_20170_72194# a_18546_72236# a_20078_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13229 a_9919_51959# a_9213_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1323 nmat.col_n[2] ANTENNA__1395__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X13230 VSS a_42769_50069# pmat.col_n[23] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13231 VDD pmat.rowon_n[13] a_19074_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13232 VDD nmat.rowon_n[4] a_51202_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13233 a_2980_29967# a_2500_30345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13234 VSS a_45019_38645# a_46636_36469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X13235 VSS cgen.dlycontrol4_in[0] a_29627_43983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X13236 a_33222_71190# a_18546_71232# a_33130_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13237 VDD pmat.rowon_n[8] a_20078_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13238 a_44174_60146# pmat.row_n[4] a_44666_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13239 a_35138_8894# a_18162_8488# a_35230_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1324 a_19074_12910# pmat.row_n[4] a_19566_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13240 VDD a_7693_22365# a_12294_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13241 a_29206_61150# a_18546_61192# a_29114_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13242 VDD a_5271_35407# a_5550_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X13243 vcm a_18162_68218# a_38242_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13244 a_30118_7890# VDD a_30610_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13245 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X13246 a_21187_28335# a_10223_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13247 VDD pmat.rowon_n[7] a_33130_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13248 VSS config_2_in[12] a_1591_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13249 VDD a_13091_52047# a_18011_50729# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1325 a_12128_32375# a_9135_60967# a_12270_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13250 a_8655_76751# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X13251 VDD a_46263_52245# pmat.col[27] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X13252 VSS a_2007_25597# a_35277_30333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13253 a_12472_35077# a_11409_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X13254 a_21082_72194# VDD a_21574_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13255 a_1757_33775# a_1591_33775# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13256 VSS pmat.row_n[2] a_27502_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13257 a_38242_11500# a_18546_11498# a_38150_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13258 a_21574_60508# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13259 a_15383_42089# a_14261_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1326 a_23582_10464# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13260 a_34134_71190# pmat.row_n[15] a_34626_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13261 a_4319_15039# a_4144_15113# a_4498_15101# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13262 a_11499_71017# a_11115_71285# a_11427_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13263 a_4503_6335# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13264 a_39246_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13265 a_2122_13779# a_2400_13763# a_2356_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13266 a_13909_68047# a_3615_71631# a_13575_68743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13267 VDD a_5579_12394# a_5779_13255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13268 a_35534_61190# pmat.rowon_n[5] a_35138_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13269 a_2873_45577# a_1683_45205# a_2764_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1327 a_45246_41167# a_35312_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13270 a_10811_77437# a_7658_71543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13271 VDD a_6424_55687# a_5955_55223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13272 a_37497_38550# a_36341_39141# a_37404_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13273 VSS a_10651_24617# a_10287_24759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X13274 a_28202_22544# a_18546_22542# a_28110_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13275 a_28131_50069# a_38851_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X13276 a_32218_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13277 a_25209_42043# a_23700_42919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13278 a_46182_18934# pmat.row_n[10] a_46674_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13279 a_43566_21906# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1328 VSS pmat.row_n[12] a_21478_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13280 VSS VDD a_46578_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13281 a_18546_55168# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13282 a_50690_16488# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13283 VSS a_39781_40157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X13284 a_40250_69182# a_18546_69224# a_40158_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13285 a_19582_46983# a_19678_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13286 a_32522_66210# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13287 VDD a_6927_30503# a_9195_58951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13288 a_36234_59142# a_18546_59184# a_36142_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13289 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1329 a_47582_59182# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13290 a_39246_7484# a_18546_7482# a_39154_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13291 VSS a_9827_53379# a_10449_53153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13292 a_14569_16367# a_10515_13967# a_14497_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13293 a_30118_23954# pmat.row_n[15] a_30610_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13294 a_30118_19938# a_18162_19532# a_30210_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13295 a_4130_77117# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13296 a_2215_8207# a_1591_8213# a_2107_8585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13297 a_11358_73309# a_11232_73211# a_10954_73195# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=360000u l=150000u
X13298 a_39550_60186# pmat.rowon_n[4] a_39154_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13299 a_39550_19898# nmat.rowon_n[4] a_39154_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X133 a_31165_29199# a_13641_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.9e+11p pd=3.8e+06u as=0p ps=0u w=650000u l=150000u
X1330 a_41162_61150# pmat.row_n[5] a_41654_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13300 VSS pmat.row_n[8] a_36538_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13301 VDD a_3577_70197# a_2944_72104# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13302 a_40554_14878# nmat.rowon_n[9] a_40158_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13303 a_33130_55126# a_18162_55166# a_33222_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13304 VDD a_2468_21959# a_2099_21237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13305 VSS pmat.row_n[7] a_49590_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13306 a_23582_18496# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13307 a_23486_24918# VSS a_23090_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13308 a_20078_15922# pmat.row_n[7] a_20570_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13309 a_38557_47381# a_38391_47381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1331 a_27198_20536# a_18546_20534# a_27106_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13310 a_3026_64061# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13311 vcm a_18162_65206# a_41254_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13312 VDD a_9581_56079# a_12021_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13313 a_41162_69182# pmat.row_n[13] a_41654_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13314 vcm a_18162_55166# a_37238_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13315 VSS _1183_.A2 a_14734_4175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13316 a_33130_14918# pmat.row_n[6] a_33622_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13317 a_37146_59142# pmat.row_n[3] a_37638_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13318 a_34134_18934# a_18162_18528# a_34226_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13319 VDD a_6835_51183# a_6914_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1332 vcm a_18162_19532# a_31214_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13320 a_26498_57174# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13321 a_10287_24759# a_9528_20407# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13322 VSS a_35007_44527# a_35113_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13323 a_12757_36950# a_12585_37179# a_12543_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13324 VSS a_77528_40202# a_77341_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13325 a_26498_15882# pmat.rowoff_n[7] a_26102_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13326 a_36634_9460# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13327 VSS VDD a_30514_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13328 a_45199_44905# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13329 VDD a_40105_47375# a_44963_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1333 VSS a_7370_27791# a_7663_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13330 a_17234_46403# a_10515_13967# a_17138_46403# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13331 vcm a_18162_24552# a_28202_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13332 vcm a_18162_66210# a_27198_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13333 a_38242_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13334 VDD nmat.rowon_n[14] a_46182_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13335 a_31214_64162# a_18546_64204# a_31122_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13336 a_31614_68540# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13337 a_27598_58500# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13338 VDD a_12263_50959# a_17183_51817# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13339 VSS a_28867_40871# a_13909_39605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1334 VSS pmat.row_n[1] a_51598_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13340 a_6451_67655# a_13158_71285# a_13884_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13341 a_7631_75895# a_6975_76823# a_7805_76001# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13342 VSS pmat.row_n[3] a_27502_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13343 a_34134_9898# pmat.row_n[1] a_34626_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13344 a_11921_10749# a_10839_11989# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13345 a_4443_62063# a_4413_62037# a_4349_62063# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X13346 VDD a_13091_28327# a_38293_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X13347 vcm a_18162_16520# a_36234_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13348 VDD vcm.sky130_fd_sc_hd__buf_4_2.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=4.74e+06u w=500000u l=500000u M=2
X13349 a_8256_20291# a_7644_16341# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1335 a_45178_16926# pmat.row_n[8] a_45670_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13350 a_40250_14512# a_18546_14510# a_40158_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13351 a_40554_71230# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13352 VSS pmat.row_n[8] a_39550_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13353 vcm a_18162_60186# a_32218_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13354 a_6649_41935# a_6369_39465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13355 vcm a_18162_15516# a_49286_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13356 a_32126_64162# pmat.row_n[8] a_32618_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13357 a_37638_21508# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13358 VDD a_12813_31029# a_12703_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13359 vcm a_18162_10496# a_50290_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1336 a_29510_8854# nmat.rowon_n[15] a_29114_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13360 a_37238_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13361 a_6884_74183# a_7092_74005# a_7026_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13362 a_2163_58941# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13363 a_8325_10901# a_1717_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13364 VSS a_2099_24746# a_1895_23610# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13365 a_44266_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13366 a_23033_28879# a_21341_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13367 a_22086_56130# pmat.row_n[0] a_22578_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13368 a_44570_70226# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13369 a_26194_15516# a_18546_15514# a_26102_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1337 VSS pmat.row_n[11] a_34530_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13370 vcm a_18162_12504# a_23182_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13371 a_42166_23954# a_18162_23548# a_42258_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13372 VSS a_2419_53351# a_2419_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X13373 VSS a_10651_44211# a_10591_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13374 a_38150_13914# a_18162_13508# a_38242_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13375 VSS a_38972_39655# a_38935_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13376 a_7797_63151# a_7321_63151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X13377 a_26102_55126# VDD a_26594_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13378 a_33765_39141# a_32072_38567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13379 a_47724_47081# ANTENNA__1197__B.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1338 VSS _1187_.A2 a_14458_5487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X13380 a_47582_61190# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13381 VSS pmat.row_n[14] a_21478_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13382 vcm a_18162_21540# a_31214_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13383 VDD a_3295_40277# a_3234_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13384 a_14475_24233# a_14287_24349# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13385 VSS pmat.row_n[10] a_51598_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13386 vcm a_18162_11500# a_27198_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13387 VSS a_41731_49525# a_28131_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13388 a_35630_24520# nmat.en_bit_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13389 VDD _1179_.X a_25590_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1339 a_24407_31375# a_44811_36469# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X13390 a_28110_24958# a_18162_24552# a_28202_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13391 a_18947_49811# a_19283_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X13392 VDD pmat.rowon_n[10] a_38150_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13393 VDD a_16113_52271# a_16863_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X13394 a_26498_10862# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13395 a_32218_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13396 a_6984_64015# a_5307_67655# a_6794_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13397 a_38242_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13398 a_1757_18005# a_1591_18005# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13399 VSS pmat.row_n[5] a_24490_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X134 VSS a_1858_25615# a_20217_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1340 a_6435_34863# a_5989_34863# a_6339_34863# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X13400 a_27531_51727# ANTENNA__1197__B.DIODE a_27313_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13401 a_9528_20407# a_12875_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X13402 VDD a_2325_36469# a_2215_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13403 VSS a_4068_25615# a_7888_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13404 vcm a_18162_70226# a_39246_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13405 a_25129_31751# a_20616_27791# a_25292_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13406 a_14261_42043# a_13227_42333# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13407 VSS a_22499_49783# a_22199_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13408 a_37542_7850# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13409 a_36142_20942# pmat.row_n[12] a_36634_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1341 VDD a_10878_58487# a_11797_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.62e+12p ps=1.524e+07u w=1e+06u l=150000u M=4
X13410 a_6619_56311# a_3339_70759# a_6793_56417# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13411 a_43662_72556# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13412 a_36142_16926# a_18162_16520# a_36234_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13413 a_8479_11484# a_8511_10422# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13414 a_39646_62516# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13415 a_40250_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13416 VDD a_30641_44743# a_31976_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X13417 VDD pmat.rowon_n[4] a_43170_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13418 vcm a_18162_59182# a_25190_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13419 a_5821_18785# a_5603_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1342 VSS a_8267_49159# a_8091_49192# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13420 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X13421 VSS VDD a_47582_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13422 a_26102_72194# a_18162_72234# a_26194_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13423 VDD a_11797_60431# a_11797_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13424 VSS pmat.row_n[4] a_28506_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13425 VSS a_4403_51701# a_1923_53055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X13426 VSS pmat.row_n[11] a_28506_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13427 a_25494_16886# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13428 a_12543_36950# a_12585_37179# a_12543_37277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13429 a_30913_39867# a_29772_40517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1343 a_36234_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13430 a_30210_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13431 a_14491_51969# a_5363_33551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13432 a_23090_10902# a_18162_10496# a_23182_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13433 VDD VDD a_20078_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13434 a_37542_69222# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13435 a_28506_9858# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13436 VDD nmat.rowon_n[1] a_29114_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13437 a_20170_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13438 vcm a_18162_58178# a_29206_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13439 VDD pmat.rowon_n[15] a_33130_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1344 a_20316_47607# a_18823_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X13440 VSS pmat.row_n[11] a_41558_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13441 vcm a_18162_18528# a_51294_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13442 a_37519_46983# a_37791_46811# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X13443 a_39307_27791# a_25879_31591# a_39089_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13444 a_18953_43493# a_17996_41831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13445 pmat.rowon_n[9] a_14734_64015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13446 a_33222_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13447 a_45133_38155# a_44444_32233# a_45047_38155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13448 a_45270_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13449 a_40650_7452# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1345 a_26355_29673# a_25315_28335# a_24374_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X13450 a_38150_58138# a_18162_58178# a_38242_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13451 VDD nmat.rowon_n[9] a_19074_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13452 a_3227_22351# a_2603_22357# a_3119_22729# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X13453 a_25718_32463# a_25688_32117# a_25423_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13454 VDD a_15101_29423# a_24959_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13455 a_8581_73461# a_8363_73865# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X13456 a_31221_32143# a_1781_9308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X13457 a_31122_21946# a_18162_21540# a_31214_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13458 VDD VDD a_50198_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13459 VDD a_22787_34165# a_11921_37462# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1346 VSS pmat.row_n[3] a_24490_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13460 a_27106_11906# a_18162_11500# a_27198_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13461 a_38150_17930# pmat.row_n[9] a_38642_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13462 a_42658_15484# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13463 VDD nmat.rowon_n[5] a_45178_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13464 VSS a_2847_63999# a_2781_64073# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X13465 a_37291_29397# a_44449_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u M=2
X13466 a_9552_67191# a_9405_66627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13467 a_31518_66210# pmat.rowon_n[10] a_31122_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13468 a_2886_25071# a_2648_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13469 VSS _1194_.B1 a_13257_4175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1347 a_1757_23445# a_1591_23445# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13470 VDD a_11927_27399# a_17047_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13471 VSS pmat.row_n[2] a_35534_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13472 a_82971_11989# _1194_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X13473 a_6583_62607# a_6175_60039# a_6777_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13474 a_7258_40303# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13475 a_32522_7850# VDD a_32126_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13476 a_46182_69182# a_18162_69222# a_46274_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13477 VSS pmat.row_n[1] a_48586_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13478 VDD a_33007_37683# a_33033_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X13479 a_50290_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1348 a_35230_12504# a_18546_12502# a_35138_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13480 VDD a_19488_52423# a_14287_69455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X13481 VDD ANTENNA__1395__A1.DIODE a_47035_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13482 a_36234_67174# a_18546_67216# a_36142_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13483 a_43170_11906# pmat.row_n[3] a_43662_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13484 a_22499_49783# a_36265_48981# a_36209_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13485 a_28506_64202# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13486 a_6976_32375# a_4128_64391# a_7118_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X13487 a_2419_69455# a_4025_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13488 VDD pmat.rowon_n[13] a_40158_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13489 a_1757_50095# a_1591_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1349 a_45178_8894# a_18162_8488# a_45270_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13490 a_49286_66170# a_18546_66212# a_49194_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13491 VDD pmat.rowon_n[3] a_36142_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13492 a_22269_40391# a_21621_40955# a_22743_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13493 VDD nmat.rowon_n[4] a_49194_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13494 a_40250_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13495 a_33130_63158# a_18162_63198# a_33222_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13496 VDD config_1_in[13] a_1591_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13497 VSS a_14641_57167# a_14839_70223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13498 a_23182_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13499 a_20078_66170# a_18162_66210# a_20170_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X135 pmat.en_bit_n[0] a_17702_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X1350 a_33309_36039# a_33489_36603# a_34611_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X13500 a_25494_57174# pmat.rowon_n[1] a_25098_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13501 a_19566_16488# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13502 VSS a_13091_52047# a_18568_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13503 a_47975_46831# a_47724_47081# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13504 vcm a_18162_63198# a_37238_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13505 a_22933_32117# a_22715_32521# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13506 a_24094_7890# a_18162_7484# a_24186_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13507 a_37146_67174# pmat.row_n[11] a_37638_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13508 a_11325_76457# a_10239_77295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X13509 a_2971_53903# a_1591_52815# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1351 a_22578_16488# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13510 a_41654_65528# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13511 VDD a_13979_65087# a_13966_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13512 a_9417_5737# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X13513 a_11317_40188# a_10979_43222# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13514 a_51202_22950# pmat.row_n[14] a_51694_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13515 a_41162_55126# a_18162_55166# a_41254_55126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13516 a_34226_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13517 a_8197_64789# a_8031_64789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13518 a_2843_11849# a_2327_11477# a_2748_11837# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13519 VSS pmat.row_n[7] a_30514_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1352 vcm a_18162_68218# a_39246_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13520 a_30189_48437# a_29076_48695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X13521 a_5935_6575# a_5654_9527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13522 VDD a_1586_50247# a_5639_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13523 a_37542_22910# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13524 a_14708_31599# a_4707_32156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13525 a_12249_71311# a_11893_71427# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13526 a_44570_23914# pmat.rowoff_n[15] a_44174_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13527 a_41162_14918# pmat.row_n[6] a_41654_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13528 VSS pmat.row_n[12] a_41558_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13529 a_7026_74031# a_2407_49289# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1353 VSS a_5363_12015# a_5012_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13530 VSS a_28915_50959# a_47407_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13531 VDD a_11091_26311# a_11041_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13532 VDD a_24867_53135# a_47861_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X13533 a_31214_72194# a_18546_72236# a_31122_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13534 a_44666_56492# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13535 a_24094_24958# VDD a_24586_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13536 VDD a_11113_38659# a_14864_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13537 a_27198_62154# a_18546_62196# a_27106_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13538 a_43720_32143# a_43543_32151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13539 a_19965_43131# a_16355_43123# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1354 a_40158_7890# VDD a_40650_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13540 a_27598_66532# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13541 pmat.rowoff_n[14] a_14839_70223# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X13542 VSS a_6612_66933# a_4298_67191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X13543 a_3480_17143# a_3688_17179# a_3622_17277# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X13544 VSS a_82789_26677# nmat.col[29] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13545 VSS a_37813_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X13546 VDD pmat.rowon_n[8] a_31122_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13547 a_34530_15882# pmat.rowoff_n[7] a_34134_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13548 a_27106_56130# a_18162_56170# a_27198_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13549 a_4312_74005# a_4601_74005# a_4535_74031# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X1355 VSS a_6611_57399# a_6559_57167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13550 VDD a_14647_51701# a_14578_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13551 vcm a_18162_24552# a_36234_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13552 VDD a_3727_66113# a_3688_65987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13553 a_14905_28585# a_14365_22351# a_14833_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13554 VDD pmat.rowon_n[0] a_21082_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13555 VSS VDD a_39550_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13556 a_48682_55488# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13557 vcm a_18162_23548# a_49286_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13558 a_32126_72194# VDD a_32618_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13559 a_43566_70226# pmat.rowon_n[14] a_43170_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1356 vcm a_18162_63198# a_40250_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13560 a_35630_58500# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13561 VDD a_5579_12394# a_6763_13103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X13562 a_28110_62154# pmat.row_n[6] a_28602_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13563 a_32618_60508# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13564 VSS pmat.row_n[3] a_35534_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13565 a_49286_11500# a_18546_11498# a_49194_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13566 a_25997_42902# a_25209_42043# a_26331_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13567 a_10979_43222# a_11021_43011# a_10979_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13568 a_8038_10927# a_1717_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13569 a_47673_51433# _1154_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1357 a_6607_75895# a_6799_75637# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X13570 a_6524_65327# a_3866_57399# a_6334_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13571 a_2672_64073# a_1591_63701# a_2325_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13572 VSS pmat.row_n[2] a_48586_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13573 a_33601_30761# a_7415_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13574 VDD a_3688_17179# a_7131_19407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13575 VSS a_19689_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X13576 a_5341_59317# a_4719_58255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13577 VDD VSS a_25098_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13578 a_14471_27497# a_11091_26311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13579 a_26194_23548# a_18546_23546# a_26102_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1358 a_40158_67174# pmat.row_n[11] a_40650_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13580 vcm a_18162_20536# a_23182_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13581 VSS a_16381_35286# a_17867_34473# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13582 a_46578_61190# pmat.rowon_n[5] a_46182_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13583 a_27623_52521# a_23395_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13584 a_9839_47679# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13585 VSS a_9963_13967# a_14458_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X13586 a_15655_50613# a_12263_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13587 a_30514_67214# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13588 a_45064_44807# a_44966_43255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13589 VDD a_13549_8181# a_13439_8207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1359 a_5692_55509# a_5784_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13590 a_3687_14735# a_3063_14741# a_3579_15113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13591 a_19166_8488# a_18546_8486# a_19074_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13592 VDD a_1781_9308# a_1725_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13593 a_51294_69182# a_18546_69224# a_51202_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13594 a_25494_10862# nmat.rowon_n[13] a_25098_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13595 a_19332_41959# a_19428_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13596 a_47278_59142# a_18546_59184# a_47186_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13597 a_5353_35407# a_4601_35727# a_5271_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13598 a_2007_49770# a_2099_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X13599 a_1757_33775# a_1591_33775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X136 VDD a_32256_44869# a_32160_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X1360 VDD a_7109_29423# a_46013_42997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X13600 a_20474_59182# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13601 a_48282_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13602 vcm a_18162_61190# a_26194_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13603 VSS pmat.row_n[8] a_47582_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13604 a_51598_14878# nmat.rowon_n[9] a_51202_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13605 a_30610_63520# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13606 VDD pmat.rowoff_n[12] a_35138_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13607 a_34626_18496# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13608 a_38242_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13609 a_2163_74173# a_1674_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1361 VSS _1154_.A a_82818_69135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X13610 vcm a_18162_55166# a_48282_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13611 a_6699_76983# a_6795_76989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X13612 a_48190_59142# pmat.row_n[3] a_48682_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13613 VDD a_1586_50247# a_1683_45205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13614 a_24490_58178# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13615 a_23395_53135# a_26891_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13616 a_4918_34319# a_4792_34435# a_4514_34451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13617 a_3684_22729# a_2603_22357# a_3337_22325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13618 a_19689_41317# a_19233_41479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13619 a_1586_63927# a_1644_57141# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X1362 a_39246_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13620 a_36142_24958# a_18162_24552# a_36234_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13621 a_31210_31751# a_31217_29429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X13622 a_39646_70548# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13623 a_40250_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13624 a_36161_37462# a_36341_38053# a_37404_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13625 vcm a_18162_67214# a_25190_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13626 a_36234_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13627 VDD a_30663_50087# ANTENNA__1395__A2.DIODE VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13628 a_36538_69222# pmat.rowon_n[13] a_36142_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13629 a_39154_60146# a_18162_60186# a_39246_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1363 a_20695_32447# a_20520_32521# a_20874_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13630 a_7578_16694# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13631 vcm a_18162_17524# a_43262_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13632 VSS a_14589_35286# a_13653_35516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X13633 a_49286_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13634 a_10747_6727# a_9668_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13635 VSS a_28704_29568# a_28626_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13636 a_17573_27791# _0467_ a_17845_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X13637 nmat.col[16] a_26891_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X13638 a_25190_10496# a_18546_10494# a_25098_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13639 a_30121_31599# a_30527_31573# a_29635_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.1125e+11p ps=1.95e+06u w=650000u l=150000u
X1364 VDD a_40837_46261# a_44389_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.44e+12p ps=2.288e+07u w=1e+06u l=150000u M=8
X13640 VDD a_36193_35805# a_35799_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13641 a_5029_45199# a_2983_48071# a_4933_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13642 a_7674_69135# a_4991_69831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13643 a_6821_18543# a_6343_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13644 a_10957_28879# a_10609_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X13645 VSS pmat.row_n[9] a_37542_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13646 a_30118_65166# pmat.row_n[9] a_30610_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13647 vcm a_18162_16520# a_47278_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13648 a_13795_10687# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13649 pmat.col_n[11] ANTENNA__1187__B1.DIODE a_30479_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1365 a_5505_53387# a_2419_53351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13650 a_51294_14512# a_18546_14510# a_51202_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13651 VDD a_3615_71631# a_4503_70455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13652 VSS a_25575_31055# a_39666_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X13653 a_50290_56130# a_18546_56172# a_50198_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13654 VSS pmat.row_n[1] a_38546_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13655 VSS a_22879_41781# a_11921_41814# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13656 a_46578_15882# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13657 a_2325_8181# a_2107_8585# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13658 VSS nmat.en_C0_n a_20474_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13659 a_14277_11471# a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1366 a_9529_51005# a_9463_50877# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13660 a_19697_28335# a_6664_26159# a_19405_28853# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X13661 VSS a_32871_49007# a_9411_2215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X13662 VDD a_34553_42658# a_34552_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13663 VSS pmat.row_n[5] a_50594_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13664 a_20078_57134# pmat.row_n[1] a_20570_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13665 a_48586_9858# nmat.rowon_n[14] a_48190_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13666 a_1925_20871# cgen.dlycontrol4_in[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13667 VDD a_35559_30209# a_35520_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13668 VSS pmat.row_n[15] a_33526_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13669 a_30514_20902# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1367 a_22825_50345# a_21371_50087# a_22753_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13670 VDD a_1674_68047# a_5547_77295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13671 VDD pmat.rowon_n[5] a_37146_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13672 a_10693_74031# a_10515_75895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X13673 a_7212_62607# a_6583_62607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X13674 a_33130_56130# pmat.row_n[0] a_33622_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13675 VSS a_1781_9308# a_1725_12342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13676 a_24186_16520# a_18546_16518# a_24094_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13677 a_5455_46831# a_5173_45993# a_5633_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X13678 a_1846_74283# a_2124_74299# a_2080_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13679 a_42258_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1368 a_6927_30503# a_10851_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X13680 VDD a_10190_60663# a_10287_61127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13681 a_10595_53361# a_10205_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X13682 a_18162_56170# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13683 a_19470_17890# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13684 a_1757_15829# a_1591_15829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13685 VDD a_3295_23060# a_2907_22522# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13686 a_24374_29941# a_25681_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13687 VSS pmat.row_n[7] a_23486_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13688 a_34828_41605# a_33765_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X13689 a_20474_12870# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1369 VSS pmat.row_n[2] a_28506_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13690 a_46763_44431# a_7109_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X13691 VSS a_2655_59317# a_1823_60949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13692 a_45574_62194# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13693 VDD a_2715_51969# a_2676_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13694 VSS a_20329_35431# a_17675_37001# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13695 a_2319_56860# a_2124_56891# a_2629_56623# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X13696 a_28506_72234# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13697 VSS a_29404_36165# a_29367_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13698 VDD a_21124_42919# a_21028_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13699 VSS pmat.row_n[14] a_32522_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X137 a_34768_47375# a_32687_46607# a_35186_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X1370 a_25494_55166# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13700 a_24094_58138# pmat.row_n[2] a_24586_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13701 VDD pmat.rowon_n[11] a_36142_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13702 a_46934_53135# ANTENNA__1197__B.DIODE a_46765_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X13703 a_24490_11866# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13704 VDD a_6799_75637# a_6699_76983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13705 a_46674_24520# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13706 a_3061_11445# a_2843_11849# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13707 a_36234_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13708 VDD nmat.rowon_n[1] a_50198_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13709 vcm a_18162_58178# a_50290_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1371 a_30210_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13710 a_19832_37253# a_18769_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13711 VSS pmat.row_n[6] a_22482_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13712 VSS a_16926_46261# a_13091_18535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X13713 VSS a_25221_46519# a_25189_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13714 a_19166_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13715 a_1644_64213# a_1823_64213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13716 a_36538_64202# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13717 a_49286_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13718 a_8625_56445# a_8581_56053# a_8459_56457# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13719 a_23033_27791# ANTENNA__1395__B1.DIODE nmat.col_n[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 a_26594_7452# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13720 a_36538_22910# nmat.rowon_n[1] a_36142_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13721 a_19268_34191# a_19091_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13722 VDD nmat.rowon_n[9] a_40158_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13723 a_7578_16367# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13724 a_9869_62581# a_9651_62985# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X13725 VSS a_30819_40191# a_30765_40513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13726 VDD VSS a_23090_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13727 a_33491_32463# a_29163_29423# a_33395_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13728 a_2250_70045# a_2124_69947# a_1846_69931# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13729 a_41162_63158# a_18162_63198# a_41254_63158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1373 a_22482_7850# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13730 a_47186_20942# pmat.row_n[12] a_47678_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13731 VDD a_24833_34191# a_26659_34967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13732 a_47186_16926# a_18162_16520# a_47278_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13733 VSS pmat.row_n[0] a_27502_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13734 a_25209_44581# a_23700_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X13735 a_11427_73180# a_11271_73085# a_11572_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X13736 a_51294_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13737 VDD a_12585_40443# a_16612_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13738 a_37146_12910# pmat.row_n[4] a_37638_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13739 VDD a_13779_36595# a_13805_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1374 a_42307_31756# a_35244_32411# a_42783_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X13740 VSS a_12449_22895# a_13013_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13741 a_10979_42895# a_10725_43222# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13742 a_10167_17277# a_9913_16950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13743 VDD nmat.rowon_n[10] a_44174_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13744 a_41654_10464# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13745 a_27198_70186# a_18546_70228# a_27106_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13746 a_29510_66210# pmat.rowon_n[10] a_29114_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13747 a_43659_28853# a_43451_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13748 a_30015_51727# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X13749 a_24586_20504# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1375 a_32836_50345# _1183_.A2 a_32371_50247# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13750 VDD pmat.rowoff_n[15] a_27106_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13751 VSS a_5351_19913# a_13955_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.554e+11p ps=1.58e+06u w=420000u l=150000u
X13752 VDD VDD a_31122_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13753 a_24186_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13754 a_11905_74895# a_10515_75895# a_11823_74895# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13755 VDD ANTENNA__1395__A1.DIODE a_22195_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13756 a_27106_64162# a_18162_64202# a_27198_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13757 a_2104_45565# a_1987_45370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13758 a_48586_69222# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13759 a_31214_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1376 a_40554_22910# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13760 VSS a_37291_29397# a_47043_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13761 VSS a_5597_44807# a_5566_44905# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13762 VDD clk_dig a_7387_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X13763 a_31869_42689# a_24833_40719# a_31783_42689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13764 a_20570_8456# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13765 VSS a_1923_69823# a_2893_72765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13766 VSS config_1_in[15] a_1591_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13767 VDD a_13432_62581# a_13205_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X13768 a_5688_52423# a_5784_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X13769 a_35230_62154# a_18546_62196# a_35138_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1377 a_37146_21946# a_18162_21540# a_37238_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13770 VDD a_28704_29568# a_43533_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13771 VSS a_3746_58487# a_9481_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X13772 a_35630_66532# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13773 a_28110_70186# pmat.row_n[14] a_28602_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13774 VSS pmat.row_n[3] a_42562_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13775 VDD nmat.rowon_n[15] a_30118_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13776 a_28202_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13777 a_25098_12910# a_18162_12504# a_25190_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13778 a_5318_13647# a_4241_13653# a_5156_14025# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13779 a_48282_61150# a_18546_61192# a_48190_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1378 VSS a_1899_35051# a_6311_42692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13780 a_18241_31698# a_20695_32447# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X13781 VDD config_2_in[14] a_1591_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13782 a_44917_43023# a_44739_43567# a_44573_45173# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X13783 a_21478_61190# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13784 a_26957_37691# a_26501_37462# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X13785 a_12381_63151# a_11883_62063# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13786 a_36142_62154# pmat.row_n[6] a_36634_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13787 a_3495_62927# a_1823_64213# a_3305_62607# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X13788 VSS a_17285_32117# nmat.rowoff_n[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13789 VSS pmat.row_n[2] a_46578_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1379 a_29206_67174# a_18546_67216# a_29114_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13790 a_40650_60508# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13791 a_43566_55166# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13792 a_34277_38550# a_33765_39141# a_34828_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13793 a_3225_74941# a_2747_74549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13794 a_7001_17027# a_3688_17179# a_6929_17027# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13795 a_28628_27247# a_9411_2215# a_28325_27221# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X13796 VSS pmat.row_n[12] a_29510_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13797 a_49194_61150# pmat.row_n[5] a_49686_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13798 a_37497_38550# a_36341_39141# a_37463_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13799 VDD a_25850_48981# a_18823_50247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X138 a_11479_18543# a_9441_20189# a_11116_18695# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1380 VSS a_7717_14735# a_37237_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13800 a_83007_26703# ANTENNA__1395__B1.DIODE a_82789_26677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13801 a_43274_47919# a_30111_47911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13802 a_47278_67174# a_18546_67216# a_47186_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13803 nmat.en_bit_n[1] a_16966_29673# a_17830_29423# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X13804 VSS a_12851_28853# a_18566_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13805 cgen.dlycontrol4_in[0] a_1626_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13806 a_20619_49551# a_20175_49667# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X13807 VDD pmat.rowon_n[13] a_51202_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13808 VDD a_23700_42919# a_23604_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13809 a_23043_28335# a_22792_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X1381 VSS a_1769_14735# a_1769_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=2
X13810 VSS a_4075_31591# a_12332_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13811 vcm a_18162_8488# a_41254_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13812 a_9313_26409# a_4339_27804# a_9217_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13813 a_23486_58178# pmat.rowon_n[2] a_23090_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13814 a_5265_14025# a_4075_13653# a_5156_14025# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13815 a_37542_71230# pmat.rowon_n[15] a_37146_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13816 a_30610_71552# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13817 a_51294_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13818 a_2007_21482# a_2099_21237# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X13819 VDD a_21981_34191# a_25647_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1382 VSS VDD a_32522_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13820 VDD pmat.rowon_n[8] a_29114_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13821 a_26594_61512# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13822 a_34226_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13823 VSS a_20534_35431# a_20329_35431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13824 a_12407_28853# a_8583_29199# a_12689_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X13825 a_5506_60751# a_5535_57993# a_5696_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13826 a_51294_8488# a_18546_8486# a_51202_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13827 a_51598_66210# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13828 a_19441_47491# a_16800_47213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13829 a_4165_67753# a_2791_57703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1383 a_4249_9615# a_2021_11043# a_4167_9615# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13830 vcm a_18162_63198# a_48282_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13831 VDD a_36324_46983# a_35540_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13832 VSS a_10751_71543# a_9279_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13833 a_48190_67174# pmat.row_n[11] a_48682_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13834 VDD pmat.rowon_n[0] a_19074_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13835 a_21007_51843# a_10515_13967# a_20911_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13836 a_42562_24918# VSS a_42166_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13837 a_36234_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13838 a_13290_50095# a_12044_49641# a_13290_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X13839 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.sky130_fd_sc_hd__buf_4_0.X vcm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X1384 a_14453_31599# a_14287_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13840 a_42658_57496# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13841 a_48586_22910# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13842 VSS a_30255_49783# pmat.col[11] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13843 VSS a_6787_47607# a_6292_65479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13844 a_14427_46519# a_14699_46377# a_14657_46403# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13845 a_23239_37217# a_14600_37607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13846 a_35138_24958# nmat.en_bit_n[2] a_35630_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13847 a_23663_44535# a_22541_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13848 VSS a_7631_75895# a_6051_74183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13849 a_25098_57134# a_18162_57174# a_25190_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1385 a_11317_40188# a_10979_43222# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13850 VSS a_12247_20175# a_12252_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13851 VDD a_30663_50087# a_35353_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13852 a_45574_15882# pmat.rowoff_n[7] a_45178_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13853 VSS pmat.row_n[4] a_42562_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13854 VSS a_12044_49641# a_12002_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13855 VDD a_4809_28577# a_4699_28701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13856 a_2781_64073# a_1591_63701# a_2672_64073# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13857 a_11877_56079# a_11835_56311# a_11793_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13858 a_12147_24233# a_7026_24527# a_11987_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13859 a_2950_74707# a_3228_74691# a_3184_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1386 VDD pmat.rowon_n[13] a_33130_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13860 VDD nmat.rowon_n[6] a_32126_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13861 vcm a_18162_24552# a_47278_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13862 a_2107_28169# a_1757_27797# a_2012_28157# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X13863 vcm a_18162_66210# a_46274_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13864 a_2219_4943# a_1775_5059# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X13865 VSS a_3305_15823# a_6621_16885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13866 a_30210_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13867 a_50290_64162# a_18546_64204# a_50198_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13868 a_50690_68540# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13869 VSS a_22063_46519# a_21837_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1387 a_47278_17524# a_18546_17522# a_47186_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13870 a_46674_58500# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13871 a_28110_9898# pmat.row_n[1] a_28602_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13872 a_6909_31061# a_6743_31061# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13873 VSS a_19689_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X13874 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X13875 a_49590_14878# nmat.rowon_n[9] a_49194_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13876 VSS pmat.row_n[3] a_46578_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13877 VDD a_41926_46983# a_42617_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13878 a_5595_19958# a_4523_21276# a_5136_19783# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13879 VSS a_6981_28879# a_7109_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1388 a_21124_36391# a_19965_36603# a_21087_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X13880 vcm a_18162_7484# a_30210_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13881 a_29114_15922# pmat.row_n[7] a_29606_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13882 VSS pmat.row_n[13] a_29510_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13883 VSS a_7578_48553# a_7373_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13884 a_24186_24552# a_18546_24550# a_24094_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13885 a_23182_66170# a_18546_66212# a_23090_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13886 a_33622_13476# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13887 a_30118_10902# pmat.row_n[2] a_30610_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13888 a_19166_56130# a_18546_56172# a_19074_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13889 vcm a_18162_60186# a_51294_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1389 a_19470_71230# pmat.rowon_n[15] a_19074_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13890 a_15393_28879# a_14943_26703# a_15299_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X13891 a_51202_64162# pmat.row_n[8] a_51694_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13892 VDD pmat.rowon_n[2] a_23090_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13893 VSS pmat.row_n[5] a_19470_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13894 a_5402_56079# a_4259_73807# a_5245_56053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X13895 a_23486_11866# nmat.rowon_n[12] a_23090_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13896 VDD a_6559_33767# a_7217_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13897 VSS a_6612_65845# a_5267_65479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X13898 ANTENNA__1184__B1.DIODE a_47212_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X13899 a_41162_56130# pmat.row_n[0] a_41654_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X139 a_4725_53359# a_4659_53738# a_4653_53359# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1390 a_33222_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13900 a_14565_3855# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13901 a_43170_70186# a_18162_70226# a_43262_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13902 vcm a_18162_62194# a_24186_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13903 a_5257_62215# a_4985_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13904 a_24094_66170# pmat.row_n[10] a_24586_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13905 a_35534_64202# pmat.rowon_n[8] a_35138_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13906 VSS a_27785_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X13907 VDD a_27579_34967# a_14600_37607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X13908 a_45270_15516# a_18546_15514# a_45178_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13909 vcm a_18162_12504# a_42258_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1391 a_30118_56130# a_18162_56170# a_30210_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13910 a_9217_49257# a_8907_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13911 a_36234_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13912 a_2935_38279# a_2847_38975# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X13913 a_24857_50959# _1224_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13914 VDD pmat.rowoff_n[12] a_46182_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13915 a_18566_30287# a_12461_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13916 a_8915_6409# a_8399_6037# a_8820_6397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13917 a_3843_17277# a_3305_15823# a_3480_17143# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13918 a_19689_34789# a_17996_35303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X13919 a_36538_72234# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1392 a_4241_28335# a_4075_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13920 a_49286_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13921 a_5012_42301# a_4432_42313# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13922 a_4705_39759# a_4351_39872# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13923 VSS pmat.row_n[14] a_40554_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13924 a_3484_58229# a_3938_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13925 a_11506_47083# a_11823_46973# a_11781_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13926 a_35534_58178# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13927 a_49590_71230# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13928 vcm a_18162_11500# a_46274_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13929 VDD pmat.rowoff_n[4] a_36142_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1393 pmat.col[30] ANTENNA__1197__B.DIODE a_47775_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X13930 a_6141_44629# a_6732_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13931 vcm a_18162_68218# a_23182_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13932 a_26272_44869# a_25209_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X13933 a_4351_55527# a_2315_44124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13934 a_47186_24958# a_18162_24552# a_47278_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13935 a_51294_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13936 a_47278_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13937 a_11071_36694# a_11041_36596# a_10999_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13938 VSS pmat.row_n[5] a_43566_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13939 a_40554_17890# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1394 a_44570_21906# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13940 vcm a_18162_13508# a_19166_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13941 a_2847_38975# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13942 a_37542_8854# nmat.rowon_n[15] a_37146_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13943 a_24719_36341# a_24895_36341# a_24847_36367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X13944 a_76962_40202# a_77058_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13945 a_23182_11500# a_18546_11498# a_23090_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13946 VSS pmat.row_n[15] a_26498_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13947 a_6412_8725# a_6872_8725# a_6830_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13948 a_10216_62985# a_9301_62613# a_9869_62581# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13949 a_24186_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1395 a_12967_58559# a_12792_58633# a_13146_58621# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13950 a_9556_62973# a_6175_60039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X13951 a_12040_16367# a_11881_16911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13952 a_9521_31353# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13953 vcm a_18162_59182# a_44266_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13954 VSS a_1923_69823# a_2985_74941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13955 a_27198_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13956 a_20474_61190# pmat.rowon_n[5] a_20078_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13957 a_14287_50345# a_14249_49525# a_14369_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X13958 a_44570_16886# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13959 a_35230_70186# a_18546_70228# a_35138_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1396 VSS a_42240_29423# a_43605_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13960 VDD a_34002_44527# a_34547_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13961 VDD a_6799_75637# a_6757_75663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X13962 a_42166_10902# a_18162_10496# a_42258_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13963 a_10405_64239# a_5363_70543# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X13964 a_11703_48156# a_11508_48187# a_12013_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X13965 a_10045_54697# a_6559_33767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13966 a_14649_29423# a_12461_29673# a_14553_29423# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X13967 a_31122_18934# pmat.row_n[10] a_31614_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13968 VSS VDD a_31518_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13969 a_25098_20942# a_18162_20536# a_25190_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1397 a_47186_57134# pmat.row_n[1] a_47678_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13970 a_28202_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13971 a_31761_52521# ANTENNA__1395__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13972 VDD a_4955_40277# a_6637_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13973 a_45529_51157# a_17139_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13974 VDD pmat.rowon_n[6] a_35138_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13975 a_4901_30753# a_4683_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13976 VDD a_32957_30287# a_33331_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13977 a_21174_59142# a_18546_59184# a_21082_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13978 VDD pmat.rowon_n[5] a_48190_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13979 VDD a_9668_10651# a_10233_7913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1398 VDD a_12445_58229# a_12335_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X13980 a_24490_60186# pmat.rowon_n[4] a_24094_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13981 a_37709_52245# a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13982 a_39246_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13983 a_24490_19898# nmat.rowon_n[4] a_24094_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13984 VSS pmat.row_n[8] a_21478_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13985 VDD ANTENNA__1190__A1.DIODE a_29187_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13986 a_36142_70186# pmat.row_n[14] a_36634_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13987 VSS pmat.row_n[7] a_34530_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13988 a_9797_9813# a_1717_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13989 a_43566_63198# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1399 a_51694_55488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13990 a_9902_18115# a_9557_17705# a_9820_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13991 a_13163_10383# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X13992 VSS a_4697_74005# a_4312_74005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13993 VDD a_24833_34191# a_26475_34343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13994 a_25190_58138# a_18546_58180# a_25098_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13995 vcm a_18162_55166# a_22178_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13996 a_22086_59142# pmat.row_n[3] a_22578_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13997 VSS a_4863_13077# a_4379_13818# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13998 a_46182_11906# a_18162_11500# a_46274_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13999 VSS a_28116_38567# a_28079_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14 VDD pmat.rowon_n[6] a_44174_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X140 a_4349_35407# a_4307_35639# a_4267_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1400 VSS a_4123_16042# a_3367_14906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14000 pmat.row_n[8] a_19675_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14001 VDD a_7037_60729# a_7067_60470# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14002 a_32126_7890# VDD a_32618_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14003 a_50594_66210# pmat.rowon_n[10] a_50198_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14004 VSS a_16745_34427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X14005 a_35138_58138# pmat.row_n[2] a_35630_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14006 VDD a_5659_38127# a_6061_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14007 a_5589_14967# a_5451_14557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14008 a_35534_11866# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14009 a_26498_7850# VDD a_26102_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1401 VSS VDD a_42562_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14010 VSS a_4257_34319# a_4267_35407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14011 VSS a_27789_36039# a_28171_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14012 VSS a_33011_29941# a_32957_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14013 VDD VDD a_29114_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14014 a_47278_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14015 VDD a_10055_31591# a_14565_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14016 a_9148_57487# a_4128_64391# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X14017 a_39127_29423# a_37827_30793# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14018 VDD a_33309_41479# a_34552_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X14019 a_10377_32509# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1402 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14020 a_7895_58294# a_5535_57993# a_7436_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14021 a_23182_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14022 a_28876_47741# a_28639_47081# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X14023 a_22365_32149# a_22199_32149# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14024 VDD a_4503_6335# a_4490_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14025 a_47582_64202# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14026 VDD a_9339_28335# a_9741_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14027 a_26576_46831# a_25681_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X14028 a_11071_36367# a_10817_36694# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14029 a_45178_21946# pmat.row_n[13] a_45670_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1403 a_31122_23954# pmat.row_n[15] a_31614_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14030 a_13768_22325# a_4523_21276# a_13717_21583# VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14031 VDD a_1923_69823# a_2464_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14032 VDD nmat.rowon_n[9] a_51202_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14033 a_45178_17930# a_18162_17524# a_45270_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14034 VSS a_4516_21531# a_9323_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14035 a_22459_28879# a_22015_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14036 a_12857_31421# a_12813_31029# a_12691_31433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X14037 VSS a_32371_47349# a_31105_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14038 VDD a_2325_63669# a_2215_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14039 a_37542_56170# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1404 a_22463_52047# ANTENNA__1195__A1.DIODE pmat.col_n[2] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X14040 a_6881_5487# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14041 a_15489_29199# a_15435_29111# a_15299_28879# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X14042 a_7436_58487# a_5535_57993# a_7578_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14043 vcm a_18162_16520# a_21174_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14044 a_44570_57174# pmat.rowon_n[1] a_44174_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14045 a_38642_16488# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14046 a_42065_50345# a_28131_50069# pmat.col[23] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X14047 a_27502_67214# pmat.rowon_n[11] a_27106_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14048 VSS pmat.row_n[8] a_24490_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14049 vcm a_18162_15516# a_34226_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1405 a_5629_24233# a_2952_25045# a_5547_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14050 VSS a_31925_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X14051 VSS a_9581_56079# a_11829_55329# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14052 a_5809_51335# a_2389_45859# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14053 a_48190_12910# pmat.row_n[4] a_48682_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14054 a_22578_21508# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14055 a_22178_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14056 a_40099_52245# ANTENNA__1187__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X14057 a_25098_65166# a_18162_65206# a_25190_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14058 a_6699_76983# a_6975_76823# a_6933_77117# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14059 nmat.col_n[4] a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X1406 a_31122_19938# a_18162_19532# a_31214_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14060 VDD a_38905_28853# a_41949_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X14061 a_17191_48981# a_17139_49551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X14062 a_2007_42644# a_2051_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X14063 a_25117_39141# a_23700_39655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X14064 a_20438_35431# a_11497_40719# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14065 VDD a_5363_33551# a_19439_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14066 VSS a_10575_15253# a_10509_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14067 VDD a_17811_39605# a_17635_39605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14068 pmat.rowon_n[5] a_11067_16359# a_14655_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14069 a_2840_55509# a_1591_54991# a_3063_55535# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X1407 a_22063_46519# a_13275_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X14070 VDD pmat.rowoff_n[7] a_28110_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14071 a_50290_72194# a_18546_72236# a_50198_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14072 a_46383_47695# a_33423_47695# a_45450_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14073 a_23090_13914# a_18162_13508# a_23182_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14074 VSS a_2683_22089# a_9135_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14075 a_31249_28879# a_19405_28853# a_31165_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14076 a_7109_29423# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X14077 a_46274_62154# a_18546_62196# a_46182_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14078 a_12658_42895# a_12481_42895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14079 VDD pmat.rowon_n[13] a_49194_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1408 a_34626_65528# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14080 a_46674_66532# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14081 a_43170_63158# pmat.row_n[7] a_43662_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14082 a_34724_44527# a_34547_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14083 VDD a_11007_58229# a_11842_59887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14084 VDD a_31425_37218# a_31976_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X14085 VSS a_19817_37692# a_19509_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14086 VSS config_1_in[13] a_1591_22351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14087 VDD a_28915_50959# a_32871_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14088 VDD pmat.rowon_n[8] a_50198_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14089 a_1644_57141# a_1674_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1409 vcm a_18162_13508# a_48282_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14090 VSS _1196_.B1 pmat.col_n[31] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14091 a_46182_56130# a_18162_56170# a_46274_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14092 a_3503_19087# a_2879_19093# a_3395_19465# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X14093 a_7004_66959# a_6970_67191# a_6749_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X14094 a_32522_61190# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14095 a_29114_66170# a_18162_66210# a_29206_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14096 VSS a_5935_46983# a_5893_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14097 vcm a_18162_71230# a_20170_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14098 a_38642_9460# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14099 a_2369_36861# a_2325_36469# a_2203_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X141 a_1683_48169# a_1739_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1410 a_8103_53903# a_7479_53909# a_7995_54281# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X14100 a_29606_11468# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14101 a_24895_38517# a_12345_39100# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14102 a_19166_64162# a_18546_64204# a_19074_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14103 VDD pmat.rowon_n[0] a_40158_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14104 a_20570_24520# nmat.en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14105 a_19566_68540# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14106 a_51202_72194# VDD a_51694_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14107 a_40250_7484# a_18546_7482# a_40158_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14108 VDD pmat.rowon_n[10] a_23090_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14109 a_47186_62154# pmat.row_n[6] a_47678_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1411 a_30210_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14110 a_33519_46831# a_33839_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14111 VDD nmat.rowon_n[14] a_48190_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14112 a_16377_38779# a_15921_38550# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X14113 a_51694_60508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14114 a_23182_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14115 VSS a_5329_54965# a_4587_53505# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X14116 VSS a_1781_9308# a_28639_47081# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14117 VSS a_54790_39198# comp.adc_nor_latch_0.R VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.65e+11p ps=1.66e+06u w=500000u l=150000u M=2
X14118 a_7534_37039# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14119 vcm a_18162_70226# a_24186_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1412 a_33423_47695# a_6664_26159# a_33515_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=2.44e+12p ps=2.288e+07u w=1e+06u l=150000u M=8
X14120 VSS a_1761_6031# a_1775_5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14121 a_11711_20725# a_7644_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14122 a_9963_54447# a_4128_64391# a_10117_54697# VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14123 vcm a_18162_9492# a_21174_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14124 VDD VSS a_44174_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14125 a_35534_72234# VDD a_35138_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14126 a_21082_20942# pmat.row_n[12] a_21574_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14127 a_45270_23548# a_18546_23546# a_45178_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14128 VSS a_9545_66567# a_11057_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X14129 a_21082_16926# a_18162_16520# a_21174_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1413 a_35230_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14130 vcm a_18162_20536# a_42258_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14131 VDD pmat.rowon_n[9] a_27106_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14132 a_24586_62516# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14133 vcm a_18162_10496# a_38242_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14134 a_48586_71230# pmat.rowon_n[15] a_48190_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14135 VSS a_9195_60039# a_7457_62037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X14136 a_31214_9492# a_18546_9490# a_31122_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14137 a_30121_31849# a_28704_29568# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X14138 a_44570_10862# nmat.rowon_n[13] a_44174_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14139 VSS a_3173_25045# a_3107_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1414 a_10207_30511# a_9761_30511# a_10111_30511# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X14140 VSS ANTENNA__1190__A2.DIODE a_83166_10703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X14141 a_2847_20479# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14142 a_2375_16532# a_2467_16341# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X14143 a_27502_20902# pmat.rowoff_n[12] a_27106_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14144 a_25628_35077# a_24565_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X14145 a_12795_17999# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X14146 a_25505_51183# a_15667_27239# a_25287_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14147 VSS a_14839_20871# a_14839_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14148 a_22482_69222# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14149 a_44561_52815# ANTENNA__1190__B1.DIODE pmat.col_n[25] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1415 a_40349_40726# a_39469_43493# a_40591_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X14150 a_46386_33231# a_45829_35407# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X14151 a_18546_15514# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14152 VDD a_13837_36893# a_13443_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14153 a_3884_55311# a_2727_58470# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14154 a_17113_41317# a_13503_43421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X14155 a_50198_15922# pmat.row_n[7] a_50690_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14156 a_2764_45577# a_1849_45205# a_2417_45173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X14157 a_47278_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14158 a_12543_40541# a_12289_40214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14159 a_34277_37462# a_33765_38053# a_34828_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1416 a_34134_55126# a_18162_55166# a_34226_55126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14160 a_4613_19087# a_4135_19391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14161 a_5323_71829# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X14162 a_23090_58138# a_18162_58178# a_23182_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14163 vcm a_18162_21540# a_19166_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14164 a_37146_71190# a_18162_71230# a_37238_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14165 a_14830_63151# a_10055_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X14166 VSS pmat.row_n[10] a_39550_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14167 VSS a_14825_50095# a_15210_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14168 a_43566_16886# nmat.rowon_n[7] a_43170_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14169 VSS a_25695_28111# a_36637_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1417 a_10383_75637# a_10515_75895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14170 a_26498_68218# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14171 VDD a_23055_41781# a_22879_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14172 a_28872_29673# a_28812_29575# a_28770_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5e+11p pd=2.5e+06u as=0p ps=0u w=1e+06u l=150000u
X14173 a_19928_37253# a_18769_36965# a_19832_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14174 a_6796_15279# a_6679_15492# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X14175 VSS a_16045_37692# a_15737_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14176 a_11202_55687# a_14163_55295# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14177 a_23090_17930# pmat.row_n[9] a_23582_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14178 a_6551_22057# nmat.sw a_6469_21813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14179 a_47236_45743# a_47147_44655# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X1418 VDD a_38627_50613# a_38575_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14180 VDD nmat.rowon_n[5] a_30118_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14181 a_33255_43777# a_24833_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14182 vcm a_18162_67214# a_44266_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14183 VSS a_11149_40188# a_24895_43957# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14184 a_44266_55126# a_18546_55168# a_44174_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14185 VDD a_9135_22057# a_8197_20871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14186 a_2007_49770# a_2099_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X14187 VSS a_2411_16101# a_3657_19453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14188 a_35084_31599# a_33869_31599# a_34895_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14189 a_44666_59504# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1419 VSS a_1858_25615# a_20217_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14190 nmat.rowoff_n[14] a_14839_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X14191 VSS pmat.row_n[2] a_20474_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14192 VSS a_10595_53361# a_10541_53387# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14193 a_2319_31836# a_2124_31867# a_2629_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X14194 VDD a_10851_30485# a_10838_30877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14195 a_29510_59182# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14196 VDD a_12128_32375# a_11299_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14197 a_31122_69182# a_18162_69222# a_31214_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14198 VSS pmat.row_n[1] a_33526_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14199 a_30641_44743# a_30913_44219# a_32035_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X142 VSS a_12248_42583# a_12061_42325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1420 a_21082_15922# pmat.row_n[7] a_21574_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14200 a_45808_45993# a_31675_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14201 a_2559_46261# a_2347_46070# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14202 VDD pmat.rowon_n[14] a_35138_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14203 a_27106_16926# pmat.row_n[8] a_27598_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14204 a_21082_9898# a_18162_9492# a_21174_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14205 a_21174_67174# a_18546_67216# a_21082_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14206 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14207 a_39550_7850# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14208 a_35230_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14209 a_34226_66170# a_18546_66212# a_34134_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1421 a_47582_12870# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14210 a_18162_70226# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14211 VDD pmat.rowon_n[3] a_21082_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14212 a_19955_32521# a_19439_32149# a_19860_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X14213 a_31214_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14214 a_37864_42693# a_36801_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X14215 a_5266_17143# a_6621_16885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14216 VSS VDD a_49590_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14217 VSS a_40951_31599# a_45705_33551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14218 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14219 a_46978_44905# a_7109_29423# a_46896_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1422 VSS pmat.row_n[13] a_21478_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14220 vcm a_18162_63198# a_22178_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14221 a_3109_52093# a_1923_53055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14222 a_2369_26159# a_2325_26401# a_2203_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X14223 vcm a_18162_18528# a_39246_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14224 a_22086_67174# pmat.row_n[11] a_22578_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14225 a_43262_16520# a_18546_16518# a_43170_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14226 vcm a_18162_13508# a_40250_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14227 VSS a_22199_30287# a_29272_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X14228 vcm a_18162_62194# a_35230_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14229 a_35138_66170# pmat.row_n[10] a_35630_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1423 a_24490_24918# VSS a_24094_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14230 a_6920_46287# a_3339_70759# a_5935_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.55e+11p pd=2.51e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X14231 a_46578_64202# pmat.rowon_n[8] a_46182_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14232 VDD a_5227_13077# a_5166_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X14233 a_28631_44265# a_27789_44743# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X14234 a_13529_39429# a_13837_39069# a_13503_39069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14235 a_2007_76970# a_2099_76725# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X14236 a_22482_22910# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14237 a_47278_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14238 a_1979_9334# a_1949_9308# a_1907_9334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14239 a_19074_21946# a_18162_21540# a_19166_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1424 a_18162_20536# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14240 a_2673_52093# a_2195_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14241 a_2347_46070# a_2389_45859# a_2347_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14242 a_36538_56170# pmat.rowon_n[0] a_36142_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14243 a_2319_54965# a_2163_55233# a_2464_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X14244 VSS a_14427_46519# a_14379_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X14245 a_47582_72234# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14246 VSS pmat.row_n[14] a_51598_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14247 a_29206_17524# a_18546_17522# a_29114_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14248 a_41422_49871# a_37820_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14249 a_5671_40097# a_4955_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1425 VSS pmat.row_n[2] a_51598_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14250 a_8859_22467# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14251 a_41558_9858# nmat.rowon_n[14] a_41162_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14252 a_26498_21906# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14253 a_22787_34165# a_22963_34165# a_22915_34191# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X14254 vcm a_18162_24552# a_21174_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14255 VSS pmat.row_n[6] a_41558_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14256 a_29114_57134# pmat.row_n[1] a_29606_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14257 a_38242_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14258 VSS VDD a_24490_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14259 a_33622_55488# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1426 a_24586_57496# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14260 vcm a_18162_23548# a_34226_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14261 a_20570_58500# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14262 nmat.col_n[7] a_14458_4399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14263 VDD a_12429_62607# a_12985_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X14264 a_40707_48783# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X14265 a_42258_71190# a_18546_71232# a_42166_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14266 a_34226_11500# a_18546_11498# a_34134_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14267 VSS pmat.row_n[3] a_20474_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14268 VDD VSS a_42166_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14269 a_29510_12870# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1427 a_8547_65161# a_8031_64789# a_8452_65149# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X14270 a_14504_37607# a_14712_37429# a_14646_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14271 VSS pmat.row_n[2] a_33526_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14272 VDD ANTENNA__1195__A1.DIODE a_47861_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X14273 VSS a_7373_48695# a_5411_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14274 a_11142_64783# a_10707_64783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X14275 a_50198_7890# a_18162_7484# a_50290_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14276 a_1857_47375# a_1769_13103# a_1775_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14277 a_31518_61190# pmat.rowon_n[5] a_31122_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14278 a_39496_30199# a_38905_28853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14279 a_46274_70186# a_18546_70228# a_46182_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1428 VSS a_18568_51959# a_18199_52789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X14280 VDD a_11067_16359# a_14287_57280# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14281 a_39154_22950# pmat.row_n[14] a_39646_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14282 a_43170_71190# pmat.row_n[15] a_43662_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14283 a_26102_7890# a_18162_7484# a_26194_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14284 a_43662_20504# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14285 VSS a_10814_29111# a_10609_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14286 VDD VDD a_50198_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14287 a_43262_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14288 VSS a_16800_47213# a_17012_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14289 a_6788_5853# a_6574_5853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1429 a_39125_48437# a_38907_48841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X14290 VDD pmat.rowon_n[6] a_46182_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14291 a_11113_39747# a_33489_44219# a_34611_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X14292 a_46182_64162# a_18162_64202# a_46274_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14293 a_16837_36603# a_13779_36595# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X14294 a_50290_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14295 a_32218_59142# a_18546_59184# a_32126_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14296 a_28506_18894# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14297 VDD a_29051_37607# a_13357_37429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X14298 a_26515_43447# a_25393_43493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X14299 a_9919_57863# a_10191_57691# a_10149_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X143 a_47278_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1430 vcm a_18162_7484# a_47278_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14300 a_33222_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14301 a_19166_72194# a_18546_72236# a_19074_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14302 VSS pmat.row_n[8] a_32522_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14303 VDD a_11021_43011# a_20752_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X14304 VSS a_13805_43990# a_15107_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X14305 a_10789_64783# a_10601_65103# a_10707_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14306 a_37238_22544# a_18546_22542# a_37146_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14307 a_47186_70186# pmat.row_n[14] a_47678_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14308 VDD nmat.rowon_n[9] a_49194_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14309 VDD pmat.rowoff_n[12] a_20078_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1431 a_34134_14918# pmat.row_n[6] a_34626_14480# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14310 VSS a_5495_65479# a_5275_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14311 a_44174_12910# a_18162_12504# a_44266_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14312 a_23182_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14313 a_45287_33231# a_30663_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.195e+12p pd=1.039e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X14314 a_20078_61150# a_18162_61190# a_20170_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14315 VSS a_2676_29941# a_2610_30345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X14316 VSS pmat.row_n[13] a_44570_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14317 vcm a_18162_55166# a_33222_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14318 a_33130_59142# pmat.row_n[3] a_33622_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14319 VDD a_21981_34191# a_28867_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1432 VSS pmat.row_n[12] a_34530_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14320 a_7970_27907# a_2952_25045# a_7888_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14321 a_21082_24958# a_18162_24552# a_21174_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14322 VDD a_7631_15253# a_4976_16091# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X14323 a_11212_14191# a_10593_15823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14324 a_24586_70548# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14325 a_10873_40693# a_30403_40747# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14326 a_21174_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14327 a_21478_69222# pmat.rowon_n[13] a_21082_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14328 VDD a_1923_61759# a_2464_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14329 a_24094_60146# a_18162_60186# a_24186_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1433 a_4341_24643# a_3325_23439# a_4259_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14330 VSS pmat.row_n[12] a_48586_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14331 a_45574_65206# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14332 a_17740_31287# nmat.en_bit_n[0] a_17882_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14333 VSS a_7263_42453# a_7197_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14334 a_34226_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14335 a_43170_18934# a_18162_18528# a_43262_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14336 a_4591_28335# a_4075_28335# a_4496_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X14337 a_11347_40541# a_11093_40214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14338 a_2203_26159# a_1757_26159# a_2107_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14339 a_11993_10749# a_9675_10396# a_11921_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1434 VSS a_9581_56079# a_11829_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X14340 VDD a_44420_45895# a_41926_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14341 VDD a_11797_60431# a_11977_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14342 VDD nmat.rowon_n[13] a_27106_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14343 VSS a_10291_77269# a_10239_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14344 a_42562_58178# pmat.rowon_n[2] a_42166_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14345 VDD a_9664_47753# a_9839_47679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14346 a_18546_23546# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14347 a_1643_58773# a_1846_59051# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14348 a_10241_54697# a_9581_56079# a_10117_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X14349 a_25494_68218# pmat.rowon_n[12] a_25098_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1435 VSS a_6872_8725# a_6956_8965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14350 VSS pmat.row_n[9] a_22482_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14351 a_45670_61512# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14352 a_48586_56170# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14353 VSS a_2744_25223# a_2191_24501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14354 vcm a_18162_16520# a_32218_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14355 a_50198_66170# a_18162_66210# a_50290_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14356 a_2781_33775# a_1591_33775# a_2672_33775# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X14357 a_39246_69182# a_18546_69224# a_39154_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14358 a_49686_16488# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14359 a_9655_6335# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1436 a_5508_32687# a_5391_32900# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X14360 a_16837_44219# a_15420_44007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X14361 a_1761_4399# a_1591_4399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X14362 a_36634_19500# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14363 a_31518_15882# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14364 VDD a_10049_60663# a_10423_64786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14365 a_22684_35303# a_21621_35515# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X14366 a_13441_70767# a_13327_70741# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14367 a_19399_48437# a_19283_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X14368 a_28506_59182# pmat.rowon_n[3] a_28110_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14369 VDD pmat.rowon_n[5] a_22086_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1437 a_27502_15882# pmat.rowoff_n[7] a_27106_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14370 nmat.rowon_n[7] a_16219_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14371 VDD nmat.rowon_n[7] a_26102_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14372 a_44266_63158# a_18546_63200# a_44174_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14373 a_22269_40391# a_21621_40955# a_22684_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14374 VSS a_15163_32375# a_14839_20871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14375 a_26331_36919# a_25209_36965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14376 VDD a_8583_29199# a_25143_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14377 a_15667_27239# a_41731_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14378 a_44666_67536# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14379 VSS a_8908_14967# a_8767_16055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1438 VSS pmat.row_n[4] a_24490_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14380 VSS a_14336_48071# a_13462_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14381 VSS a_5967_5461# a_5558_9527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14382 VDD a_2215_47375# a_7937_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X14383 VSS a_43315_48437# a_44976_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X14384 a_44174_57134# a_18162_57174# a_44266_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14385 a_20439_27247# a_11927_27399# a_20267_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14386 a_30514_62194# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14387 a_27106_67174# a_18162_67214# a_27198_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14388 VSS VDD a_29510_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14389 a_9581_76207# a_6975_76823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X1439 VDD a_28116_37479# a_28189_37981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X14390 a_20682_32143# a_19605_32149# a_20520_32521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14391 a_20520_30511# a_19439_30511# a_20173_30753# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X14392 VSS pmat.row_n[14] a_44570_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14393 VSS a_10781_42869# a_11200_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14394 a_2467_35015# a_2659_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X14395 VSS a_3295_23060# a_2907_22522# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14396 a_8259_10927# a_8111_11209# a_7896_11079# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X14397 a_3983_49911# a_2983_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14398 a_20170_8488# a_18546_8486# a_20078_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14399 VDD pmat.rowon_n[11] a_21082_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X144 a_28202_64162# a_18546_64204# a_28110_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1440 VSS pmat.row_n[7] a_36538_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14400 VDD pmat.rowon_n[0] a_51202_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14401 comp.adc_nor_latch_0.QN comp_latch VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14402 a_31614_24520# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14403 VSS a_16837_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X14404 a_21174_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14405 a_37542_17890# nmat.rowon_n[6] a_37146_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14406 VSS a_14773_43746# a_13837_43421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X14407 VSS a_6884_74183# a_5931_74183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14408 a_82788_9991# ANTENNA__1184__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14409 a_22915_34191# a_11317_36924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1441 VSS _1196_.B1 nmat.col[30] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X14410 a_21478_64202# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14411 a_34226_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14412 VDD a_8481_10396# a_10047_8751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14413 a_15021_31841# a_14803_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14414 a_21478_22910# nmat.rowon_n[1] a_21082_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14415 VDD a_1899_35051# a_2882_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14416 a_16911_51959# a_17183_51817# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X14417 VSS pmat.row_n[13] a_48586_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14418 a_12815_26409# a_8013_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X14419 a_43262_24552# a_18546_24550# a_43170_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1442 a_9835_15279# a_9485_15279# a_9740_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X14420 VSS a_34277_37462# a_33341_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X14421 vcm a_18162_21540# a_40250_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14422 vcm a_18162_70226# a_35230_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14423 a_39246_14512# a_18546_14510# a_39154_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14424 a_6608_60663# a_6816_60699# a_6750_60797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14425 a_38242_56130# a_18546_56172# a_38150_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14426 a_14833_29967# a_14365_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14427 a_46578_72234# VDD a_46182_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14428 a_25691_52521# ANTENNA__1190__B1.DIODE a_25473_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14429 VDD a_24270_49783# a_23971_50228# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1443 VDD a_28901_48437# a_28573_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=2
X14430 a_32126_20942# pmat.row_n[12] a_32618_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14431 a_32126_16926# a_18162_16520# a_32218_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14432 VDD pmat.rowon_n[2] a_42166_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14433 VDD vcm.sky130_fd_sc_hd__inv_1_4.Y vcm.sky130_fd_sc_hd__nand2_1_1.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14434 VSS pmat.row_n[5] a_38546_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14435 VDD a_12228_40693# a_27566_43805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14436 a_4031_40455# a_2839_38101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14437 a_42562_11866# nmat.rowon_n[12] a_42166_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14438 a_43261_51727# a_16311_28327# pmat.col[24] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X14439 a_25590_15484# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1444 a_13896_8585# a_12981_8213# a_13549_8181# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X14440 a_25494_21906# nmat.rowon_n[2] a_25098_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14441 a_22086_12910# pmat.row_n[4] a_22578_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14442 a_7001_13103# a_5173_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14443 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14444 VDD pmat.rowon_n[1] a_28110_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14445 a_31879_34191# a_31702_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14446 VSS a_1586_50247# a_5639_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14447 a_7004_65871# a_5595_65301# a_6749_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14448 VDD a_4124_28023# a_2283_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14449 VDD a_11271_73085# a_11232_73211# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1445 a_5043_57399# a_4025_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X14450 result_out[5] a_1644_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14451 a_17113_34789# a_15144_36165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X14452 a_37754_30838# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X14453 a_18272_35077# a_17113_34789# a_18176_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14454 a_50594_59182# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14455 a_24895_37429# a_13357_37429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14456 VDD a_7129_57685# a_7159_58038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14457 a_12895_53359# a_9581_56079# a_12806_53359# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14458 a_33526_69222# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14459 a_6330_18909# a_5253_18543# a_6168_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1446 vcm a_18162_24552# a_29206_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14460 VSS a_13697_47349# a_12604_47080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14461 a_8547_77129# a_8197_76757# a_8452_77117# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X14462 a_28506_12870# pmat.rowoff_n[4] a_28110_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14463 VSS pmat.row_n[4] a_37542_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14464 a_26102_11906# pmat.row_n[3] a_26594_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14465 a_17739_50871# a_16083_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X14466 a_9195_7423# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14467 VSS pmat.row_n[11] a_37542_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14468 a_20170_62154# a_18546_62196# a_20078_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14469 a_5612_9295# a_5558_9527# a_5510_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1447 VSS pmat.row_n[6] a_49590_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14470 a_7939_31591# a_31263_32117# a_31221_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14471 a_41321_30511# a_40967_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14472 a_20570_66532# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14473 VSS a_30111_47911# a_45432_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X14474 a_48190_71190# a_18162_71230# a_48282_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14475 VDD pmat.rowon_n[3] a_19074_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14476 VSS a_2683_22089# a_7665_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X14477 VSS a_11852_49783# a_11803_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14478 a_27603_34191# cgen.dlycontrol2_in[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14479 a_33222_61150# a_18546_61192# a_33130_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1448 VSS a_11421_17455# a_11711_16911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14480 a_28049_50613# a_28131_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14481 a_10693_24233# a_5991_23983# a_10597_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14482 vcm a_18162_68218# a_42258_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14483 VDD nmat.rowon_n[1] a_38150_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14484 vcm a_18162_58178# a_38242_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14485 a_37146_8894# pmat.row_n[0] a_37638_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14486 a_10953_38341# a_11261_37981# a_10927_37981# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14487 a_3885_77129# a_2695_76757# a_3776_77129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X14488 VSS a_8305_20871# a_11903_20969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14489 a_5547_24233# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X1449 a_51294_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14490 a_5081_53135# a_2315_44124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X14491 VSS a_3576_17143# a_6795_18319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X14492 a_42258_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14493 a_11235_26159# a_10791_26409# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14494 a_43566_8854# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14495 a_47678_8456# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14496 VSS a_11007_58229# a_10090_58093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14497 a_21082_62154# pmat.row_n[6] a_21574_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14498 VSS pmat.row_n[2] a_31518_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14499 VSS pmat.row_n[15] a_45574_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X145 vcm a_18162_61190# a_25190_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1450 a_37238_72194# a_18546_72236# a_37146_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14500 VDD a_7717_14735# a_13275_48783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X14501 a_34134_61150# pmat.row_n[5] a_34626_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14502 VDD a_11697_56775# a_8749_57141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X14503 a_43262_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14504 a_19470_8854# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14505 a_40158_21946# a_18162_21540# a_40250_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14506 a_2926_45199# a_1849_45205# a_2764_45577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14507 a_8471_56079# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14508 VDD pmat.rowon_n[14] a_46182_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14509 vcm a_18162_69222# a_28202_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1451 a_14369_11177# a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=0p ps=0u w=1e+06u l=150000u
X14510 a_39246_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14511 a_8105_7125# a_7939_7125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X14512 a_32218_67174# a_18546_67216# a_32126_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14513 a_25098_19938# pmat.row_n[11] a_25590_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14514 a_4514_34451# a_4831_34561# a_4789_34685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14515 a_46274_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14516 a_14645_28381# a_10589_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14517 VSS pmat.row_n[0] a_29510_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14518 a_22343_50613# a_22475_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14519 VSS a_20616_27791# a_27355_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1452 VDD a_2847_8511# a_2834_8207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14520 VDD a_11487_69653# a_11391_69831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14521 a_29206_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14522 a_22482_71230# pmat.rowon_n[15] a_22086_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14523 a_2325_63669# a_2107_64073# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X14524 a_28202_12504# a_18546_12502# a_28110_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14525 a_19860_30511# a_9307_31068# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14526 VSS a_21147_49525# pmat.row_n[13] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X14527 a_10864_68565# a_10391_69653# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14528 a_6823_58951# a_6559_57167# a_7168_58799# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X14529 vcm a_18162_19532# a_37238_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1453 a_45193_50639# a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14530 a_44174_20942# a_18162_20536# a_44266_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14531 a_11397_76457# a_11023_76359# a_11325_76457# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14532 a_50198_57134# pmat.row_n[1] a_50690_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14533 a_19166_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14534 a_40250_59142# a_18546_59184# a_40158_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14535 vcm a_18162_63198# a_33222_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14536 a_33130_67174# pmat.row_n[11] a_33622_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14537 a_36538_18894# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14538 VSS a_22725_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X14539 VSS pmat.row_n[8] a_40554_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1454 a_13239_65161# a_12723_64789# a_13144_65149# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X14540 a_25139_27497# _1192_.A2 a_24921_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14541 a_18162_67214# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X14542 a_49590_17890# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14543 a_20474_23914# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14544 VSS a_5497_62839# a_5445_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X14545 cgen.enable_dlycontrol_in a_1591_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X14546 a_50594_12870# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14547 a_21174_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14548 a_33526_22910# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14549 vcm a_18162_55166# a_41254_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1455 a_28602_58500# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14550 a_3909_17209# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14551 a_27198_18528# a_18546_18526# a_27106_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14552 a_41162_59142# pmat.row_n[3] a_41654_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14553 VDD nmat.rowon_n[15] a_32126_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14554 VSS a_1858_25615# a_2511_34319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X14555 a_29510_61190# pmat.rowon_n[5] a_29114_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14556 VSS pmat.row_n[9] a_26498_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14557 VDD a_45119_32661# a_45396_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.195e+12p ps=1.039e+07u w=1e+06u l=150000u M=2
X14558 a_1895_38842# a_2283_39189# a_2241_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14559 a_30514_15882# pmat.rowoff_n[7] a_30118_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1456 VSS a_11927_27399# a_20439_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X14560 a_37007_52521# a_34942_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14561 a_7799_16367# a_4976_16091# a_7436_16519# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X14562 a_5462_30006# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X14563 a_36234_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14564 VSS a_10190_60663# a_10191_57691# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14565 nmat.rowoff_n[11] a_10515_61839# a_14370_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X14566 vcm a_18162_24552# a_32218_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14567 a_16552_46805# a_16403_46831# a_16848_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14568 vcm a_18162_66210# a_31214_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14569 a_9747_69679# a_9301_69679# a_9651_69679# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X1457 a_22377_51727# _1194_.A2 pmat.col_n[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X14570 a_5253_32687# a_5087_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X14571 vcm a_18162_14512# a_28202_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14572 a_49286_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14573 vcm a_18162_56170# a_27198_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14574 VDD a_2500_30345# a_2676_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14575 a_13427_18303# a_13252_18377# a_13606_18365# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X14576 VDD a_24719_35253# a_11921_35286# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14577 a_31614_58500# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14578 a_27502_13874# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14579 a_12561_57167# a_6927_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1458 a_1757_36501# a_1591_36501# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14580 VSS a_38531_51348# pmat.col[19] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14581 VSS pmat.row_n[3] a_31518_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14582 a_10388_17277# a_8305_20871# a_10167_16950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X14583 VSS a_4031_20884# a_3183_19258# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14584 a_33386_30485# a_6664_26159# a_33601_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14585 a_28202_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14586 VSS a_7563_63303# a_7796_62723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14587 a_39246_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14588 VSS a_29685_34954# a_20534_35431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14589 VDD a_44444_32233# a_46897_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1459 VDD a_6643_5724# a_6574_5853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14590 a_30118_8894# a_18162_8488# a_30210_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14591 a_13529_38341# a_13837_37981# a_13503_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14592 a_39550_66210# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14593 VDD a_3879_42997# a_2263_43719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X14594 a_7937_61839# a_5784_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14595 VSS pmat.row_n[8] a_43566_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14596 a_37146_23954# pmat.row_n[15] a_37638_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14597 a_36459_29673# a_36453_29199# a_36895_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14598 a_37146_19938# a_18162_19532# a_37238_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14599 a_22276_46831# a_21797_47081# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X146 VSS a_7693_22365# a_11897_21813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X1460 a_44174_9898# pmat.row_n[1] a_44666_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14600 a_41654_21508# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14601 a_41254_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14602 a_44174_65166# a_18162_65206# a_44266_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14603 pmat.col_n[18] a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14604 VSS a_28281_41245# a_27973_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14605 VSS a_13837_43421# a_13529_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14606 a_2356_13647# a_1687_13621# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14607 nmat.col[1] _1196_.B1 a_13283_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14608 a_21970_48071# a_19283_49783# a_22273_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14609 a_3814_65871# a_3727_66113# a_3410_66003# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X1461 VSS pmat.row_n[3] a_28506_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14610 VSS pmat.row_n[7] a_29510_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14611 VSS a_7436_16519# a_7387_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14612 VDD nmat.rowon_n[7] a_34134_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14613 a_19470_69222# pmat.rowon_n[13] a_19074_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14614 a_2781_50095# a_1591_50095# a_2672_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X14615 a_15543_31573# a_15368_31599# a_15722_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X14616 VSS a_10811_77437# a_10772_77563# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14617 vcm a_18162_17524# a_26194_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14618 a_20474_64202# pmat.rowon_n[8] a_20078_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14619 a_1846_69931# a_2163_69821# a_2121_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1462 a_41254_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14620 a_30210_15516# a_18546_15514# a_30118_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14621 a_4737_23957# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14622 VDD pmat.rowoff_n[7] a_47186_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14623 a_14287_12015# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14624 a_44666_12472# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14625 a_4446_65871# a_3727_66113# a_3883_65845# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X14626 VDD a_2683_22089# a_9201_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14627 a_12925_60431# a_9135_60967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X14628 a_2464_56989# a_2250_56989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14629 a_42166_13914# a_18162_13508# a_42258_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1463 VSS a_30571_50959# a_46815_37013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.9975e+11p ps=3.83e+06u w=650000u l=150000u
X14630 VSS a_2683_22089# a_8951_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14631 a_18162_20536# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X14632 a_21174_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14633 a_27598_22512# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14634 a_35786_47893# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14635 a_9195_58951# a_1769_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14636 VDD pmat.rowoff_n[12] a_31122_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14637 a_37820_30485# a_40125_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u M=2
X14638 VDD a_24374_29941# a_28803_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X14639 a_10449_53153# a_6559_33767# a_10363_53153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1464 a_9759_62607# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X14640 a_21478_72234# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14641 a_34226_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14642 a_23821_35279# a_23655_35279# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14643 a_51598_61190# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14644 a_5715_16911# a_5463_17027# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14645 VDD a_11435_58791# a_14287_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14646 a_34530_71230# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14647 a_8471_56079# a_7847_56085# a_8363_56457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14648 vcm a_18162_11500# a_31214_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14649 a_18162_18528# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X1465 a_12243_16733# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X14650 VDD pmat.rowoff_n[4] a_21082_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14651 a_38242_64162# a_18546_64204# a_38150_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14652 a_48682_11468# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14653 a_38642_68540# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14654 a_43495_47919# a_43261_48783# a_43132_48071# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X14655 a_3026_23805# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14656 a_32126_24958# a_18162_24552# a_32218_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14657 nmat.col[10] _1187_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=0p ps=0u w=650000u l=150000u M=2
X14658 VDD pmat.rowon_n[10] a_42166_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14659 a_28110_14918# a_18162_14512# a_28202_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1466 a_45187_38129# a_46815_37013# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14660 a_6661_21583# a_3351_27249# a_6579_21583# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14661 VDD a_18241_31698# a_34243_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14662 a_32218_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14663 a_4779_30511# a_4333_30511# a_4683_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14664 VDD a_33617_42333# a_33223_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14665 a_35138_60146# a_18162_60186# a_35230_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14666 VDD a_20520_30511# a_20695_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14667 VDD a_78448_40202# a_78261_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14668 a_25190_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14669 a_44763_34293# a_44647_35520# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1467 a_26498_62194# pmat.rowon_n[6] a_26102_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14670 a_5989_40303# a_5823_40303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X14671 VDD nmat.rowon_n[12] a_25098_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14672 vcm a_18162_60186# a_39246_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14673 vcm a_18162_7484# a_32218_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14674 a_26583_34343# cgen.dlycontrol1_in[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14675 a_6607_75895# a_6051_74183# a_7005_75983# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X14676 a_39154_64162# pmat.row_n[8] a_39646_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14677 a_43662_62516# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14678 VDD a_9581_73487# a_9685_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14679 a_13005_66665# a_12217_66389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1468 a_41558_71230# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14680 a_2319_67740# a_2163_67645# a_2464_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X14681 nmat.rowoff_n[5] a_10515_61839# a_14277_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X14682 a_8439_10422# a_8257_10422# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14683 VSS a_7840_27247# a_19697_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14684 VDD a_11759_10615# a_11051_8903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14685 a_20170_70186# a_18546_70228# a_20078_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14686 a_47678_19500# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14687 a_20253_46287# a_20076_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14688 vcm a_18162_71230# a_29206_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14689 VDD pmat.rowon_n[11] a_19074_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1469 VSS a_6787_47607# a_12081_62723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X14690 VDD nmat.rowon_n[14] a_41162_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14691 VDD pmat.rowon_n[0] a_49194_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14692 VDD pmat.rowon_n[6] a_20078_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14693 a_41558_69222# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14694 VDD _1184_.A2 a_11897_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14695 a_7465_53359# a_6559_33767# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X14696 VSS a_3688_17179# a_9820_18115# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14697 VSS a_43132_48071# a_42292_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14698 a_29606_63520# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14699 a_20961_30305# a_20895_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X147 a_7259_31433# a_6909_31061# a_7164_31421# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1470 pmat.rowon_n[3] a_10239_14183# a_14471_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X14700 VDD pmat.rowon_n[5] a_33130_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14701 VSS a_4675_54599# a_3199_53877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14702 a_10589_22351# a_10209_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X14703 a_5156_14025# a_4241_13653# a_4809_13621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X14704 a_19470_22910# nmat.rowon_n[1] a_19074_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14705 a_21082_70186# pmat.row_n[14] a_21574_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14706 a_42166_58138# a_18162_58178# a_42258_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14707 a_25098_68178# a_18162_68218# a_25190_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14708 a_13285_70767# a_12809_69679# a_13203_70767# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14709 a_12862_16733# a_11785_16367# a_12700_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1471 a_38150_72194# VDD a_38642_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14710 VDD a_4025_54965# a_4535_56623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14711 a_2610_30345# a_2217_29973# a_2500_30345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X14712 VSS a_39505_38780# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X14713 a_42166_17930# pmat.row_n[9] a_42658_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14714 VSS pmat.row_n[15] a_42562_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14715 a_31122_11906# a_18162_11500# a_31214_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14716 a_39246_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14717 a_4461_46805# a_4128_46983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14718 a_12517_51183# a_11807_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14719 VDD a_31263_28309# a_31015_29111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.25e+11p ps=2.85e+06u w=1e+06u l=150000u
X1472 a_4032_26311# a_2952_25045# a_4174_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14720 VSS a_77882_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_4.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14721 VDD a_2417_45173# a_2307_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14722 a_35534_18894# nmat.rowon_n[5] a_35138_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14723 a_28110_59142# a_18162_59182# a_28202_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14724 a_29768_39429# a_28705_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14725 a_11877_58261# a_11711_58261# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14726 a_32218_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14727 a_28202_20536# a_18546_20534# a_28110_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14728 VSS a_2411_43301# a_8625_56445# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14729 a_17559_51157# a_17033_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X1473 a_19332_41959# a_19428_41781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14730 a_48586_17890# nmat.rowon_n[6] a_48190_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14731 vcm a_18162_69222# a_36234_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14732 a_46182_16926# pmat.row_n[8] a_46674_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14733 a_39550_8854# nmat.rowon_n[15] a_39154_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14734 a_12581_69455# a_12067_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14735 a_51598_8854# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14736 a_40250_67174# a_18546_67216# a_40158_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14737 a_9871_53903# a_4128_64391# a_9953_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14738 a_32522_64202# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14739 a_23329_37462# a_22725_38053# a_23847_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1474 a_38642_21508# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14740 a_5597_44807# a_5921_44629# a_5843_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X14741 a_36234_57134# a_18546_57176# a_36142_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14742 VDD comp_latch a_55914_40254# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14743 a_30118_21946# pmat.row_n[13] a_30610_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14744 a_45815_36815# a_43776_30287# a_45625_36495# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X14745 a_30118_17930# a_18162_17524# a_30210_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14746 a_5785_48463# a_5383_48783# a_5621_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X14747 VDD a_6179_65479# a_5495_65479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X14748 VDD pmat.rowon_n[3] a_40158_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14749 a_37612_30663# a_37827_30793# a_37754_30838# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X1475 vcm a_18162_10496# a_51294_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14750 VSS pmat.row_n[6] a_36538_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14751 VSS a_7693_22365# a_10932_21959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X14752 a_49286_56130# a_18546_56172# a_49194_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14753 a_33331_31599# a_32771_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14754 a_11798_62063# a_10049_60663# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14755 a_2672_64073# a_1757_63701# a_2325_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14756 a_6794_64015# a_5081_53135# a_6984_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14757 VSS pmat.row_n[3] a_25494_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14758 a_22482_56170# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14759 a_19074_18934# pmat.row_n[10] a_19566_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1476 a_38242_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14760 VSS VDD a_19470_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14761 a_10570_62973# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14762 a_6615_37039# a_6265_37039# a_6520_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X14763 VSS a_28525_43655# a_28907_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X14764 VSS a_12197_38306# a_11261_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X14765 a_20078_13914# pmat.row_n[5] a_20570_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14766 VSS pmat.row_n[5] a_49590_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14767 a_23582_16488# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14768 VSS a_14336_46983# a_13830_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14769 result_out[1] a_1644_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1477 a_42658_70548# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14770 a_7631_55687# a_1769_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14771 a_3746_58487# a_4043_33535# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X14772 VSS a_12069_38517# a_16339_43745# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14773 a_5907_23145# a_3351_27249# a_5825_22901# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14774 vcm a_18162_63198# a_41254_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14775 a_8038_11254# a_1717_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14776 a_41162_67174# pmat.row_n[11] a_41654_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14777 a_33130_12910# pmat.row_n[4] a_33622_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14778 a_3331_59317# a_3136_59459# a_3641_59709# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X14779 a_3434_51727# a_2715_51969# a_2871_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1478 a_12038_55687# a_10955_55687# a_12175_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14780 a_5633_71631# a_5779_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14781 VSS a_10697_75218# a_11905_74895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14782 VSS nmat.sample a_18546_8486# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X14783 a_4175_49667# a_3983_49911# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14784 a_40677_48437# a_40949_48437# a_41348_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X14785 a_14071_8511# a_13896_8585# a_14250_8573# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X14786 a_26498_55166# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14787 a_26498_13874# nmat.rowon_n[10] a_26102_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14788 VDD a_4984_41935# a_5558_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14789 VSS a_40467_46261# a_11948_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1479 a_34611_43177# a_34553_42658# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X14790 a_4357_51433# a_2389_45859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14791 a_36634_7452# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14792 a_6836_24527# a_4523_21276# a_6752_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14793 a_44774_40821# a_46013_42997# a_46043_43343# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u M=2
X14794 a_41558_22910# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14795 a_11337_25071# a_5991_23983# a_11505_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14796 VSS _1224_.X a_82735_2223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X14797 a_35230_18528# a_18546_18526# a_35138_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14798 VDD a_14491_51969# a_14452_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14799 VDD a_30489_36893# a_30095_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X148 a_28602_68540# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1480 VSS a_4259_65103# a_4445_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14800 a_44183_27497# a_27763_27221# a_43965_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14801 vcm a_18162_64202# a_27198_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14802 nmat.col[10] a_10883_3303# a_13546_5263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14803 VSS a_9441_20189# a_10478_25045# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14804 VSS _1183_.A2 a_32740_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14805 VDD VDD a_46182_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14806 VSS VDD a_42562_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14807 a_27020_49007# a_25839_49783# a_25850_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X14808 a_27106_68178# pmat.row_n[12] a_27598_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14809 a_38546_66210# pmat.rowon_n[10] a_38150_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1481 a_11067_64015# a_24775_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X14810 a_31214_62154# a_18546_62196# a_31122_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14811 a_4533_38279# a_7355_37013# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14812 a_40645_46519# a_11067_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.728e+11p pd=1.82e+06u as=0p ps=0u w=640000u l=150000u
X14813 a_31614_66532# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14814 a_48282_17524# a_18546_17522# a_48190_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14815 VDD a_9963_28111# a_15857_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14816 VDD pmat.rowoff_n[15] a_36142_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14817 a_23883_34165# a_11057_35836# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14818 VDD a_5749_57685# a_5779_58038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14819 a_31122_56130# a_18162_56170# a_31214_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1482 VSS a_11711_50959# a_38601_49035# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14820 a_13459_28111# a_41731_49525# a_46487_49871# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14821 a_34134_7890# VDD a_34626_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14822 a_22523_31094# pmat.en_bit_n[2] a_22064_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14823 a_4149_44431# a_3325_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14824 VDD a_9213_53903# a_9953_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14825 pmat.col[28] ANTENNA__1395__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14826 VDD a_14773_43746# a_13837_43421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X14827 a_23486_9858# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14828 VDD a_9303_22351# a_10097_22895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14829 a_36617_42043# a_34924_41605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X1483 a_10795_47893# a_11230_48171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14830 a_12453_63151# a_11797_60431# a_12381_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14831 vcm a_18162_14512# a_36234_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14832 VDD a_9092_31287# a_7619_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14833 a_28506_7850# VDD a_28110_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14834 VSS VDD a_43566_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14835 a_13483_37782# a_13301_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14836 vcm a_18162_13508# a_49286_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14837 VSS a_12092_42895# a_12198_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14838 a_32126_62154# pmat.row_n[6] a_32618_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14839 a_40250_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1484 a_45270_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14840 a_37238_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14841 a_11435_58791# a_15655_50613# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X14842 a_22064_31287# pmat.en_bit_n[2] a_22206_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14843 VSS a_2847_23743# a_2781_23817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X14844 VSS a_24643_51959# pmat.col_n[3] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14845 a_11165_67753# a_9545_66567# a_10975_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X14846 a_25590_57496# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14847 a_9385_26409# a_4516_21531# a_9313_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14848 a_20474_72234# VDD a_20078_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14849 a_3331_59317# a_3175_59585# a_3476_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X1485 a_42166_60146# a_18162_60186# a_42258_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14850 a_9112_77129# a_8031_76757# a_8765_76725# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14851 a_30210_23548# a_18546_23546# a_30118_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14852 a_50594_61190# pmat.rowon_n[5] a_50198_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14853 a_26194_13508# a_18546_13506# a_26102_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14854 vcm a_18162_10496# a_23182_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14855 VDD a_3793_47479# a_3799_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14856 a_9274_64783# a_8197_64789# a_9112_65161# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14857 a_33526_71230# pmat.rowon_n[15] a_33130_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14858 VSS pmat.row_n[4] a_25494_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14859 vcm a_18162_19532# a_48282_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1486 a_14792_51727# a_14578_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X14860 a_2973_10089# a_2021_9563# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14861 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14862 a_51294_59142# a_18546_59184# a_51202_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14863 a_26041_36374# a_25209_36965# a_26331_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X14864 a_47582_18894# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14865 a_38242_72194# a_18546_72236# a_38150_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14866 a_10233_50639# a_9463_50877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14867 VSS pmat.row_n[8] a_51598_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14868 a_14691_29575# a_14751_28341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X14869 vcm a_18162_9492# a_48282_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1487 VDD a_28525_43655# a_28848_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X14870 a_7937_61519# a_1823_66941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14871 a_17046_52521# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X14872 a_35630_22512# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14873 a_28110_22950# a_18162_22544# a_28202_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14874 VDD pmat.rowon_n[8] a_38150_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14875 a_5320_30199# a_5535_29980# a_5462_30006# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X14876 a_32218_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14877 a_18546_18526# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X14878 VSS a_22085_38550# a_23479_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14879 a_44791_43541# a_7109_29423# a_45009_43817# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1488 a_25098_70186# a_18162_70226# a_25190_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14880 a_7865_58553# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14881 a_9597_53609# a_7521_47081# a_9502_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X14882 a_9415_24233# a_6829_26703# a_9217_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X14883 a_22086_71190# a_18162_71230# a_22178_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14884 a_27502_62194# pmat.rowon_n[6] a_27106_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14885 VSS pmat.row_n[10] a_24490_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14886 a_46130_34319# a_29937_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14887 a_6806_63695# a_4985_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X14888 a_4956_59317# a_5341_59317# a_5085_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X14889 a_39154_72194# VDD a_39646_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1489 a_8215_69929# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14890 VDD a_38711_37683# a_38737_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X14891 a_43662_70548# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14892 a_36142_14918# a_18162_14512# a_36234_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14893 a_11292_36367# a_11041_36596# a_11071_36694# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X14894 VDD a_20173_30753# a_20063_30877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14895 VSS a_10781_42364# a_23055_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14896 a_39646_60508# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14897 a_40250_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14898 a_47278_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14899 a_40554_69222# pmat.rowon_n[13] a_40158_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X149 VDD pmat.rowon_n[10] a_32126_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1490 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14900 vcm a_18162_57174# a_25190_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14901 VDD a_6553_53047# a_5784_52423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14902 a_26102_70186# a_18162_70226# a_26194_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14903 VSS a_1957_43567# a_12277_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X14904 a_27687_34967# cgen.dlycontrol1_in[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14905 VSS a_7865_58553# a_7799_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14906 a_25494_14878# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14907 VDD a_5565_19605# a_5595_19958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14908 a_26833_35073# a_26767_34967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14909 VDD pmat.rowon_n[14] a_20078_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1491 a_3339_59879# a_3891_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X14910 a_29606_71552# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14911 a_37542_67214# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14912 a_6772_62927# a_3866_57399# a_6681_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X14913 a_9303_22351# a_8859_22467# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14914 a_3431_57167# a_3770_57399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14915 VDD pmat.rowoff_n[12] a_29114_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14916 a_20170_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14917 a_44570_68218# pmat.rowon_n[12] a_44174_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14918 VSS pmat.row_n[9] a_41558_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14919 a_11795_26819# a_9777_26935# a_11713_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1492 vcm a_18162_12504# a_24186_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14920 VSS a_9777_26935# a_11713_26819# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X14921 VSS a_22199_30287# a_41600_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X14922 vcm a_18162_16520# a_51294_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14923 VDD nmat.rowon_n[6] a_41162_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14924 a_1642_20871# a_1738_20693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14925 a_39392_28111# ANTENNA__1395__A1.DIODE a_39089_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X14926 VSS a_24937_36039# a_25687_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14927 a_29114_61150# a_18162_61190# a_29206_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14928 VSS a_11067_27239# nmat.col_n[0] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14929 a_1881_71855# a_1846_72107# a_1643_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1493 a_12257_8527# a_12133_9001# a_12269_8207# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14930 a_33222_9492# a_18546_9490# a_33130_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14931 VDD a_47223_38671# _1192_.B1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X14932 VDD a_7563_63303# a_7878_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14933 a_12795_17999# a_12171_18005# a_12687_18377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14934 a_48190_23954# pmat.row_n[15] a_48682_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14935 a_48190_19938# a_18162_19532# a_48282_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14936 VDD pmat.rowoff_n[4] a_19074_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14937 VDD a_18660_47607# a_18083_47593# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X14938 a_7129_57685# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14939 VSS a_10781_42364# a_10725_42390# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1494 VDD a_2021_9563# a_4357_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14940 a_6334_65327# a_5462_62215# a_6524_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14941 a_37828_27247# ANTENNA__1190__A1.DIODE a_37525_27221# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14942 vcm a_18162_18528# a_24186_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14943 a_47582_59182# pmat.rowon_n[3] a_47186_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14944 VSS pmat.row_n[0] a_44570_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14945 a_38150_15922# pmat.row_n[7] a_38642_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14946 a_48190_9898# a_18162_9492# a_48282_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14947 VDD nmat.sw a_10383_13077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14948 VDD nmat.rowon_n[7] a_45178_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14949 a_19865_46983# nmat.rowon_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1495 a_39154_13914# a_18162_13508# a_39246_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14950 a_42658_13476# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14951 VSS pmat.row_n[10] a_27502_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14952 a_31518_64202# pmat.rowon_n[8] a_31122_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14953 VDD a_9545_66567# a_10057_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14954 a_37680_37479# a_37776_37479# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X14955 a_78165_39738# a_78261_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14956 VSS a_2983_48071# a_4167_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X14957 VDD a_12003_52815# a_12723_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14958 a_3241_47919# a_2971_48285# a_3151_48285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14959 a_8213_53877# a_7995_54281# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1496 VDD nmat.rowon_n[13] a_45178_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14960 VDD cgen.enable_dlycontrol_in a_24667_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14961 a_32218_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14962 a_14741_56873# a_10515_15055# a_14657_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14963 a_20411_51157# a_19584_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X14964 a_21478_56170# pmat.rowon_n[0] a_21082_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14965 a_46182_67174# a_18162_67214# a_46274_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14966 VSS VDD a_48586_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14967 a_32522_72234# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14968 a_36234_65166# a_18546_65208# a_36142_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14969 a_36634_69544# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1497 a_18162_65206# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14970 VDD a_1586_33927# a_6099_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14971 a_19970_46287# a_19793_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14972 VSS a_10055_31591# a_17403_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14973 vcm a_18162_71230# a_50290_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14974 VDD pmat.rowon_n[11] a_40158_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14975 VDD a_4075_31591# a_14369_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14976 a_29206_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14977 a_49286_64162# a_18546_64204# a_49194_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14978 a_18546_63200# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X14979 a_36142_59142# a_18162_59182# a_36234_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1498 a_11849_50095# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14980 a_49686_68540# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14981 VSS a_77882_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_2.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14982 a_40250_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14983 a_18546_10494# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14984 a_19074_69182# a_18162_69222# a_19166_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14985 VDD a_2163_61761# a_2124_61635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14986 a_2387_70483# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14987 a_23182_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14988 a_25494_55166# VSS a_25098_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14989 a_40554_22910# nmat.rowon_n[1] a_40158_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1499 VDD pmat.rowoff_n[12] a_28110_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14990 a_37146_65166# pmat.row_n[9] a_37638_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14991 a_13805_43990# a_13985_44581# a_15048_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14992 a_2319_31836# a_2163_31741# a_2464_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X14993 a_22895_47893# a_22459_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X14994 VDD pmat.rowon_n[12] a_26102_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14995 a_51202_20942# pmat.row_n[12] a_51694_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14996 VDD a_1899_35051# a_6641_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14997 a_51202_16926# a_18162_16520# a_51294_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14998 a_26498_63198# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14999 VDD a_5266_17143# a_6835_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15 a_13443_38007# a_13503_37981# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.19408e+15p ps=1.06986e+10u w=800000u l=150000u M=2
X150 VSS a_76962_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_3.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1500 VSS a_1923_69823# a_1881_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15000 a_33222_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15001 VSS a_9075_28023# a_11159_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15002 a_37542_20902# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15003 VSS a_10927_43421# a_10985_44220# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X15004 a_4351_39872# a_3325_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X15005 a_41162_12910# pmat.row_n[4] a_41654_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15006 a_44570_21906# nmat.rowon_n[2] a_44174_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15007 vcm a_18162_72234# a_27198_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15008 VSS a_8264_11703# a_7283_11484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15009 VDD a_10927_37981# a_10953_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1501 a_43566_68218# pmat.rowon_n[12] a_43170_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15010 a_43274_48246# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X15011 a_12764_40541# a_11565_39061# a_12543_40214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X15012 a_31214_70186# a_18546_70228# a_31122_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15013 a_5423_67191# a_5651_66975# a_5597_67297# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15014 VDD pmat.rowon_n[1] a_47186_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15015 a_24094_22950# pmat.row_n[14] a_24586_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15016 a_6244_71829# a_3339_70759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15017 vcm a_18162_22544# a_45270_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15018 a_27198_60146# a_18546_60188# a_27106_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15019 a_27598_64524# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1502 vcm a_18162_16520# a_50290_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15020 a_35353_50639# a_30571_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15021 VSS a_14533_39631# a_19233_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X15022 VSS a_33382_46983# a_31152_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15023 VDD pmat.rowon_n[6] a_31122_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15024 a_34530_13874# nmat.rowon_n[10] a_34134_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15025 a_31122_64162# a_18162_64202# a_31214_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15026 a_12020_39783# a_12228_39605# a_12162_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15027 a_30479_52271# ANTENNA__1184__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15028 a_4503_70455# a_2419_53351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15029 a_47582_12870# pmat.rowoff_n[4] a_47186_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1503 VDD a_1586_50247# a_1591_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15030 a_7953_67753# a_7899_67477# a_7435_68021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15031 a_30100_52047# a_11067_27239# a_29797_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X15032 VSS a_1591_13103# a_1769_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X15033 a_12605_28879# a_10957_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X15034 VDD a_3688_17179# a_9902_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15035 VSS pmat.row_n[14] a_39550_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15036 a_22178_22544# a_18546_22542# a_22086_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15037 a_32126_70186# pmat.row_n[14] a_32618_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15038 vcm a_18162_21540# a_49286_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15039 a_40158_18934# pmat.row_n[10] a_40650_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1504 a_28110_61150# a_18162_61190# a_28202_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15040 a_6829_25731# a_6641_25731# a_6747_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15041 a_2012_43389# a_1895_43194# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15042 a_28110_60146# pmat.row_n[4] a_28602_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15043 a_37238_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15044 a_4697_74005# a_4225_71311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15045 pmat.col_n[13] a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15046 VSS VDD a_50594_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15047 VSS a_3339_59879# a_10529_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15048 a_14963_37782# a_14712_37429# a_14504_37607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15049 a_6404_5853# a_5967_5461# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1505 VDD a_13739_51701# a_13432_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15050 a_43566_9858# nmat.rowon_n[14] a_43170_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15051 a_21867_34709# a_22043_35041# a_21995_35101# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X15052 a_26194_21540# a_18546_21538# a_26102_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15053 a_44266_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15054 a_41049_30511# a_17842_27497# a_40967_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15055 a_10785_30511# a_9595_30511# a_10676_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15056 result_out[6] a_1644_62581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15057 a_46578_18894# nmat.rowon_n[5] a_46182_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15058 VSS pmat.row_n[2] a_50594_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15059 a_10449_32509# a_10070_32143# a_10377_32509# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X1506 nmat.col_n[9] a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15060 VDD a_7865_58553# a_7895_58294# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15061 a_19470_9858# nmat.rowon_n[14] a_19074_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15062 a_17049_48579# a_16800_47213# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X15063 VSS a_4025_54965# a_4535_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15064 VDD a_24747_29967# a_40785_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X15065 a_31518_9858# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15066 a_30955_42689# a_24833_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15067 VDD a_13329_47893# a_12328_48168# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15068 VSS pmat.row_n[12] a_33526_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15069 a_30514_65206# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1507 a_6835_14735# a_7295_14441# a_7085_15055# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.39e+12p pd=1.278e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15070 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15071 a_12875_16341# a_12700_16367# a_13054_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15072 vcm a_18162_69222# a_47278_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15073 a_20520_30511# a_19605_30511# a_20173_30753# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X15074 a_51294_67174# a_18546_67216# a_51202_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15075 a_44174_19938# pmat.row_n[11] a_44666_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15076 VSS a_11823_46973# a_11784_47099# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15077 VDD a_1586_50247# a_12907_54997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15078 a_47278_57134# a_18546_57176# a_47186_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15079 a_9367_14774# a_8305_20871# a_8908_14967# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1508 a_5682_56311# a_12341_57141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15080 a_20474_57174# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15081 a_2557_65327# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15082 a_1959_10615# a_1979_11254# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15083 VDD pmat.rowon_n[3] a_51202_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15084 a_48282_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15085 a_8507_57487# a_4128_64391# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X15086 VSS pmat.row_n[6] a_47582_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15087 VDD a_9583_10121# a_10943_8903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15088 VSS a_7435_68021# a_6970_67191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15089 a_22449_44219# a_21124_42919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X1509 VDD ANTENNA__1195__A1.DIODE a_23849_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X15090 a_29404_44869# a_28245_44581# a_29367_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X15091 a_26102_63158# pmat.row_n[7] a_26594_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15092 a_12155_27791# a_11711_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15093 a_30610_61512# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15094 a_33526_56170# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15095 VDD VDD a_38150_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15096 VSS a_31469_40726# a_32035_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X15097 a_24186_69182# a_18546_69224# a_24094_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15098 a_34626_16488# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15099 VSS a_38851_28327# a_47043_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X151 a_13717_21263# a_5351_19913# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u
X1510 a_33925_29199# a_31339_31787# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.9e+11p pd=3.8e+06u as=0p ps=0u w=650000u l=150000u
X15100 VSS a_12152_66415# a_12809_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15101 a_38242_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15102 a_21574_19500# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15103 a_12559_51325# a_5363_33551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X15104 a_13361_56399# a_13091_54447# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15105 VSS a_24737_30485# a_24160_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15106 VDD a_2839_38101# a_4351_39872# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15107 VSS a_2149_45717# a_2568_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15108 a_6641_43023# a_6554_43255# a_6311_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15109 a_1644_34293# a_1591_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1511 VDD a_22628_30485# a_28803_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15110 a_36142_22950# a_18162_22544# a_36234_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15111 a_11813_8751# a_11051_8903# a_11731_8751# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15112 VDD a_25287_32117# a_6007_33767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15113 a_40250_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15114 a_28202_68178# a_18546_68220# a_28110_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15115 a_4031_20884# a_4123_20693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15116 VSS a_12345_39100# a_12289_39126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15117 vcm a_18162_65206# a_25190_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15118 a_46994_34639# a_46522_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X15119 VSS pmat.row_n[0] a_22482_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1512 vcm a_18162_71230# a_36234_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15120 VDD nmat.rowon_n[15] a_26102_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15121 VDD a_14149_39747# a_20337_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15122 a_25098_69182# pmat.row_n[13] a_25590_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15123 a_49194_21946# a_18162_21540# a_49286_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15124 a_2592_29423# a_1781_9308# a_2289_29397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X15125 a_36538_67214# pmat.rowon_n[11] a_36142_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15126 a_2250_56989# a_2163_56765# a_1846_56875# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15127 vcm a_18162_15516# a_43262_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15128 a_46274_18528# a_18546_18526# a_46182_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15129 a_6832_67279# a_5779_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X1513 a_7797_63151# a_7321_63151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.34e+11p pd=2.02e+06u as=0p ps=0u w=650000u l=150000u
X15130 VSS pmat.row_n[9] a_45574_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15131 a_7413_63151# a_7563_63303# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15132 a_12132_12925# a_10845_12559# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15133 a_1979_11254# a_2021_11043# a_1979_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15134 VSS a_1899_35051# a_2882_74397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X15135 a_2882_61519# a_2163_61761# a_2319_61493# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X15136 a_26194_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15137 a_13205_62607# a_12429_62607# a_5462_62215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15138 VSS a_2021_11043# a_7009_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15139 vcm a_18162_24552# a_51294_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1514 VSS a_8583_29199# a_25481_29245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15140 VDD a_4308_24135# a_3387_22869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15141 vcm a_18162_14512# a_47278_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15142 a_38071_30838# a_37820_30485# a_37612_30663# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15143 VSS a_14933_37429# a_14867_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15144 vcm a_18162_56170# a_46274_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15145 a_13985_41317# a_10651_42035# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X15146 a_11756_50461# a_11542_50461# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15147 VSS a_5497_73719# a_5725_76207# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15148 a_50690_58500# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15149 a_22482_17890# nmat.rowon_n[6] a_22086_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1515 a_5257_62215# a_5462_62215# a_5420_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15150 a_46578_13874# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15151 a_13459_4943# ANTENNA__1187__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15152 VSS pmat.row_n[3] a_50594_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15153 a_20078_55126# pmat.en_C0_n a_20570_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15154 a_27437_28995# a_27249_28995# a_27355_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15155 a_29510_23914# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15156 a_26695_51183# a_13091_28327# pmat.col[7] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15157 vcm a_18162_8488# a_37238_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15158 VSS pmat.row_n[13] a_33526_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15159 VSS a_17927_48437# pmat.row_n[4] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X1516 a_20170_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15160 a_38150_66170# a_18162_66210# a_38242_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15161 a_24186_14512# a_18546_14510# a_24094_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15162 VDD a_9528_20407# a_9477_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15163 a_33489_43131# a_32072_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15164 VDD a_35036_32375# a_31263_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15165 a_23182_56130# a_18546_56172# a_23090_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15166 a_18546_59184# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X15167 a_31518_72234# VDD a_31122_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15168 a_19470_15882# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15169 a_47278_8488# a_18546_8486# a_47186_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1517 VDD a_22895_47893# pmat.row_n[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15170 VSS a_2389_45859# a_4927_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X15171 VSS pmat.row_n[5] a_23486_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15172 a_20474_10862# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15173 VSS pmat.row_n[7] a_48586_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15174 a_13015_62927# a_12985_62581# a_5462_62215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X15175 a_45574_60186# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15176 a_45574_19898# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15177 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot vcm.sky130_fd_sc_hd__buf_4_1.X VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X15178 a_18169_31353# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X15179 VSS a_24197_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X1518 a_29114_24958# a_18162_24552# a_29206_24552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15180 VSS pmat.row_n[10] a_35534_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15181 a_12255_34473# a_11133_34427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15182 a_9099_47753# a_8749_47381# a_9004_47741# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15183 a_28506_70226# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15184 VDD _1224_.X a_44561_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15185 a_7343_74358# a_7092_74005# a_6884_74183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15186 a_26149_27247# a_15667_27239# a_25931_27221# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15187 VSS a_26460_40517# a_26423_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15188 a_18546_71232# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X15189 VDD config_2_in[3] a_1591_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1519 VDD pmat.rowon_n[10] a_39154_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15190 a_49286_72194# a_18546_72236# a_49194_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15191 VDD pmat.rowon_n[9] a_36142_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15192 VSS _1187_.A2 a_83092_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15193 a_40250_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15194 a_46674_22512# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15195 a_8560_54281# a_7645_53909# a_8213_53877# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X15196 VDD a_29076_48695# a_30833_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X15197 a_36234_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15198 VDD pmat.rowoff_n[12] a_50198_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15199 VSS a_30523_41245# a_30463_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X152 a_37238_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1520 VSS a_4533_38279# a_5741_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X15200 a_20078_72194# a_18162_72234# a_20170_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15201 a_25494_63198# pmat.rowon_n[7] a_25098_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15202 VSS pmat.row_n[4] a_22482_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15203 VSS pmat.row_n[11] a_22482_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15204 VSS a_19083_28879# a_19541_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X15205 pmat.col_n[22] a_13091_28327# a_41418_53135# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15206 VSS a_11681_35823# a_11317_36924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X15207 a_50198_61150# a_18162_61190# a_50290_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15208 VSS ANTENNA_fanout52_A.DIODE a_31419_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15209 a_36634_14480# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1521 a_36634_63520# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15210 VDD nmat.rowon_n[6] a_39154_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15211 a_36538_20902# pmat.rowoff_n[12] a_36142_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15212 a_33130_71190# a_18162_71230# a_33222_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15213 VDD pmat.rowoff_n[4] a_40158_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15214 a_19566_24520# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15215 a_3413_6037# a_3247_6037# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15216 a_11568_40541# a_11317_40188# a_11347_40214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X15217 VDD nmat.rowon_n[1] a_23090_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15218 a_51202_24958# a_18162_24552# a_51294_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15219 vcm a_18162_58178# a_23182_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1522 vcm a_18162_18528# a_23182_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15220 a_47186_14918# a_18162_14512# a_47278_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15221 a_51294_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15222 a_51598_69222# pmat.rowon_n[13] a_51202_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15223 VSS a_1923_31743# a_2369_28157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15224 a_37146_10902# pmat.row_n[2] a_37638_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15225 VSS pmat.row_n[15] a_30514_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15226 a_2099_76725# a_1899_76001# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15227 VDD nmat.rowon_n[12] a_44174_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15228 a_29510_64202# pmat.rowon_n[8] a_29114_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15229 a_12175_27221# a_12075_24847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.35e+11p pd=2.67e+06u as=0p ps=0u w=1e+06u l=150000u
X1523 a_33222_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15230 VDD pmat.rowon_n[12] a_34134_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15231 a_14250_74941# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15232 a_27598_72556# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15233 a_15549_39867# a_15093_39638# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15234 VDD nmat.rowon_n[2] a_27106_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15235 VDD pmat.rowon_n[14] a_31122_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15236 a_24186_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15237 a_2781_23817# a_1591_23445# a_2672_23817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15238 VSS a_6619_56311# a_5730_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X15239 a_27106_62154# a_18162_62194# a_27198_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1524 a_27355_28995# a_27249_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X15240 VDD a_10147_29415# a_36278_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15241 a_19689_42405# a_18272_42693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15242 a_48586_67214# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15243 a_31214_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15244 a_3909_17209# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15245 a_19470_56170# pmat.rowon_n[0] a_19074_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15246 a_3319_76751# a_2695_76757# a_3211_77129# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15247 a_2244_20871# config_1_in[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15248 a_40567_32403# a_40903_32375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X15249 a_35230_60146# a_18546_60188# a_35138_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1525 a_46578_59182# pmat.rowon_n[3] a_46182_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15250 a_35630_64524# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15251 a_38546_59182# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15252 VSS a_30913_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X15253 a_30155_42583# a_24833_40719# a_30329_42689# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15254 vcm a_18162_19532# a_22178_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15255 a_40158_69182# a_18162_69222# a_40250_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15256 VSS pmat.row_n[1] a_42562_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15257 a_28202_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15258 a_13055_10761# a_12705_10389# a_12960_10749# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15259 a_23090_9898# pmat.row_n[1] a_23582_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1526 VDD pmat.rowon_n[5] a_40158_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15260 a_48682_63520# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15261 a_5785_60431# a_5535_57993# a_5351_60663# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15262 a_7048_23277# a_7479_22467# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15263 vcm a_18162_18528# a_35230_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15264 a_21478_18894# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15265 VSS a_8919_71615# a_8853_71689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X15266 a_19615_41959# a_12658_42895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15267 a_5939_60137# a_6175_60039# a_6133_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X15268 a_34530_17890# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15269 VDD nmat.rowon_n[4] a_43170_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1527 a_29206_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15270 a_25190_71190# a_18546_71232# a_25098_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15271 VDD a_9195_7423# a_9182_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15272 a_36142_60146# pmat.row_n[4] a_36634_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15273 a_44174_68178# a_18162_68218# a_44266_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15274 a_2672_33775# a_1757_33775# a_2325_34017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15275 VDD a_77245_39738# a_77058_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15276 VDD pmat.rowon_n[7] a_25098_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15277 VDD a_10195_30186# a_9899_30724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15278 a_47278_65166# a_18546_65208# a_47186_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15279 VDD a_2163_55233# a_2124_55107# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1528 a_31388_27247# ANTENNA__1190__A1.DIODE a_31085_27221# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X15280 VDD a_38851_28327# a_47298_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15281 a_47678_69544# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15282 a_39154_8894# pmat.row_n[0] a_39646_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15283 VSS a_25393_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X15284 a_6242_67503# a_6451_67655# a_6432_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X15285 VDD a_28116_39655# a_28020_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15286 VDD pmat.rowon_n[11] a_51202_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15287 VSS pmat.row_n[2] a_19470_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15288 a_26102_71190# pmat.row_n[15] a_26594_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15289 a_21174_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1529 a_25505_51183# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X15290 a_47186_59142# a_18162_59182# a_47278_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15291 a_6173_22895# a_5825_22901# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15292 a_51294_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15293 a_49686_8456# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15294 a_45574_8854# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15295 VSS a_23455_32447# a_23933_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X15296 VDD pmat.rowon_n[6] a_29114_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15297 a_4541_64561# a_4259_65103# a_4032_64391# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.344e+11p ps=1.48e+06u w=420000u l=150000u
X15298 a_22541_43131# a_22085_42902# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15299 a_34226_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X153 a_25802_48169# a_24602_48169# a_25466_47919# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X1530 VSS pmat.row_n[5] a_25494_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15300 a_9217_22057# a_8507_20175# a_9135_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15301 a_51598_64202# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15302 VSS a_33775_29111# a_33011_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X15303 a_1979_10927# a_1725_11254# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15304 a_51598_22910# nmat.rowon_n[1] a_51202_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15305 a_11276_55785# a_11202_55687# a_10815_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15306 a_43132_48071# a_43261_48783# a_43274_48246# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X15307 a_48190_65166# pmat.row_n[9] a_48682_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15308 a_1674_68047# a_1644_68021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X15309 VSS a_11921_37462# a_10985_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X1531 a_8268_73853# a_5403_67655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X15310 a_24186_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15311 a_5043_57399# a_4075_68583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15312 a_41558_56170# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15313 VSS VDD a_38546_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15314 a_37680_36391# a_37129_36130# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15315 a_30947_47919# a_30111_47911# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15316 a_38851_28327# a_47499_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X15317 a_24490_66210# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15318 a_38150_57134# pmat.row_n[1] a_38642_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15319 VDD a_9135_60967# a_9305_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X1532 a_7168_58799# a_7299_58951# a_6978_58799# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X15320 a_42658_55488# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15321 a_28543_27497# a_18243_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15322 a_48586_20902# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15323 a_22086_23954# pmat.row_n[15] a_22578_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15324 a_17739_50871# a_18011_50729# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15325 a_22086_19938# a_18162_19532# a_22178_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15326 vcm a_18162_23548# a_43262_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15327 a_13437_26703# a_13479_26935# a_13013_27023# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15328 VDD a_9463_50877# a_10045_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15329 a_10223_26703# a_9779_26819# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1533 a_22482_17890# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15330 VDD a_3305_27791# a_7177_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15331 a_9129_7497# a_7939_7125# a_9020_7497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15332 a_35138_22950# pmat.row_n[14] a_35630_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15333 a_28981_43493# a_28525_43655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X15334 a_28202_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15335 a_25098_55126# a_18162_55166# a_25190_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15336 a_7153_15279# a_7109_15521# a_6987_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15337 a_38546_12870# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15338 VDD a_13335_31359# a_13322_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15339 a_45574_13874# nmat.rowon_n[10] a_45178_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1534 a_20411_51157# a_19584_52423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15340 VSS pmat.row_n[2] a_42562_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15341 a_41475_31751# a_26479_32117# a_41709_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15342 a_25098_14918# pmat.row_n[6] a_25590_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15343 a_28602_17492# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15344 a_28506_23914# pmat.rowoff_n[15] a_28110_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15345 a_2012_36861# a_1895_36666# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15346 VDD a_45277_32687# a_47039_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u M=3
X15347 VSS a_39981_37462# a_40591_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15348 a_10781_42364# a_30955_42689# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X15349 a_14449_52093# a_13739_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1535 VSS a_5682_56311# a_6128_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X15350 pmat.col[26] a_17139_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15351 a_26102_18934# a_18162_18528# a_26194_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15352 VDD pmat.rowoff_n[7] a_32126_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15353 a_9317_47349# a_9099_47753# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X15354 vcm a_18162_64202# a_46274_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15355 VDD a_12197_43746# a_11261_43421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X15356 a_46182_68178# pmat.row_n[12] a_46674_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15357 VSS a_4127_37013# a_4073_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15358 a_50290_62154# a_18546_62196# a_50198_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15359 a_17503_32143# pmat.rowon_n[7] a_17285_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1536 a_20752_38341# a_20848_38341# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X15360 a_50690_66532# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15361 VSS a_4031_53034# a_3496_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X15362 VSS a_10498_19631# a_10779_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X15363 a_8456_69135# a_4991_69831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X15364 a_24501_49667# a_18823_50247# a_24405_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15365 VDD pmat.rowon_n[3] a_49194_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15366 VSS pmat.row_n[0] a_30514_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15367 a_28110_7890# VDD a_28602_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15368 VDD a_24867_53135# a_45193_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15369 VSS a_33007_37683# a_32947_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X1537 a_9528_20407# a_12875_16341# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X15370 a_11572_73309# a_11358_73309# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15371 vcm a_18162_66210# a_19166_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15372 a_29114_13914# pmat.row_n[5] a_29606_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15373 a_10703_50069# a_11138_50347# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15374 a_4253_42479# a_2419_69455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15375 a_42258_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15376 a_23182_64162# a_18546_64204# a_23090_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15377 a_33622_11468# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15378 vcm a_18162_61190# a_20170_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15379 a_23582_68540# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1538 a_26779_47197# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15380 a_1644_76181# a_1823_76181# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15381 a_3613_19061# a_3395_19465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X15382 a_18162_62194# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X15383 VSS a_2791_57703# a_3591_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X15384 a_19566_58500# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15385 a_51202_62154# pmat.row_n[6] a_51694_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15386 a_2200_12015# a_1761_11471# a_1979_12342# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X15387 a_4703_24527# a_4259_24643# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15388 a_26475_34343# a_26583_34343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15389 VDD a_2192_49159# a_2099_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1539 VDD a_2944_72104# a_2882_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X15390 VDD a_12345_39100# a_12757_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X15391 VSS pmat.row_n[3] a_19470_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15392 VDD a_12651_35823# a_12757_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15393 a_2319_67740# a_2124_67771# a_2629_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X15394 VDD a_7180_37039# a_7355_37013# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15395 a_2557_58799# a_1923_53055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15396 a_5737_76457# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15397 a_4514_34451# a_4792_34435# a_4748_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15398 VSS a_29937_31055# a_44665_45519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15399 vcm a_18162_60186# a_24186_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X154 VDD cgen.dlycontrol2_in[0] a_28431_34735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1540 a_11067_22057# a_4523_21276# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15400 VSS a_16689_43132# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X15401 a_24094_64162# pmat.row_n[8] a_24586_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15402 VDD a_3325_36495# a_4135_37815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15403 a_32126_8894# a_18162_8488# a_32218_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15404 a_19551_34191# a_19374_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15405 VSS a_39079_40947# a_39019_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15406 a_4267_35407# a_4307_35639# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15407 a_3776_77129# a_2861_76757# a_3429_76725# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15408 a_45270_13508# a_18546_13506# a_45178_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15409 vcm a_18162_10496# a_42258_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1541 a_45178_67174# a_18162_67214# a_45270_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15410 a_29051_39783# a_29159_39783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15411 a_36234_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15412 a_16163_43413# a_12237_38772# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X15413 a_21478_7850# VDD a_21082_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15414 a_4165_67753# a_1591_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15415 a_13717_21583# a_5351_19913# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15416 a_36538_70226# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15417 a_49286_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15418 a_32618_19500# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15419 a_3776_77129# a_2695_76757# a_3429_76725# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1542 VDD pmat.rowon_n[4] a_44174_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15420 a_19505_38779# a_17536_38567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X15421 a_14261_42043# a_13227_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15422 a_46804_51433# _1196_.B1 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15423 VSS a_35715_29941# a_35646_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X15424 a_11413_50095# a_10703_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15425 VDD nmat.rowon_n[13] a_36142_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15426 a_23663_38825# a_22541_38779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15427 VDD a_13091_50095# a_13278_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15428 a_50594_23914# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15429 a_2969_55535# a_2791_57703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1543 vcm a_18162_59182# a_26194_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15430 a_19488_52423# a_19584_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X15431 a_47186_22950# a_18162_22544# a_47278_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15432 a_25647_34343# a_24833_34191# a_25821_34219# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X15433 a_44266_19532# a_18546_19530# a_44174_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15434 a_51294_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15435 VDD a_11067_30287# a_15660_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X15436 a_28725_52271# ANTENNA__1197__A.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15437 a_9480_6409# a_8565_6037# a_9133_6005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15438 a_11829_55329# a_4128_64391# a_11743_55329# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X15439 a_45943_47375# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X1544 VSS VDD a_47582_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15440 a_39550_61190# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15441 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15442 VDD a_40105_47375# a_44791_43541# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15443 a_41162_71190# a_18162_71230# a_41254_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15444 a_40554_15882# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15445 VSS pmat.row_n[10] a_43566_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15446 vcm a_18162_11500# a_19166_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15447 a_29510_72234# VDD a_29114_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15448 a_9183_76359# a_6795_76989# a_9581_76207# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15449 VSS ANTENNA__1197__B.DIODE a_34030_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1545 a_17317_31849# a_10055_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X15450 VDD a_16339_43745# a_16163_43413# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15451 a_24186_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15452 VDD ANTENNA__1190__A1.DIODE a_83094_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15453 a_13985_34789# a_13529_34951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X15454 a_9305_58229# a_9577_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15455 a_36234_7484# a_18546_7482# a_36142_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15456 vcm a_18162_57174# a_44266_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15457 a_13269_31433# a_12079_31061# a_13160_31433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15458 VDD a_6639_23413# nmat.sw VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15459 VDD a_11927_27399# a_22138_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1546 VDD a_14589_40726# a_13653_40956# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X15460 a_35715_43447# a_34593_43493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X15461 a_9135_26409# a_4516_21531# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15462 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top vcm.sky130_fd_sc_hd__buf_4_2.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X15463 VDD a_11067_64015# a_17317_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15464 a_20474_18894# nmat.rowon_n[5] a_20078_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15465 a_44570_14878# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15466 a_36459_29673# a_36453_29199# a_36723_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15467 a_28591_36519# a_23821_35279# a_28765_36395# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X15468 VDD a_24895_35253# a_24719_35253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X15469 a_20848_39429# a_19689_39141# a_20811_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1547 a_9664_47753# a_8749_47381# a_9317_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X15470 a_27502_24918# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15471 a_11233_76207# a_10239_77295# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15472 a_35630_72556# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15473 VSS a_26891_28327# a_35224_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15474 nmat.rowon_n[6] a_14460_12265# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X15475 a_33526_17890# nmat.rowon_n[6] a_33130_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15476 VDD a_1643_61493# a_1591_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15477 vcm a_18162_69222# a_21174_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15478 a_31122_16926# pmat.row_n[8] a_31614_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15479 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1548 VDD a_10383_75637# a_6795_76989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15480 a_25575_31055# a_25042_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15481 a_8749_47381# a_8583_47381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15482 VDD pmat.rowon_n[4] a_35138_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15483 a_48682_71552# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15484 a_5779_13255# a_4895_12559# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15485 vcm a_18162_7484# a_34226_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15486 a_21174_57134# a_18546_57176# a_21082_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15487 a_5603_32687# a_5253_32687# a_5508_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15488 a_10041_74281# a_9581_73487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15489 a_44382_41167# a_35312_31599# a_44382_40847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X1549 a_30210_57134# a_18546_57176# a_30118_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15490 a_27198_9492# a_18546_9490# a_27106_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15491 a_34948_50069# a_26891_28327# a_35077_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X15492 VSS pmat.row_n[6] a_21478_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15493 a_34226_56130# a_18546_56172# a_34134_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15494 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15495 a_12925_60431# a_11007_58229# a_11797_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X15496 VSS a_4508_65845# a_4446_65871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15497 VSS pmat.row_n[5] a_34530_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15498 a_1907_11254# a_1725_11254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15499 a_6832_66191# a_5687_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X155 VSS ANTENNA__1184__B1.DIODE nmat.col[19] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X1550 VSS a_25695_28111# a_35161_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X15500 VDD pmat.rowon_n[15] a_25098_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15501 a_15839_49525# a_13091_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15502 VDD nmat.rowon_n[14] a_43170_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15503 a_13073_54997# a_12907_54997# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15504 a_10117_54697# a_9581_56079# a_9963_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15505 VDD a_3583_11775# a_3570_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15506 VSS a_27763_27221# nmat.col[8] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15507 a_19717_49257# a_16083_50069# a_19622_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X15508 a_11057_67503# a_10499_67503# a_10975_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15509 a_25190_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1551 VSS a_47591_35407# _1192_.A2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X15510 a_49590_69222# pmat.rowon_n[13] a_49194_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15511 VSS pmat.row_n[10] a_46578_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15512 a_50594_64202# pmat.rowon_n[8] a_50198_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15513 VDD nmat.rowon_n[14] a_19074_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15514 a_44666_23516# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15515 a_31122_9898# pmat.row_n[1] a_31614_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15516 a_44266_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15517 a_26983_31849# a_23933_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15518 VSS a_22059_37683# a_21999_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15519 a_51294_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1552 VDD a_77882_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_2.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15520 VSS a_11979_47068# a_11910_47197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15521 VDD a_10391_62911# a_10378_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15522 VDD pmat.rowon_n[14] a_29114_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15523 a_47278_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15524 a_19074_11906# a_18162_11500# a_19166_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15525 a_20170_18528# a_18546_18526# a_20078_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15526 a_40554_56170# pmat.rowon_n[0] a_40158_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15527 VDD nmat.rowon_n[5] a_37146_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15528 VDD a_10287_61127# a_10195_59861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15529 a_23486_66210# pmat.rowon_n[10] a_23090_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1553 a_26498_16886# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15530 a_10765_24233# a_9075_28023# a_10693_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15531 a_33222_17524# a_18546_17522# a_33130_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15532 VSS a_17927_47349# pmat.row_n[0] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X15533 a_47678_14480# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15534 VDD pmat.rowoff_n[15] a_21082_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15535 a_45178_15922# a_18162_15516# a_45270_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15536 a_48282_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15537 a_33489_42043# a_30523_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15538 a_9415_51433# a_9319_50639# a_9319_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15539 VDD pmat.rowoff_n[4] a_51202_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1554 a_21147_49525# a_20619_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15540 a_2847_41151# a_2672_41225# a_3026_41213# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15541 VSS a_20776_51959# a_19579_52789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X15542 a_2672_50095# a_1757_50095# a_2325_50337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15543 VDD a_5363_33551# a_12079_31061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15544 VDD a_6904_40303# a_7079_40277# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15545 a_78448_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_1.X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15546 vcm a_18162_14512# a_21174_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15547 a_44570_55166# VSS a_44174_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15548 a_27502_65206# pmat.rowon_n[9] a_27106_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15549 VDD a_9195_60039# a_7457_62037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X1555 VSS a_9460_10615# a_8111_11209# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15550 vcm a_18162_13508# a_34226_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15551 VDD nmat.rowon_n[7] a_14460_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15552 a_48190_10902# pmat.row_n[2] a_48682_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15553 a_22178_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15554 a_42258_61150# a_18546_61192# a_42166_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15555 VDD pmat.rowon_n[12] a_45178_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15556 a_25098_63158# a_18162_63198# a_25190_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15557 a_39634_48463# a_38557_48469# a_39472_48841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15558 a_10339_21263# a_8197_20871# a_10441_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15559 VSS a_10049_60663# a_10423_64786# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1556 a_1925_20871# cgen.dlycontrol4_in[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15560 a_27198_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15561 a_8263_20969# a_8197_20871# a_8155_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15562 a_4791_30877# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15563 a_2107_39049# a_1757_38677# a_2012_39037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15564 a_14372_4399# ANTENNA__1190__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15565 a_6917_27907# a_4516_21531# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15566 a_6251_49007# a_5805_49007# a_6155_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15567 vcm a_18162_72234# a_46274_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15568 a_6524_69679# a_5497_62839# a_6334_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15569 VDD nmat.rowon_n[10] a_28110_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1557 VSS pmat.row_n[6] a_30514_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15570 a_24847_35279# a_11041_36596# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15571 a_50290_70186# a_18546_70228# a_50198_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15572 a_8363_73865# a_8013_73493# a_8268_73853# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15573 VDD a_32687_46607# a_33986_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X15574 a_46274_60146# a_18546_60188# a_46182_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15575 nmat.rowoff_n[1] a_14839_7119# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X15576 VSS a_3325_20175# a_8859_22467# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15577 VDD pmat.rowon_n[11] a_49194_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15578 a_46674_64524# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15579 a_43170_61150# pmat.row_n[5] a_43662_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1558 a_24197_42405# a_23741_42567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X15580 vcm a_18162_19532# a_33222_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15581 a_40837_46261# a_46897_40303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X15582 VDD pmat.rowon_n[6] a_50198_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15583 a_22537_36911# a_22111_36950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15584 a_32522_18894# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15585 a_23182_72194# a_18546_72236# a_23090_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15586 a_36634_56492# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15587 a_38642_7452# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15588 a_2195_51701# a_2398_51859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15589 a_19166_62154# a_18546_62196# a_19074_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1559 a_17336_43439# a_17159_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15590 a_8831_24501# a_8399_18115# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15591 a_49590_22910# nmat.rowon_n[1] a_49194_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15592 a_20570_22512# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15593 a_19566_66532# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15594 a_41254_22544# a_18546_22542# a_41162_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15595 a_51202_70186# pmat.row_n[14] a_51694_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15596 VDD pmat.rowon_n[8] a_23090_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15597 a_37238_12504# a_18546_12502# a_37146_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15598 a_47186_60146# pmat.row_n[4] a_47678_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15599 VDD VDD a_48190_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X156 VSS a_1586_8439# a_3247_6037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1560 a_24094_10902# a_18162_10496# a_24186_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15600 VSS VDD a_44570_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15601 a_19074_56130# a_18162_56170# a_19166_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15602 VSS a_1957_43567# a_11173_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15603 a_3227_22351# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15604 cgen.dlycontrol1_in[4] a_1591_35951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15605 VDD a_12792_12937# a_12967_12863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15606 a_24094_72194# VDD a_24586_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15607 a_8861_24527# a_7415_29397# a_8333_24847# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X15608 VDD a_13091_28327# a_26437_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X15609 a_35534_70226# pmat.rowon_n[14] a_35138_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1561 a_19409_40719# a_19143_41085# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15610 a_2099_25236# a_2191_25045# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15611 a_21082_14918# a_18162_14512# a_21174_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15612 a_45270_21540# a_18546_21538# a_45178_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15613 a_25494_9858# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15614 a_10562_15645# a_9485_15279# a_10400_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15615 a_24586_60508# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15616 a_32218_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15617 VSS a_1781_9308# a_2200_9661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15618 VDD a_2375_63316# a_1895_63866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15619 a_22097_28995# a_10441_21263# a_22015_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1562 VSS a_7111_74575# a_2149_45717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X15620 cgen.dlycontrol3_in[4] a_1591_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X15621 a_12461_19881# a_9441_20189# a_11892_21959# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15622 a_17459_37143# a_17675_37001# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15623 a_11542_50461# a_11455_50237# a_11138_50347# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X15624 VDD a_3305_17999# a_5979_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15625 a_5415_71543# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15626 VDD a_34949_52245# pmat.col_n[14] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15627 a_18777_51183# a_18429_51189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X15628 a_1757_43029# a_1591_43029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X15629 a_38546_61190# pmat.rowon_n[5] a_38150_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1563 a_49194_7890# VDD a_49686_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15630 a_29735_40183# a_28613_40229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X15631 a_77245_40202# a_77341_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15632 a_32072_38567# a_30913_38779# a_32035_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X15633 a_4719_30287# a_5423_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X15634 a_9466_77117# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15635 a_22482_67214# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15636 a_11961_27907# a_5991_23983# a_11889_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15637 a_18546_13506# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X15638 VDD a_5579_12394# a_5411_12167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15639 a_49194_18934# pmat.row_n[10] a_49686_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1564 a_35230_20536# a_18546_20534# a_35138_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15640 VSS VDD a_49590_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15641 a_43262_69182# a_18546_69224# a_43170_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15642 vcm a_18162_66210# a_40250_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15643 a_8305_20871# a_12047_14165# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X15644 a_50198_13914# pmat.row_n[5] a_50690_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15645 a_35534_66210# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15646 a_12985_62581# a_13432_62581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15647 a_39246_59142# a_18546_59184# a_39154_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15648 a_40650_19500# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15649 VDD a_4492_32375# a_4123_32661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1565 VDD nmat.sample a_18546_8486# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X15650 a_33130_23954# pmat.row_n[15] a_33622_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15651 a_13699_72777# a_13349_72405# a_13604_72765# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15652 VSS a_7436_58487# a_7299_58951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15653 a_33130_19938# a_18162_19532# a_33222_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15654 a_11212_14191# a_10593_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15655 VSS pmat.row_n[8] a_39550_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15656 VDD a_34724_44527# a_34830_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15657 VSS a_12228_40693# a_27566_43805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15658 a_6891_15279# a_6375_15279# a_6796_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X15659 a_43566_14878# nmat.rowon_n[9] a_43170_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1566 VDD pmat.sample_n a_18162_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X15660 a_37238_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15661 VDD a_8583_29199# a_25327_28992# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15662 VDD a_18241_31698# a_32319_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X15663 a_32522_59182# pmat.rowon_n[3] a_32126_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15664 a_10159_52047# a_9463_50877# a_10052_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X15665 a_23090_15922# pmat.row_n[7] a_23582_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15666 a_26594_18496# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15667 a_26498_24918# VSS a_26102_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15668 VDD a_37612_30663# a_37143_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15669 VDD nmat.rowon_n[7] a_30118_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1567 a_12461_29673# a_8583_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15670 VSS a_4429_76751# a_4993_77071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X15671 vcm a_18162_65206# a_44266_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15672 VDD a_7373_49007# a_8121_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X15673 a_8853_71689# a_7663_71317# a_8744_71689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15674 a_44174_69182# pmat.row_n[13] a_44666_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15675 VDD a_2021_26677# a_2879_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X15676 a_29404_36165# a_28245_35877# a_29308_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X15677 VSS a_14011_19087# a_10515_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X15678 a_11693_70767# a_11345_70773# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15679 VDD a_3305_15823# a_6623_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1568 a_38546_9858# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15680 a_45251_53047# _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X15681 a_14917_23983# a_14475_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15682 a_28774_30287# a_18563_27791# a_28336_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X15683 a_29510_57174# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15684 VDD a_26041_36374# a_26272_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15685 VDD a_39079_40947# a_39321_42333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X15686 a_4700_44655# a_4257_34319# a_4525_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15687 a_31122_67174# a_18162_67214# a_31214_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15688 VSS VDD a_33526_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15689 a_19083_28879# a_18973_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.225e+11p pd=3.9e+06u as=0p ps=0u w=650000u l=150000u
X1569 a_22178_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15690 a_21082_7890# a_18162_7484# a_21174_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15691 a_21174_65166# a_18546_65208# a_21082_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15692 a_45270_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15693 VSS a_22493_31353# a_22427_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15694 a_21574_69544# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15695 a_34226_64162# a_18546_64204# a_34134_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15696 a_7845_67503# a_7803_67655# a_7435_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X15697 a_21082_59142# a_18162_59182# a_21174_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15698 a_31214_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15699 a_34626_68540# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X157 pmat.row_n[5] a_21883_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1570 VDD a_36561_38780# a_36167_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X15700 VSS a_3305_17999# a_6661_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15701 a_4791_30877# a_4167_30511# a_4683_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15702 a_30913_43131# a_30140_43781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15703 a_41703_29423# a_38905_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15704 a_45884_38377# a_45866_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15705 VSS vcm.sky130_fd_sc_hd__nand2_1_1.A a_77980_40594# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15706 a_22086_65166# pmat.row_n[9] a_22578_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15707 vcm a_18162_16520# a_39246_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15708 a_8268_73853# a_5403_67655# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15709 a_43262_14512# a_18546_14510# a_43170_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1571 pmat.row_n[12] a_19491_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15710 a_43566_71230# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15711 vcm a_18162_11500# a_40250_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15712 a_15667_28111# a_13479_26935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X15713 a_2099_24746# a_2191_24501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15714 VSS a_2046_30184# a_2051_29973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15715 VSS a_24374_29941# a_27976_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X15716 a_50594_72234# VDD a_50198_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15717 vcm a_18162_60186# a_35230_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15718 a_26671_46831# a_26155_46831# a_26576_46831# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X15719 a_35138_64162# pmat.row_n[8] a_35630_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1572 VDD _1154_.X a_83196_3561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.955e+12p ps=1.791e+07u w=1e+06u l=150000u M=4
X15720 a_5043_37191# a_4257_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15721 a_22482_20902# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15722 VSS pmat.row_n[15] a_25494_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15723 a_47278_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15724 a_25098_56130# pmat.row_n[0] a_25590_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15725 VDD pmat.rowon_n[1] a_32126_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15726 a_16607_36911# a_16430_36911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15727 a_47582_70226# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15728 vcm a_18162_22544# a_30210_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15729 a_7067_53511# a_7163_53333# a_7465_53359# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1573 VDD a_1591_58799# a_2603_58368# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X15730 a_29206_15516# a_18546_15514# a_29114_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15731 VSS a_8443_20719# a_18795_28882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15732 a_45178_23954# a_18162_23548# a_45270_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15733 a_45196_47695# a_45112_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15734 a_17874_50755# a_16083_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15735 a_5417_11445# a_5768_9527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15736 a_37542_62194# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15737 VDD a_23823_47679# a_23810_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15738 a_2107_20553# a_1757_20181# a_2012_20541# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15739 VDD a_6608_70455# a_6559_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1574 a_9217_23983# a_8291_23983# a_9217_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.65e+11p pd=2.93e+06u as=2.25e+11p ps=2.45e+06u w=1e+06u l=150000u
X15740 a_32522_12870# pmat.rowoff_n[4] a_32126_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15741 a_44570_63198# pmat.rowon_n[7] a_44174_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15742 VSS pmat.row_n[4] a_41558_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15743 a_23815_48981# a_23971_49140# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X15744 a_29114_55126# VDD a_29606_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15745 VDD a_9827_53379# a_10363_53153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15746 VSS pmat.row_n[11] a_41558_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15747 VSS pmat.row_n[14] a_24490_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15748 VSS a_13327_70741# a_13285_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15749 a_7865_58553# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1575 a_25280_46831# a_25189_46287# a_25180_46831# VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X15750 vcm a_18162_21540# a_34226_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15751 VDD a_12967_58559# a_11007_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15752 vcm a_18162_71230# a_38242_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15753 VDD a_11067_27239# a_28267_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15754 a_22178_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15755 a_13728_59663# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15756 a_38642_24520# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15757 VSS a_2199_13887# a_2369_8573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15758 a_3609_9615# a_3415_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15759 VDD nmat.rowon_n[1] a_42166_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1576 a_13439_8207# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15760 vcm a_18162_58178# a_42258_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15761 a_29510_10862# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15762 VDD a_4535_38377# a_4979_38127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15763 VSS pmat.row_n[5] a_27502_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15764 a_12397_16367# a_12353_16609# a_12231_16367# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15765 a_17113_42405# a_16657_42567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15766 a_35312_31599# a_35084_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15767 VSS _1183_.A2 a_39949_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15768 a_31518_18894# nmat.rowon_n[5] a_31122_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15769 a_20267_27497# a_8568_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X1577 a_1757_26159# a_1591_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15770 VSS config_2_in[3] a_1591_33231# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X15771 a_8551_7497# a_8105_7125# a_8455_7497# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X15772 VDD a_10975_18231# a_10975_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15773 a_1644_68021# a_1674_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X15774 a_43261_51727# a_23395_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15775 a_39154_20942# pmat.row_n[12] a_39646_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15776 VSS a_6975_76823# a_9225_76207# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X15777 a_46674_72556# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15778 a_39154_16926# a_18162_16520# a_39246_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15779 VDD pmat.rowon_n[14] a_50198_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1578 VDD a_13503_36893# a_13529_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X15780 vcm a_18162_69222# a_32218_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15781 a_43262_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15782 a_40158_11906# a_18162_11500# a_40250_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15783 VDD a_10329_30753# a_10219_30877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15784 VSS a_25061_43132# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X15785 a_32771_31599# a_9963_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X15786 VDD pmat.rowon_n[4] a_46182_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15787 vcm a_18162_59182# a_28202_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15788 VSS a_3339_70759# a_6829_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15789 a_46182_62154# a_18162_62194# a_46274_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1579 VSS a_2163_71997# a_2124_72123# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15790 a_32218_57134# a_18546_57176# a_32126_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15791 a_50290_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15792 a_29114_72194# a_18162_72234# a_29206_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15793 a_28506_16886# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15794 a_33222_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15795 a_19166_70186# a_18546_70228# a_19074_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15796 VSS pmat.row_n[6] a_32522_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15797 VDD a_6975_76823# a_7631_75895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15798 VDD pmat.rowoff_n[15] a_19074_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15799 a_5979_23145# nmat.sw a_5907_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 VSS a_29076_48695# a_28629_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X1580 a_39154_58138# a_18162_58178# a_39246_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15800 VDD VDD a_23090_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15801 a_37238_20536# a_18546_20534# a_37146_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15802 VDD pmat.rowoff_n[4] a_49194_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15803 vcm a_18162_19532# a_41254_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15804 a_11077_76207# a_11023_76359# a_10995_76207# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15805 a_19074_64162# a_18162_64202# a_19166_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15806 VSS a_2319_61493# a_2250_61519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X15807 VSS a_16800_47213# a_16911_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15808 VDD a_10239_14183# a_13277_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15809 a_23182_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1581 a_50198_20942# pmat.row_n[12] a_50690_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15810 pmat.col_n[9] a_18243_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X15811 VSS pmat.row_n[11] a_44570_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15812 vcm.sky130_fd_sc_hd__nand2_1_1.Y vcm.sky130_fd_sc_hd__nand2_1_1.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15813 a_21082_22950# a_18162_22544# a_21174_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15814 comp.adc_inverter_1.out comp.adc_inverter_1.in VDD VDD sky130_fd_pr__pfet_01v8 ad=2.394e+11p pd=2.82e+06u as=0p ps=0u w=420000u l=150000u M=2
X15815 vcm.sky130_fd_sc_hd__buf_4_1.X a_77980_40594# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X15816 a_34134_21946# a_18162_21540# a_34226_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15817 a_21478_67214# pmat.rowon_n[11] a_21082_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15818 VDD pmat.rowon_n[7] a_44174_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15819 a_31214_18528# a_18546_18526# a_31122_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1582 VDD a_38905_28853# a_37827_30793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15820 VDD a_19268_34191# a_19374_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15821 a_51598_56170# pmat.rowon_n[0] a_51202_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15822 VDD nmat.rowon_n[5] a_48190_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15823 VDD ANTENNA__1196__A2.DIODE pmat.col_n[29] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X15824 VSS pmat.row_n[1] a_35534_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15825 a_12813_31029# a_12595_31433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15826 VSS pmat.row_n[9] a_30514_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15827 VDD a_22493_31353# a_22523_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15828 VDD a_2199_13887# a_5967_5461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15829 VSS pmat.row_n[2] a_38546_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1583 a_50198_16926# a_18162_16520# a_50290_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15830 a_45574_9858# nmat.rowon_n[14] a_45178_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15831 a_31767_47919# a_30999_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X15832 a_40250_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15833 a_18546_21538# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X15834 a_13555_37782# a_11497_38543# a_13483_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X15835 VSS a_23707_40693# a_12197_41570# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15836 a_49194_69182# a_18162_69222# a_49286_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15837 a_10867_41271# a_10927_41245# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15838 vcm a_18162_14512# a_32218_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15839 a_3325_23439# a_2847_23743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1584 VSS a_2411_16101# a_5865_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15840 a_6829_57487# a_4025_54965# a_6611_57399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15841 vcm a_18162_56170# a_31214_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15842 a_45432_46983# a_33423_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15843 a_39246_67174# a_18546_67216# a_39154_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15844 a_23757_47753# a_22567_47381# a_23648_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15845 VSS a_3571_13627# a_10791_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15846 VDD pmat.rowon_n[13] a_43170_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15847 a_31518_13874# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15848 VDD a_5363_70543# a_11165_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15849 a_43262_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1585 a_25494_63198# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15850 a_40158_56130# a_18162_56170# a_40250_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15851 a_2215_40847# a_1591_40853# a_2107_41225# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15852 a_6795_18319# a_3305_17999# a_6467_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X15853 a_26194_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15854 a_28506_57174# pmat.rowon_n[1] a_28110_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15855 a_23090_66170# a_18162_66210# a_23182_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15856 VDD a_13620_10761# a_13795_10687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15857 a_15477_31599# a_14287_31599# a_15368_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15858 a_41162_23954# pmat.row_n[15] a_41654_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15859 a_3977_33609# a_2787_33237# a_3868_33609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1586 a_6909_28879# a_4516_21531# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15860 a_20848_36165# a_19689_35877# a_20752_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X15861 a_41162_19938# a_18162_19532# a_41254_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15862 VDD a_3175_59585# a_3136_59459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15863 VSS a_12449_39605# a_12383_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15864 a_44666_65528# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15865 a_2464_54991# a_2250_54991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15866 VSS a_3111_53333# a_2944_52789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15867 a_7250_42845# a_6173_42479# a_7088_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15868 a_42658_8456# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15869 VSS a_15101_29423# a_28803_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X1587 a_2203_23817# a_1757_23445# a_2107_23817# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X15870 a_23700_42919# a_22541_43131# a_23663_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X15871 a_30863_46831# a_29076_48695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X15872 a_44174_55126# a_18162_55166# a_44266_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15873 VDD a_29036_41831# a_28940_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15874 VSS pmat.row_n[7] a_33526_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15875 a_34530_24918# nmat.en_bit_n[1] a_34134_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15876 a_30514_60186# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15877 a_30514_19898# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15878 VSS pmat.row_n[10] a_20474_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15879 a_14933_37429# a_14600_37607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1588 VSS a_33467_46261# a_45450_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X15880 a_11391_69831# a_10864_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15881 a_47582_23914# pmat.rowoff_n[15] a_47186_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15882 a_44174_14918# pmat.row_n[6] a_44666_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15883 VSS pmat.row_n[12] a_44570_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15884 a_34226_72194# a_18546_72236# a_34134_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15885 VDD pmat.rowon_n[9] a_21082_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15886 a_47678_56492# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15887 a_27106_24958# VDD a_27598_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15888 VSS pmat.row_n[0] a_24490_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15889 VDD nmat.rowon_n[15] a_28110_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1589 VSS a_10058_60431# a_10045_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X15890 a_44741_36201# a_43533_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15891 a_31614_22512# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15892 a_13985_41317# a_10651_42035# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15893 VSS a_1586_33927# a_6099_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15894 VSS a_7779_22583# a_7479_22467# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15895 a_21174_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15896 a_9367_53511# a_9639_53339# a_9597_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15897 VDD a_7415_29397# a_9415_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15898 a_20184_46983# a_20267_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15899 a_37542_15882# pmat.rowoff_n[7] a_37146_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X159 a_23486_58178# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1590 a_39154_17930# pmat.row_n[9] a_39646_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15900 VDD a_9133_6005# a_9023_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15901 a_6639_63927# a_6451_67655# a_6806_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X15902 pmat.en_bit_n[2] a_15753_28879# a_22576_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X15903 VDD nmat.rowon_n[6] a_24094_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15904 vcm a_18162_24552# a_39246_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15905 a_21574_14480# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15906 a_21478_20902# pmat.rowoff_n[12] a_21082_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15907 VDD a_17536_38567# a_17440_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15908 a_35138_72194# VDD a_35630_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15909 a_38907_47753# a_38557_47381# a_38812_47741# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X1591 VSS pmat.row_n[15] a_39550_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15910 a_46578_70226# pmat.rowon_n[14] a_46182_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15911 a_38642_58500# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15912 a_32126_14918# a_18162_14512# a_32218_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15913 VSS pmat.row_n[3] a_38546_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15914 a_13555_37455# a_13301_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15915 a_36538_62194# pmat.rowon_n[6] a_36142_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15916 a_25590_13476# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15917 a_4496_14013# a_4379_13818# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X15918 a_22086_10902# pmat.row_n[2] a_22578_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15919 VSS _1184_.A2 a_38379_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1592 VDD a_7085_15055# a_7717_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15920 VDD VSS a_28110_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15921 VSS a_4036_67477# a_3983_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X15922 a_4399_48169# a_4128_46983# a_4291_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15923 a_20474_68218# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15924 a_29206_23548# a_18546_23546# a_29114_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15925 vcm a_18162_8488# a_39246_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15926 a_50594_57174# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15927 a_11867_26819# a_5991_23983# a_11795_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15928 VDD a_26659_34967# a_12069_36341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X15929 a_33765_35877# a_33309_36039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X1593 VDD a_16381_35286# a_17808_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X15930 a_16848_47081# a_16800_47213# a_16764_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15931 a_33526_67214# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15932 a_14553_27247# a_5351_19913# a_14471_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15933 VDD a_2046_30184# a_5087_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15934 a_49286_8488# a_18546_8486# a_49194_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15935 a_13798_22351# a_14005_22589# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15936 a_13801_34427# a_12568_35077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15937 a_28506_10862# nmat.rowon_n[13] a_28110_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15938 a_10676_30511# a_9761_30511# a_10329_30753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15939 a_51694_19500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1594 a_43662_15484# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15940 a_20170_60146# a_18546_60188# a_20078_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15941 a_20570_64524# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15942 a_23486_59182# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15943 a_2012_8573# a_1895_8378# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15944 a_7796_62723# a_7212_62607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15945 vcm a_18162_61190# a_29206_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15946 VDD a_19582_46983# a_19531_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15947 a_24638_49159# a_22499_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15948 a_20659_49140# a_20267_50345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15949 a_33622_63520# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1595 a_43566_21906# nmat.rowon_n[2] a_43170_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15950 a_9957_26819# a_9485_27247# a_9861_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15951 a_9953_53903# a_6559_33767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15952 VDD pmat.rowoff_n[12] a_38150_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15953 VSS a_9485_27247# a_9779_26819# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15954 VDD a_2659_35015# a_6651_44661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15955 VSS a_1781_9308# a_2200_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15956 a_38150_61150# a_18162_61190# a_38242_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15957 VSS _1194_.B1 a_23844_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15958 a_27887_41271# a_28281_41245# a_27947_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X15959 a_19689_44581# a_17996_44007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X1596 a_40158_12910# pmat.row_n[4] a_40650_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15960 a_14933_37429# a_14600_37607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15961 a_12237_38772# a_12543_39126# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15962 a_12174_50461# a_11416_50363# a_11611_50332# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15963 a_22725_40229# a_22269_40391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X15964 a_27502_58178# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15965 a_21082_60146# pmat.row_n[4] a_21574_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15966 a_4801_58255# a_2419_69455# a_4885_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15967 VSS a_35039_29941# a_31263_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15968 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15969 VDD a_10699_72943# a_11499_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1597 VSS a_22787_34165# a_11921_37462# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15970 a_2012_64061# a_1895_63866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15971 a_29797_51701# a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15972 VSS a_9797_9813# a_9731_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15973 a_39154_24958# a_18162_24552# a_39246_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15974 VDD a_16607_36911# a_16713_36911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15975 a_43262_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15976 vcm a_18162_67214# a_28202_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15977 a_39246_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15978 a_32218_65166# a_18546_65208# a_32126_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15979 VSS a_10239_14183# a_14287_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1598 a_32522_66210# pmat.rowon_n[10] a_32126_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15980 VSS a_36617_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X15981 VSS pmat.row_n[5] a_35534_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15982 a_32618_69544# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15983 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15984 VDD a_3305_27791# a_4627_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.05e+11p ps=7.61e+06u w=1e+06u l=150000u M=2
X15985 VSS a_43720_32143# a_46522_34293# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X15986 a_2561_46070# a_2389_45859# a_2347_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X15987 a_32126_59142# a_18162_59182# a_32218_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15988 VDD a_5245_56053# a_3967_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X15989 a_4154_47695# a_2315_44124# a_3987_47375# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X1599 VDD pmat.rowon_n[1] a_46182_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15990 a_46578_24918# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15991 a_28202_10496# a_18546_10494# a_28110_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15992 vcm a_18162_7484# a_28202_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15993 a_46934_53135# ANTENNA__1197__A.DIODE a_46848_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15994 vcm a_18162_59182# a_36234_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15995 VDD a_7658_71543# a_7663_71317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15996 a_19166_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15997 a_40250_57134# a_18546_57176# a_40158_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15998 a_5331_53511# a_2419_53351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15999 a_33130_65166# pmat.row_n[9] a_33622_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u M=887
X160 a_37542_71230# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1600 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16000 a_36538_16886# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16001 VSS a_11892_21959# a_11987_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16002 VSS a_13718_68591# a_14289_66421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16003 a_4135_61225# a_4081_61127# a_4041_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X16004 VSS a_11883_62063# a_11883_66191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16005 VSS pmat.row_n[6] a_40554_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16006 a_12368_35823# a_12191_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16007 a_31847_52271# _1154_.X pmat.col[1] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16008 a_18162_65206# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X16009 a_10991_68591# a_10740_68841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X1601 a_23090_22950# pmat.row_n[14] a_23582_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16010 a_49590_15882# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16011 a_1757_20181# a_1591_20181# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16012 a_20474_21906# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16013 VSS VDD a_23486_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16014 a_50594_10862# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16015 a_13915_47375# a_13830_47607# a_13697_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16016 a_23090_57134# pmat.row_n[1] a_23582_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16017 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16018 VDD pmat.rowon_n[15] a_44174_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16019 a_33526_20902# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1602 VDD pmat.rowoff_n[15] a_30118_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16020 a_2369_64061# a_2325_63669# a_2203_64073# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16021 a_27198_16520# a_18546_16518# a_27106_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16022 a_1644_68565# a_1823_68565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16023 VDD a_6651_33239# a_2046_30184# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16024 a_38793_49007# a_38515_49035# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X16025 a_18169_31353# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16026 a_25098_9898# pmat.row_n[1] a_25590_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16027 VSS pmat.row_n[7] a_26498_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16028 a_29510_18894# nmat.rowon_n[5] a_29114_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16029 a_23486_12870# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1603 a_9589_6409# a_8399_6037# a_9480_6409# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X16030 a_45295_44905# a_43720_32143# a_45199_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16031 a_30514_13874# nmat.rowon_n[10] a_30118_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16032 VDD a_8443_20719# a_18795_28882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16033 a_30913_42043# a_29036_41831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16034 a_5070_27023# a_2952_25045# a_5320_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16035 pmat.rowoff_n[6] a_14458_58799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16036 a_48586_62194# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16037 a_23541_52245# _1192_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16038 a_4865_12533# a_5331_13951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16039 a_9393_17455# a_8305_20871# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X1604 cgen.dlycontrol3_in[0] a_1591_44655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16040 VSS a_2122_17455# a_2228_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16041 a_50198_72194# a_18162_72234# a_50290_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16042 vcm a_18162_64202# a_31214_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16043 a_31122_68178# pmat.row_n[12] a_31614_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16044 VDD ANTENNA__1395__A2.DIODE a_46765_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16045 VDD ANTENNA__1195__A1.DIODE a_40041_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16046 a_42562_66210# pmat.rowon_n[10] a_42166_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16047 a_82735_2223# _1183_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16048 a_27106_58138# pmat.row_n[2] a_27598_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16049 VDD pmat.rowoff_n[15] a_40158_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1605 a_9227_20291# a_9441_20189# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16050 VDD a_2847_16127# a_2834_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16051 a_13559_23439# a_7026_24527# a_13641_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X16052 a_27502_11866# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16053 a_49686_24520# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16054 VSS a_11910_43047# a_11915_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16055 a_40158_64162# a_18162_64202# a_40250_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16056 a_83741_26409# ANTENNA__1395__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16057 a_39246_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16058 VSS a_29937_31055# a_46994_34639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16059 VDD a_3305_15823# a_7407_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1606 a_30118_64162# a_18162_64202# a_30210_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16060 a_18703_51843# a_16083_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16061 a_39550_64202# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16062 VDD a_6168_32687# a_6343_32661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16063 VSS a_2021_11043# a_3142_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16064 a_47582_8854# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16065 a_6975_34538# a_7067_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16066 a_37146_21946# pmat.row_n[13] a_37638_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16067 a_37146_17930# a_18162_17524# a_37238_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16068 VDD nmat.rowon_n[9] a_43170_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16069 a_41254_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1607 a_29206_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16070 VDD VSS a_26102_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16071 a_10781_42869# a_31783_42689# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X16072 a_44174_63158# a_18162_63198# a_44266_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16073 a_17996_40743# a_16837_40955# a_17959_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16074 a_6205_5487# a_6170_5739# a_5967_5461# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16075 VDD a_9337_15033# a_9367_14774# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16076 VDD a_10379_8439# a_9731_8439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16077 a_19470_67214# pmat.rowon_n[11] a_19074_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16078 vcm a_18162_15516# a_26194_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16079 a_49590_56170# pmat.rowon_n[0] a_49194_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1608 a_42562_7850# VDD a_42166_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16080 a_23880_41605# a_22817_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X16081 a_11803_20535# a_8305_20871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16082 a_30210_13508# a_18546_13506# a_30118_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16083 VDD nmat.rowon_n[10] a_47186_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16084 a_44666_10464# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16085 a_21174_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16086 a_27598_20504# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16087 VSS pmat.row_n[12] a_42562_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16088 a_27198_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16089 a_2107_8585# a_1591_8213# a_2012_8573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1609 a_31535_49525# a_25879_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16090 a_21478_70226# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16091 a_34226_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16092 a_5621_48783# a_5411_48695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16093 a_9481_49007# a_8907_48437# a_9135_49257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X16094 a_2007_76970# a_2099_76725# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16095 a_14553_62313# a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16096 a_34530_8854# nmat.rowon_n[15] a_34134_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16097 a_51598_18894# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16098 a_50690_8456# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16099 a_10932_21959# a_4523_21276# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X161 vcm a_18162_60186# a_29206_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1610 a_13604_72765# a_6451_67655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X16100 a_25688_32117# a_26479_32117# a_26425_32463# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16101 VDD a_12328_48168# a_12266_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16102 VDD a_4659_53738# a_4491_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16103 a_2672_23817# a_1757_23445# a_2325_23413# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16104 VDD nmat.rowon_n[13] a_21082_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16105 VDD a_11711_50959# a_38515_49035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16106 a_38242_62154# a_18546_62196# a_38150_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16107 a_12107_62037# a_11842_59887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16108 a_38642_66532# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16109 a_32126_22950# a_18162_22544# a_32218_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1611 a_12353_16609# a_12135_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X16110 VDD pmat.rowon_n[8] a_42166_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16111 a_28110_12910# a_18162_12504# a_28202_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16112 a_7037_60729# a_4351_55527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16113 a_17996_44007# a_16837_44219# a_17900_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16114 VSS a_3866_57399# a_5506_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16115 VDD a_1923_61759# a_1643_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16116 a_24490_61190# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16117 VDD config_2_in[0] a_1591_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X16118 a_9217_28879# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16119 a_11872_14191# a_10791_14191# a_11525_14433# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X1612 a_35730_47919# a_33423_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X16120 a_41348_48783# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16121 a_13151_23957# a_12463_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X16122 a_39154_62154# pmat.row_n[6] a_39646_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16123 VSS pmat.row_n[2] a_49590_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16124 a_43662_60508# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16125 VDD a_1586_8439# a_3247_6037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X16126 VDD a_38041_30485# a_38071_30838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16127 a_51294_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16128 a_37238_68178# a_18546_68220# a_37146_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16129 a_17619_43439# a_17442_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1613 VDD a_24775_50095# a_11067_64015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X16130 VSS a_35752_43781# a_35715_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16131 a_36234_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16132 VDD a_2867_43541# a_2411_43301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X16133 VDD _1192_.B1 a_23763_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16134 a_83005_26159# _1192_.B1 a_82787_26133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16135 a_20570_72556# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16136 VDD a_13763_67191# a_12597_68279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16137 a_12723_68367# a_10991_68591# a_12629_68367# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X16138 VDD pmat.rowon_n[9] a_19074_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16139 VDD VDD a_41162_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1614 VDD pmat.rowoff_n[7] a_20078_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16140 VDD a_8928_73865# a_9103_73791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16141 a_26498_58178# pmat.rowon_n[2] a_26102_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16142 VDD pmat.rowon_n[4] a_20078_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16143 VSS a_33957_48437# a_36265_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X16144 a_33622_71552# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16145 a_41558_67214# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16146 a_29606_61512# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16147 a_34134_8894# a_18162_8488# a_34226_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16148 a_29968_30083# a_25681_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16149 a_19470_20902# pmat.rowoff_n[12] a_19074_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1615 a_46578_12870# pmat.rowoff_n[4] a_46182_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16150 a_1761_2767# a_1591_2767# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16151 a_23486_7850# VDD a_23090_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16152 a_3434_51727# a_2676_51843# a_2871_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X16153 a_5331_28309# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X16154 a_77882_39738# a_77978_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16155 a_84090_3087# ANTENNA__1196__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16156 a_38546_23914# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16157 VSS a_7631_55687# a_3345_62839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16158 a_42166_15922# pmat.row_n[7] a_42658_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16159 a_45670_18496# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1616 a_4255_66959# a_4396_66933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X16160 a_45574_24918# VSS a_45178_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16161 VSS pmat.row_n[13] a_42562_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16162 a_39246_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16163 a_1959_12791# a_1979_12342# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16164 VSS pmat.row_n[10] a_31518_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16165 a_5221_45199# a_4745_45519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X16166 VSS a_7533_19087# a_7847_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16167 a_2744_25223# a_2952_25045# a_2886_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16168 a_11681_35823# a_11255_35862# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16169 a_5134_41909# a_4984_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X1617 a_44174_11906# pmat.row_n[3] a_44666_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16170 a_35534_16886# nmat.rowon_n[7] a_35138_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16171 a_24214_30287# a_24160_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X16172 a_2529_44409# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16173 a_47731_36103# a_40837_46261# a_47965_35951# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16174 a_28110_57134# a_18162_57174# a_28202_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16175 VDD a_2727_58470# a_4165_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X16176 a_32218_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16177 a_27498_32117# a_27340_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X16178 VDD a_4319_15039# a_4306_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16179 a_48586_15882# pmat.rowoff_n[7] a_48190_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1618 a_29510_64202# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16180 VDD nmat.rowon_n[5] a_22086_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16181 pmat.col_n[20] ANTENNA__1187__B1.DIODE a_39219_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16182 vcm a_18162_67214# a_36234_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16183 a_3841_15101# a_3797_14709# a_3675_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16184 a_11759_10615# a_10839_11989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X16185 a_43996_31599# a_42240_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X16186 a_36783_47158# a_36532_46805# a_36324_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16187 a_40250_65166# a_18546_65208# a_40158_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16188 a_6872_8725# a_1586_8439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16189 pmat.col[3] a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X1619 _1184_.A2 a_44888_33205# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u M=4
X16190 a_2672_23817# a_1591_23445# a_2325_23413# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16191 a_40650_69544# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16192 a_36234_55126# a_18546_55168# a_36142_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16193 a_24667_43177# a_25061_43132# a_11389_40443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X16194 a_32618_14480# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16195 vcm a_18162_66210# a_49286_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16196 a_36634_59504# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16197 a_3503_19087# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16198 a_6373_49249# a_6155_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X16199 a_30118_15922# a_18162_15516# a_30210_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X162 a_44570_72234# VDD a_44174_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1620 a_27106_21946# pmat.row_n[13] a_27598_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16200 a_33222_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16201 a_5602_11791# a_1717_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16202 VSS a_5497_73719# a_5445_73807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X16203 VSS a_6639_63927# a_4266_63303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16204 vcm a_18162_61190# a_50290_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16205 a_38242_7484# a_18546_7482# a_38150_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16206 VSS a_7840_27247# a_8292_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16207 a_49686_58500# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16208 VSS pmat.row_n[1] a_25494_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16209 a_19074_16926# pmat.row_n[8] a_19566_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1621 a_27106_17930# a_18162_17524# a_27198_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16210 vcm a_18162_9492# a_43262_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16211 a_28971_47753# a_28455_47381# a_28876_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X16212 a_6179_65479# a_5081_53135# a_6346_65577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X16213 a_36617_36603# a_34924_36165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X16214 VSS pmat.row_n[3] a_49590_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16215 a_20078_11906# pmat.row_n[3] a_20570_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16216 a_41162_65166# pmat.row_n[9] a_41654_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16217 a_27198_24552# a_18546_24550# a_27106_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16218 vcm a_18162_9492# a_19166_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16219 a_17478_46805# a_16800_47213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1622 VSS a_19488_52423# a_14287_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16220 a_26194_66170# a_18546_66212# a_26102_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16221 a_33130_10902# pmat.row_n[2] a_33622_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16222 a_14321_39958# a_14149_39747# a_14107_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X16223 VDD pmat.rowon_n[12] a_30118_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16224 a_17323_28111# a_7415_29397# a_17845_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16225 VDD pmat.rowon_n[2] a_26102_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16226 a_29206_9492# a_18546_9490# a_29114_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16227 VDD a_11207_31764# a_10764_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X16228 a_20451_47491# a_18823_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16229 a_26498_11866# nmat.rowon_n[12] a_26102_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1623 VDD nmat.rowon_n[9] a_33130_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16230 a_4314_19453# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16231 a_41558_20902# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16232 a_35630_9460# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16233 a_34611_42089# a_33489_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X16234 VSS a_4399_51157# a_5809_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16235 vcm a_18162_72234# a_31214_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16236 a_44174_56130# pmat.row_n[0] a_44666_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16237 a_35230_16520# a_18546_16518# a_35138_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16238 a_12353_19631# a_12311_19783# a_11892_21959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X16239 vcm a_18162_62194# a_27198_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1624 vcm a_18162_21540# a_48282_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16240 VSS a_34204_27765# a_34883_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16241 a_17959_41001# a_16837_40955# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16242 VSS a_13091_52047# a_16863_47428# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16243 a_27106_66170# pmat.row_n[10] a_27598_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16244 a_38546_64202# pmat.rowon_n[8] a_38150_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16245 a_31214_60146# a_18546_60188# a_31122_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16246 a_48282_15516# a_18546_15514# a_48190_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16247 VDD nmat.rowon_n[14] a_45178_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16248 VDD a_5423_69367# a_4265_71543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X16249 a_31614_64524# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1625 VSS a_12328_48168# a_12266_48285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X16250 VDD a_5497_62839# a_5785_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16251 vcm a_18162_12504# a_45270_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16252 VDD a_37519_46983# a_36539_47113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X16253 a_8820_6397# a_8703_6202# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16254 VDD nmat.rowon_n[2] a_36142_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16255 a_13533_71017# a_13327_70741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16256 a_46950_43719# a_46936_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16257 VSS a_7435_68021# a_5307_67655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X16258 a_39246_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16259 nmat.col_n[0] ANTENNA__1197__B.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1626 VDD a_4043_59861# a_1923_61759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X16260 a_21574_56492# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16261 a_39550_72234# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16262 VSS pmat.row_n[14] a_43566_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16263 a_43273_48463# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X16264 a_38905_28853# a_38727_32447# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16265 a_12002_49917# a_12044_49641# a_12002_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16266 a_22178_12504# a_18546_12502# a_22086_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16267 VDD a_2149_45717# a_2561_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16268 a_32126_60146# pmat.row_n[4] a_32618_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16269 vcm a_18162_11500# a_49286_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1627 VDD pmat.rowon_n[3] a_37146_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16270 a_41254_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16271 a_83090_26409# _1192_.A2 a_82787_26133# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16272 a_37238_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16273 VDD a_46130_34319# a_35244_32411# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16274 vcm.sky130_fd_sc_hd__buf_4_3.A vcm.sky130_fd_sc_hd__buf_4_2.A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16275 a_7896_11079# comp_latch a_8038_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16276 a_40467_46261# a_40837_46261# a_40694_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.624e+11p pd=2.1e+06u as=4.576e+11p ps=2.71e+06u w=640000u l=150000u
X16277 a_11115_71285# a_10190_60663# a_11058_62063# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X16278 a_25590_55488# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16279 VDD a_9675_10396# a_11759_10615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1628 a_23663_43177# a_23700_42919# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X16280 a_4341_65103# a_1591_65327# a_4259_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16281 vcm a_18162_23548# a_26194_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16282 a_20474_70226# pmat.rowon_n[14] a_20078_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16283 VSS pmat.row_n[5] a_46578_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16284 a_2464_67869# a_2250_67869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16285 a_43170_9898# a_18162_9492# a_43262_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16286 a_43566_17890# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16287 a_34552_44007# a_33489_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X16288 a_30210_21540# a_18546_21538# a_30118_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16289 a_5320_27023# a_4712_27023# a_5070_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1629 a_21797_47081# a_21837_46983# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X16290 a_50594_18894# nmat.rowon_n[5] a_50198_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16291 a_8569_60405# a_5651_66975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16292 a_14657_56873# a_11067_16359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16293 VSS pmat.row_n[15] a_29510_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16294 a_26194_11500# a_18546_11498# a_26102_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16295 VDD nmat.en_bit_n[1] a_34134_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16296 a_14646_19881# a_10239_14183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16297 a_27198_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16298 a_19074_9898# a_18162_9492# a_19166_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16299 cgen.dlycontrol1_in[4] a_1591_35951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X163 a_29114_64162# pmat.row_n[8] a_29606_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1630 a_31214_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16300 vcm a_18162_69222# a_51294_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16301 VDD a_6927_30503# a_11276_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16302 VSS pmat.row_n[2] a_25494_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16303 nmat.col_n[1] a_13354_2223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16304 a_8565_6037# a_8399_6037# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16305 vcm a_18162_59182# a_47278_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16306 a_15657_52317# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16307 a_5627_12879# a_5579_12394# a_5227_13077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16308 a_51294_57134# a_18546_57176# a_51202_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16309 VSS a_37820_30485# a_45911_36815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X1631 VSS a_5046_67655# a_3838_70455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16310 a_29206_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16311 a_23486_61190# pmat.rowon_n[5] a_23090_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16312 a_47582_16886# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16313 VDD a_40951_31599# a_45475_35520# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16314 a_38242_70186# a_18546_70228# a_38150_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16315 VSS pmat.row_n[6] a_51598_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16316 a_45178_10902# a_18162_10496# a_45270_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16317 a_2163_55233# a_1586_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16318 VSS a_6412_8725# a_6548_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+11p ps=1.6e+06u w=540000u l=150000u
X16319 a_35630_20504# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1632 a_51294_61150# a_18546_61192# a_51202_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16320 VDD VDD a_42166_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16321 a_35230_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16322 a_34134_18934# pmat.row_n[10] a_34626_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16323 VSS nmat.en_bit_n[1] a_34530_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16324 a_28110_20942# a_18162_20536# a_28202_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16325 a_35108_39655# a_33949_39867# a_35012_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16326 VDD pmat.rowon_n[6] a_38150_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16327 a_4831_40303# a_4705_39759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X16328 a_18546_16518# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X16329 a_24186_59142# a_18546_59184# a_24094_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1633 VSS pmat.row_n[1] a_23486_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X16330 a_2250_54991# a_2163_55233# a_1846_55123# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16331 VDD a_14825_50095# a_15210_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16332 a_2250_72221# a_2124_72123# a_1846_72107# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X16333 VSS a_7521_47081# a_9871_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X16334 a_25190_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16335 a_27502_60186# pmat.rowon_n[4] a_27106_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16336 a_27502_19898# nmat.rowon_n[4] a_27106_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16337 a_40951_31599# a_40678_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16338 VSS pmat.row_n[8] a_24490_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16339 a_2672_50095# a_1591_50095# a_2325_50337# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1634 a_35885_36165# a_36193_35805# a_11297_36091# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X16340 VSS a_36617_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X16341 a_22178_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16342 a_10381_16950# a_9528_20407# a_10167_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X16343 a_39154_70186# pmat.row_n[14] a_39646_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16344 a_36142_12910# a_18162_12504# a_36234_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16345 a_36538_7850# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16346 VSS a_11337_25071# a_14753_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16347 VSS pmat.row_n[13] a_36538_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16348 a_8381_46287# a_3746_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X16349 a_28202_58138# a_18546_58180# a_28110_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1635 a_34134_63158# a_18162_63198# a_34226_63158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16350 a_40554_67214# pmat.rowon_n[11] a_40158_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16351 vcm a_18162_55166# a_25190_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16352 VDD a_2529_44409# a_2559_44150# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16353 a_5597_67297# a_2419_53351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16354 a_49194_11906# a_18162_11500# a_49286_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16355 a_50290_18528# a_18546_18526# a_50198_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16356 a_25098_59142# pmat.row_n[3] a_25590_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16357 VSS a_13655_26703# a_14829_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16358 a_24573_49667# a_21371_50087# a_24501_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16359 VSS VDD a_46578_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1636 a_19470_56170# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16360 a_2847_26133# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16361 a_47767_30761# a_37291_29397# a_47685_30517# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16362 VDD a_18869_46831# a_19474_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16363 a_8908_14967# a_8305_20871# a_9050_15101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16364 a_37238_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16365 VDD pmat.rowoff_n[15] a_51202_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16366 VSS a_2972_9991# a_4249_9615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16367 a_37542_65206# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16368 a_30210_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16369 vcm a_18162_17524# a_20170_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1637 a_3408_11849# a_2327_11477# a_3061_11445# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16370 a_37638_17492# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16371 VDD a_34277_38550# a_34828_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16372 a_26194_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16373 a_27502_9858# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16374 vcm a_18162_14512# a_51294_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16375 VDD pmat.rowoff_n[7] a_41162_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16376 VDD ANTENNA__1190__A1.DIODE a_83094_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16377 a_2121_56623# a_1643_56597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16378 VDD a_3571_13627# a_12539_10389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X16379 a_48190_21946# pmat.row_n[13] a_48682_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1638 VSS a_8831_24501# a_8333_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.4365e+12p ps=1.222e+07u w=650000u l=150000u M=2
X16380 a_48190_17930# a_18162_17524# a_48282_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16381 VDD nmat.rowon_n[13] a_19074_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16382 a_4601_74005# a_4351_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.85e+11p pd=3.57e+06u as=0p ps=0u w=1e+06u l=150000u
X16383 a_34530_58178# pmat.rowon_n[2] a_34134_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16384 a_9405_28879# a_9217_28879# a_9323_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16385 a_8907_48437# a_9839_47679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16386 VSS a_11927_27399# a_22056_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16387 a_28704_29568# a_31399_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X16388 vcm a_18162_16520# a_24186_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16389 a_45270_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1639 a_21082_66170# a_18162_66210# a_21174_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16390 a_42166_66170# a_18162_66210# a_42258_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16391 a_47582_57174# pmat.rowon_n[1] a_47186_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16392 a_38150_13914# pmat.row_n[5] a_38642_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16393 a_48190_7890# a_18162_7484# a_48282_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16394 VSS a_22064_31287# a_20895_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16395 a_42658_11468# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16396 VSS pmat.row_n[8] a_27502_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16397 a_34924_41605# a_33765_41317# a_34828_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16398 VSS a_11019_71543# a_10969_71631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16399 a_6612_66933# a_3339_70759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X164 vcm a_18162_20536# a_51294_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1640 VDD a_33084_40743# a_32988_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X16400 a_11740_47197# a_11071_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16401 a_4679_28853# a_3351_27249# a_4898_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16402 a_28110_65166# a_18162_65206# a_28202_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16403 VDD a_10287_24759# a_9777_26935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X16404 a_19505_38779# a_17536_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16405 a_32218_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16406 a_2882_56989# a_2163_56765# a_2319_56860# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16407 VDD a_2648_29397# a_6559_8527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16408 a_32522_70226# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16409 a_14005_74953# a_12815_74581# a_13896_74953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1641 a_2215_47375# a_1775_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X16410 a_36234_63158# a_18546_63200# a_36142_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16411 VSS a_4135_19391# a_4069_19465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X16412 a_36634_67536# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16413 a_30118_23954# a_18162_23548# a_30210_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16414 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16415 VDD pmat.rowon_n[9] a_40158_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16416 a_46182_24958# VDD a_46674_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16417 VDD a_16911_51959# a_14839_66103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X16418 a_49286_62154# a_18546_62196# a_49194_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16419 a_14369_57711# a_11067_16359# a_14287_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1642 a_21574_11468# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16420 a_36142_57134# a_18162_57174# a_36234_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16421 a_50690_22512# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16422 a_49686_66532# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16423 a_22482_62194# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16424 a_12809_69679# a_12067_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16425 a_40250_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16426 a_19074_67174# a_18162_67214# a_19166_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16427 a_49194_56130# a_18162_56170# a_49286_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16428 VDD a_9675_10396# a_11249_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X16429 VSS pmat.row_n[14] a_36538_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1643 a_33526_9858# nmat.rowon_n[14] a_33130_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16430 a_35534_61190# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16431 a_37743_27497# a_34204_27765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16432 a_40650_14480# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16433 a_7436_16519# a_7644_16341# a_7578_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16434 a_40554_20902# pmat.rowoff_n[12] a_40158_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16435 a_23741_42567# a_22817_41317# a_23939_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16436 VDD a_11731_8751# a_12133_9001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X16437 vcm a_18162_71230# a_23182_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16438 a_33715_48783# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16439 VDD pmat.rowon_n[0] a_43170_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1644 a_6829_49007# a_5639_49007# a_6720_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X16440 a_3476_59343# a_3262_59343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16441 a_23582_24520# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16442 a_12889_64789# a_12723_64789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16443 VDD pmat.rowon_n[10] a_26102_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16444 a_51202_14918# a_18162_14512# a_51294_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16445 a_26194_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16446 a_33222_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16447 VDD a_2648_29397# a_4815_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16448 VSS a_31675_47695# a_43267_47081# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16449 a_12437_74281# a_12225_74575# a_6292_65479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1645 a_13563_24527# a_12463_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.344e+11p pd=1.48e+06u as=0p ps=0u w=420000u l=150000u
X16450 VDD a_4516_21531# a_6579_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X16451 a_43533_30761# a_28336_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16452 a_35230_24552# a_18546_24550# a_35138_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16453 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16454 a_10167_16950# a_9528_20407# a_10167_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16455 a_41162_10902# pmat.row_n[2] a_41654_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16456 vcm a_18162_70226# a_27198_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16457 VDD nmat.rowon_n[15] a_21082_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16458 vcm a_18162_9492# a_51294_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16459 VDD a_12069_36341# a_12013_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1646 a_10601_65103# a_5651_66975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16460 VDD VSS a_47186_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16461 a_38546_72234# VDD a_38150_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16462 a_24094_20942# pmat.row_n[12] a_24586_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16463 a_31614_72556# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16464 a_24094_16926# a_18162_16520# a_24186_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16465 vcm a_18162_20536# a_45270_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16466 a_48282_23548# a_18546_23546# a_48190_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16467 a_14486_48169# a_11067_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16468 VDD pmat.rowon_n[2] a_34134_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16469 a_27598_62516# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1647 cgen.dlycontrol2_in[2] a_1591_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16470 VDD a_15543_31573# a_15530_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16471 VDD pmat.rowon_n[4] a_31122_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16472 a_31122_62154# a_18162_62194# a_31214_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16473 a_34530_11866# nmat.rowon_n[12] a_34134_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16474 a_76962_39738# a_77058_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16475 VDD a_2319_65564# a_2250_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16476 VSS a_28131_50069# pmat.col[8] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16477 a_21970_48071# a_20475_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16478 nmat.col[28] _1194_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16479 a_47582_10862# nmat.rowon_n[13] a_47186_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1648 a_34626_10464# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16480 a_31117_27791# a_21739_29415# nmat.col_n[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X16481 VDD a_37497_38550# a_37404_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16482 VSS a_34204_27765# a_36723_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16483 a_1979_11254# a_1761_9839# a_1907_11254# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X16484 a_2743_38279# a_2839_38101# a_3141_38127# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X16485 a_42562_59182# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16486 a_22178_20536# a_18546_20534# a_22086_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16487 a_4865_8181# a_4503_6335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16488 a_5779_71285# a_8283_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X16489 a_40158_16926# pmat.row_n[8] a_40650_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1649 VDD a_11521_64239# a_11867_64899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16490 a_25494_69222# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16491 a_19487_49159# a_19759_48987# a_19717_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16492 a_20063_30877# a_19439_30511# a_19955_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16493 VSS a_3615_71631# a_14365_68743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16494 a_9217_23983# a_8831_24501# a_9135_23983# VSS sky130_fd_pr__nfet_01v8 ad=1.8525e+11p pd=1.87e+06u as=0p ps=0u w=650000u l=150000u
X16495 a_36288_44527# a_36111_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16496 a_8937_15823# a_8767_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16497 VSS a_26475_34343# a_11057_35836# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16498 VSS a_36801_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X16499 a_14778_26409# a_8861_24527# a_14696_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X165 a_33622_62516# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1650 a_4707_32156# a_1781_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16500 VDD a_29163_38545# a_29023_38571# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16501 a_3591_62927# a_2215_47375# a_3495_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16502 a_46578_58178# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16503 VSS a_8695_12801# a_8656_12675# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16504 a_25190_61150# a_18546_61192# a_25098_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16505 a_46578_16886# nmat.rowon_n[7] a_46182_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16506 a_29510_68218# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16507 a_42258_8488# a_18546_8486# a_42166_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16508 a_6339_40303# a_5823_40303# a_6244_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X16509 a_21239_50613# a_21395_50857# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X1651 a_6833_37281# a_6615_37039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X16510 VSS a_34204_27765# a_34148_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16511 VDD nmat.rowon_n[5] a_33130_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16512 a_43132_48071# a_43267_47081# a_43274_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16513 vcm a_18162_67214# a_47278_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16514 a_46023_32937# a_43533_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16515 a_9184_51335# a_9457_51163# a_9415_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16516 a_51294_65166# a_18546_65208# a_51202_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16517 a_51694_69544# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16518 VDD a_13909_39605# a_14321_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16519 a_47278_55126# a_18546_55168# a_47186_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1652 a_25647_38695# a_25755_38695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X16520 a_47678_59504# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16521 a_83170_5263# ANTENNA__1190__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16522 VSS pmat.row_n[2] a_23486_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16523 a_12449_22895# a_12247_20175# a_12533_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X16524 a_51202_59142# a_18162_59182# a_51294_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16525 VSS a_13503_36893# a_13443_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16526 a_26102_61150# pmat.row_n[5] a_26594_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16527 a_35230_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16528 a_8744_71689# a_7829_71317# a_8397_71285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X16529 a_6173_6575# a_5654_9527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1653 a_6559_8527# a_5654_9527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X16530 a_34134_69182# a_18162_69222# a_34226_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16531 a_22925_28111# a_13091_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16532 VDD pmat.rowon_n[14] a_38150_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16533 a_39193_43131# a_37960_42693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16534 a_51202_9898# a_18162_9492# a_51294_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16535 a_24186_67174# a_18546_67216# a_24094_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16536 VSS nmat.rowon_n[14] a_19793_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16537 a_42987_50345# a_28131_50069# a_42769_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16538 VSS a_1586_50247# a_7479_53909# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16539 a_38242_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1654 a_10216_62985# a_9135_62613# a_9869_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16540 a_12646_51549# a_12520_51451# a_12242_51435# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X16541 a_42258_17524# a_18546_17522# a_42166_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16542 a_31021_28585# a_21365_27247# a_30699_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16543 a_7005_75983# a_6799_75637# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16544 a_3978_48071# a_3987_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16545 VSS a_12069_36341# a_12013_36694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16546 VSS a_6467_29415# a_14249_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16547 a_36142_20942# a_18162_20536# a_36234_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16548 a_43351_31599# a_41949_30761# a_42307_31756# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16549 cgen.enable_dlycontrol_in a_1591_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1655 a_44266_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16550 a_42166_57134# pmat.row_n[1] a_42658_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16551 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16552 vcm a_18162_63198# a_25190_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16553 a_25098_67174# pmat.row_n[11] a_25590_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16554 a_36538_65206# pmat.rowon_n[9] a_36142_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16555 a_46274_16520# a_18546_16518# a_46182_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16556 VDD a_11927_27399# a_12403_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16557 vcm a_18162_13508# a_43262_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16558 a_14371_25071# a_9441_20189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X16559 VSS a_2563_34837# a_4535_38377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1656 VDD a_9668_10651# a_10897_6825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X16560 a_6087_67655# a_5081_53135# a_6254_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X16561 a_35353_50639# _1154_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16562 VSS pmat.row_n[7] a_45574_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16563 a_42562_12870# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16564 VDD ANTENNA__1196__A2.DIODE a_47764_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16565 a_25494_22910# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16566 a_32522_23914# pmat.rowoff_n[15] a_32126_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16567 a_6087_67655# a_2879_57487# a_6432_67503# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X16568 VSS a_5131_13255# a_5081_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16569 a_19166_18528# a_18546_18526# a_19074_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1657 VDD a_1923_69823# a_2464_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X16570 a_9301_62613# a_9135_62613# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16571 a_41786_28111# a_18243_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16572 a_32618_56492# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16573 a_47212_29673# a_37291_29397# a_47126_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16574 a_30329_42689# a_29627_43983# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16575 result_out[7] a_1644_64213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X16576 a_46182_58138# pmat.row_n[2] a_46674_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16577 a_22482_15882# pmat.rowoff_n[7] a_22086_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16578 a_2464_31965# a_2250_31965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16579 a_36617_37691# a_36161_37462# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1658 VSS pmat.row_n[12] a_32522_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X16580 a_1644_60949# a_1823_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16581 a_46578_11866# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16582 VSS comp.adc_comp_circuit_0.adc_comp_buffer_0.in a_54790_39936# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.55e+11p ps=1.62e+06u w=500000u l=150000u
X16583 a_19965_36603# a_17996_36391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16584 VDD a_11525_14433# a_11415_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16585 a_29510_21906# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16586 vcm a_18162_24552# a_24186_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16587 VSS a_13837_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X16588 VSS a_11067_30287# a_25221_46519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16589 a_11200_42717# a_10949_42364# a_10979_42390# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1659 a_39469_38053# a_37776_37479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16590 VSS pmat.row_n[6] a_44570_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16591 a_47582_9858# nmat.rowon_n[14] a_47186_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16592 vcm a_18162_56170# a_19166_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16593 VSS VDD a_27502_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16594 a_18546_57176# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X16595 VDD a_20411_51157# a_14653_53458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16596 a_31518_70226# pmat.rowon_n[14] a_31122_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16597 a_23582_58500# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16598 a_19470_13874# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16599 a_16324_36911# a_16147_36911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X166 vcm a_18162_10496# a_47278_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1660 a_43170_19938# pmat.row_n[11] a_43662_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16600 VDD a_9528_20407# a_12461_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16601 VSS pmat.row_n[3] a_23486_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16602 VSS pmat.rowon_n[7] pmat.rowoff_n[12] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X16603 a_13717_5263# a_10883_3303# nmat.col[10] VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X16604 VDD VSS a_45178_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16605 a_23939_41271# a_22817_41317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16606 VDD a_6830_22895# a_12437_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16607 a_21478_62194# pmat.rowon_n[6] a_21082_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16608 a_10097_15279# a_10053_15521# a_9931_15279# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X16609 VSS a_4337_22351# a_5271_23447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1661 a_22988_47741# a_22276_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X16610 a_23442_32143# a_22365_32149# a_23280_32521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16611 VSS pmat.row_n[8] a_35534_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16612 a_21215_48071# a_28901_48437# a_28849_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16613 result_out[2] a_1644_56053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16614 a_49286_70186# a_18546_70228# a_49194_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16615 VDD a_2648_29397# a_10381_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16616 a_36142_65166# a_18162_65206# a_36234_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16617 VDD pmat.rowoff_n[15] a_49194_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16618 a_40250_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16619 a_46674_20504# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1662 VSS a_9303_22351# a_10097_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X16620 VSS a_45866_38279# a_46513_39009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16621 a_46274_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16622 a_6343_18517# a_6168_18543# a_6522_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16623 VSS a_15667_27239# a_45279_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16624 a_33141_51727# _1184_.A2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16625 a_20078_70186# a_18162_70226# a_20170_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16626 a_49194_64162# a_18162_64202# a_49286_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16627 a_12269_8207# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16628 a_30641_44743# a_30913_44219# a_31976_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16629 a_40554_8854# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1663 a_45670_56492# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16630 a_44666_8456# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16631 a_30181_37253# a_30489_36893# a_30155_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X16632 VDD a_24867_53135# a_40685_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16633 VDD pmat.rowoff_n[7] a_39154_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16634 VDD a_3339_59879# a_11112_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16635 a_5275_65327# a_5399_65479# a_5138_65479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16636 a_36634_12472# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16637 VDD nmat.rowon_n[13] a_40158_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16638 a_19566_22512# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16639 a_19611_27247# a_6829_26703# a_19522_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1664 VSS a_28704_29568# a_41703_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X16640 pmat.rowon_n[3] a_10239_14183# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X16641 a_51202_22950# a_18162_22544# a_51294_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16642 VDD pmat.rowoff_n[12] a_23090_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16643 a_47186_12910# a_18162_12504# a_47278_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16644 VDD a_40105_47375# a_46013_42997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16645 a_26194_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16646 a_23090_61150# a_18162_61190# a_23182_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16647 VSS pmat.row_n[13] a_47582_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16648 VSS pmat.row_n[0] a_26498_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16649 a_5462_57711# a_4351_55527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1665 VSS a_47207_35951# a_47453_36815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16650 a_51598_67214# pmat.rowon_n[11] a_51202_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16651 a_4038_22717# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16652 a_26498_71230# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16653 VDD config_1_in[1] a_1591_9839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X16654 VDD a_5351_19913# a_9339_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X16655 a_3149_40303# a_2419_69455# a_2931_40277# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16656 a_24094_24958# a_18162_24552# a_24186_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16657 a_33765_39141# a_32072_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16658 VDD pmat.rowon_n[10] a_34134_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16659 a_2847_33749# a_2672_33775# a_3026_33775# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1666 a_47278_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16660 VSS cgen.dlycontrol2_in[0] a_28431_34735# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X16661 a_27598_70548# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16662 a_41558_59182# pmat.rowon_n[3] a_41162_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16663 VDD a_2325_23413# a_2215_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16664 VSS a_12133_9001# a_12257_8527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16665 VSS a_35186_47375# a_37649_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16666 a_24186_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16667 a_27106_60146# a_18162_60186# a_27198_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16668 a_7444_9117# a_7176_8751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.89e+11p pd=1.74e+06u as=0p ps=0u w=420000u l=150000u
X16669 a_48586_65206# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1667 a_28202_62154# a_18546_62196# a_28110_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16670 VDD a_2935_38279# a_6920_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16671 VSS pmat.row_n[5] a_20474_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16672 a_2507_29673# a_2422_29575# a_2289_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16673 a_12266_48285# a_11547_48061# a_11703_48156# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16674 a_33327_52521# a_24591_28327# a_33109_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16675 a_14745_29423# a_14691_29575# a_14649_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16676 a_31518_24918# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16677 a_14460_60137# nmat.rowon_n[7] a_14287_59887# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16678 a_12371_57487# a_12341_57141# a_5682_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X16679 a_38546_57174# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1668 a_40554_71230# pmat.rowon_n[15] a_40158_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16680 a_35630_62516# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16681 a_29053_31375# a_22628_30485# a_28803_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16682 VSS a_25325_29125# a_25315_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16683 ctopp clk_ena ctopp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u M=2
X16684 a_40158_67174# a_18162_67214# a_40250_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16685 a_45574_58178# pmat.rowon_n[2] a_45178_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16686 VSS VDD a_42562_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16687 vcm a_18162_59182# a_21174_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16688 a_14460_11177# a_10239_14183# a_14369_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16689 a_28110_8894# a_18162_8488# a_28202_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1669 VSS a_3325_26159# a_4259_24643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X16690 a_10443_12879# a_10471_12791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X16691 a_23090_7890# VDD a_23582_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16692 a_28506_68218# pmat.rowon_n[12] a_28110_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16693 a_48682_61512# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16694 vcm a_18162_16520# a_35230_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16695 a_21478_16886# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16696 a_6733_45199# a_4399_51157# a_5921_44629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16697 a_39646_19500# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16698 VSS ANTENNA__1395__B1.DIODE a_22925_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16699 a_44733_44431# a_31675_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X167 a_2847_63999# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1670 a_4121_66237# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16700 a_34530_15882# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16701 _1224_.X a_82863_64213# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=8
X16702 VSS a_27049_35515# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X16703 a_23648_47753# a_22733_47381# a_23301_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X16704 a_4748_34319# a_4227_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16705 VDD pmat.rowon_n[5] a_25098_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16706 VDD a_4491_53511# a_4123_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16707 a_2743_38279# a_2935_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16708 a_9779_26819# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16709 a_10953_41605# a_11261_41245# a_10927_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1671 a_28602_66532# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16710 a_4135_37815# a_4127_37013# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16711 a_7037_60729# a_4351_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16712 VSS pmat.row_n[10] a_50594_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16713 VSS a_10383_75637# a_6795_76989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16714 a_47278_63158# a_18546_63200# a_47186_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16715 VDD a_34277_37462# a_34828_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16716 a_47678_67536# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16717 a_20474_63198# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16718 VDD pmat.rowon_n[9] a_51202_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16719 a_17336_43439# a_17159_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1672 a_25098_63158# pmat.row_n[7] a_25590_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16720 a_47186_57134# a_18162_57174# a_47278_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16721 a_15368_31599# a_14453_31599# a_15021_31841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16722 a_14391_26703# a_12987_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16723 VDD a_10047_8751# a_10379_8439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16724 a_7589_33749# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16725 VDD a_21031_37217# a_20855_36885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X16726 a_33526_62194# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16727 a_51294_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16728 a_25287_32117# a_11067_30287# a_25505_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X16729 a_3868_33609# a_2953_33237# a_3521_33205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1673 a_20078_8894# pmat.row_n[0] a_20570_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16730 VDD pmat.rowon_n[4] a_29114_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16731 VDD pmat.rowon_n[1] a_41162_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16732 VSS a_8723_67191# a_7899_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16733 VSS pmat.row_n[14] a_47582_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16734 a_12934_35823# a_12757_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16735 a_51694_14480# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16736 a_51598_20902# pmat.rowoff_n[12] a_51202_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16737 VDD a_12038_55687# a_11835_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X16738 a_50290_8488# a_18546_8486# a_50198_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16739 a_13776_37455# a_11497_38543# a_13555_37782# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1674 a_50290_22544# a_18546_22542# a_50198_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16740 VSS vcm.sky130_fd_sc_hd__buf_4_0.A a_77428_40594# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16741 a_5687_71829# a_12131_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X16742 a_34626_24520# nmat.en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16743 VDD a_10190_60663# a_10141_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16744 a_15585_29199# a_14691_29575# a_15489_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16745 a_24186_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16746 VSS _1187_.A2 a_28725_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16747 a_6612_65845# a_3339_70759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16748 VSS a_2835_13077# a_12397_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16749 a_41558_12870# pmat.rowoff_n[4] a_41162_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1675 a_12809_69679# a_12152_66415# a_12821_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16750 a_2250_67869# a_2163_67645# a_1846_67755# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16751 a_24490_64202# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16752 a_38150_55126# VDD a_38642_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16753 VDD a_10286_60405# a_10975_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16754 a_22086_21946# pmat.row_n[13] a_22578_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16755 a_46274_24552# a_18546_24550# a_46182_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16756 a_22086_17930# a_18162_17524# a_22178_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16757 vcm a_18162_21540# a_43262_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16758 a_45270_66170# a_18546_66212# a_45178_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16759 a_16111_40183# a_16505_40157# a_16171_40157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X1676 a_11530_77661# a_10811_77437# a_10967_77532# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X16760 pmat.row_n[11] a_10055_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16761 a_35138_20942# pmat.row_n[12] a_35630_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16762 a_50594_68218# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16763 a_35138_16926# a_18162_16520# a_35230_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16764 a_46481_52271# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16765 a_17996_36391# a_16837_36603# a_17900_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16766 VDD pmat.rowon_n[2] a_45178_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16767 a_38546_10862# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16768 a_14150_54991# a_13073_54997# a_13988_55369# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X16769 a_45574_11866# nmat.rowon_n[12] a_45178_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1677 VDD pmat.rowon_n[8] a_32126_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16770 VSS a_13467_21263# a_13768_22325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16771 VSS a_7717_14735# a_36453_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16772 a_28602_15484# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16773 a_28506_21906# nmat.rowon_n[2] a_28110_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16774 VSS a_3225_55509# a_2840_55509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16775 a_25098_12910# pmat.row_n[4] a_25590_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16776 VDD nmat.rowon_n[10] a_32126_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16777 VSS a_10239_77295# a_11077_76207# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16778 a_31015_29111# a_21365_27247# a_31249_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16779 vcm a_18162_62194# a_46274_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1678 VDD a_4351_55527# a_5402_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X16780 a_46182_66170# pmat.row_n[10] a_46674_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16781 a_9282_56445# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16782 a_50290_60146# a_18546_60188# a_50198_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16783 VSS a_29051_39783# a_12345_39100# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16784 vcm.sky130_fd_sc_hd__buf_4_0.A vcm.sky130_fd_sc_hd__dlymetal6s6s_1_3.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16785 a_50690_64524# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16786 a_35802_27791# a_25695_28111# a_35499_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16787 pmat.row_n[15] a_17191_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16788 a_27106_9898# pmat.row_n[1] a_27598_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16789 a_2529_44409# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1679 a_46274_12504# a_18546_12502# a_46182_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16790 VDD a_2325_50337# a_2215_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16791 a_39473_40517# a_39781_40157# a_12309_38659# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X16792 a_29189_47349# a_28971_47753# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X16793 a_10147_29415# pmat.sw a_36541_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16794 a_38150_72194# a_18162_72234# a_38242_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16795 vcm a_18162_64202# a_19166_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16796 a_40650_56492# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16797 a_29114_11906# pmat.row_n[3] a_29606_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16798 a_19074_68178# pmat.row_n[12] a_19566_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16799 a_42258_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X168 a_38150_60146# a_18162_60186# a_38242_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1680 a_29404_44869# a_28245_44581# a_29308_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X16800 a_18546_65208# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X16801 a_23182_62154# a_18546_62196# a_23090_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16802 a_23582_66532# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16803 a_20078_63158# pmat.row_n[7] a_20570_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16804 a_22178_9492# a_18546_9490# a_22086_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16805 a_41254_12504# a_18546_12502# a_41162_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16806 VSS a_8695_63937# a_8656_63811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16807 a_31976_44007# a_30913_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16808 a_51202_60146# pmat.row_n[4] a_51694_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16809 vcm a_18162_68218# a_45270_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1681 a_8413_12925# a_8378_12691# a_8175_12533# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16810 a_14486_47081# a_11067_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16811 VDD a_4075_50087# a_4627_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X16812 a_6641_8527# a_5654_9527# a_6559_8527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16813 VSS a_1899_35051# a_1775_35113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16814 a_12757_40214# a_12585_40443# a_12543_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16815 cgen.dlycontrol3_in[3] a_2235_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16816 VSS VDD a_35534_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16817 nmat.col[3] _1194_.A2 a_12999_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16818 a_12237_60431# a_10049_60663# a_11797_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16819 a_2847_18303# a_2672_18377# a_3026_18365# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1682 a_37238_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16820 VDD a_2315_44124# a_4075_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16821 a_24094_62154# pmat.row_n[6] a_24586_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16822 a_3641_72765# a_3262_72399# a_3569_72765# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16823 VDD a_36161_37462# a_37404_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16824 VSS pmat.row_n[15] a_48586_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16825 a_12132_58621# a_5535_57993# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16826 VSS pmat.row_n[2] a_34530_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16827 a_45270_11500# a_18546_11498# a_45178_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16828 a_10378_62607# a_9301_62613# a_10216_62985# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16829 a_22178_68178# a_18546_68220# a_22086_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1683 a_48282_9492# a_18546_9490# a_48190_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16830 a_49590_8854# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16831 a_43170_21946# a_18162_21540# a_43262_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16832 a_46274_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16833 VSS a_2871_51701# a_2802_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16834 a_5498_56399# a_4351_55527# a_5408_56399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16835 a_2193_11254# a_2021_11043# a_1979_11254# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X16836 a_28110_19938# pmat.row_n[11] a_28602_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16837 a_24937_36039# a_24565_34789# a_25628_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16838 a_19491_47893# a_19647_48052# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X16839 a_49286_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1684 VSS a_12651_35823# a_12757_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16840 a_4357_9295# a_2972_9991# a_4167_9615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X16841 a_42562_61190# pmat.rowon_n[5] a_42166_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16842 a_37463_38007# a_36341_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16843 a_25494_71230# pmat.rowon_n[15] a_25098_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16844 a_7079_40277# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16845 a_28629_48437# a_28901_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16846 a_8507_20175# a_8256_20291# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16847 a_2121_31599# a_1643_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16848 VDD a_24867_53135# a_36545_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16849 a_50594_21906# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1685 VDD cgen.dlycontrol4_in[4] a_30819_40191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16850 a_47186_20942# a_18162_20536# a_47278_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16851 VSS a_2411_33749# a_2369_39037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16852 a_43262_59142# a_18546_59184# a_43170_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16853 vcm a_18162_56170# a_40250_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16854 VSS a_12345_39100# a_24895_38517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16855 VSS a_7072_62037# a_5595_65301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X16856 VDD a_20787_30199# a_20591_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X16857 a_39550_18894# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16858 VSS a_11948_49783# a_38569_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16859 a_13139_54599# a_12895_53359# a_13537_54447# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X1686 a_28629_48437# a_28901_48437# a_29300_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.05e+11p ps=7.61e+06u w=1e+06u l=150000u M=2
X16860 VSS pmat.row_n[8] a_43566_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16861 a_40554_13874# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16862 a_29510_70226# pmat.rowon_n[14] a_29114_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16863 VDD a_10932_21959# a_10814_29111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X16864 a_41254_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16865 a_23486_23914# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16866 VDD a_4809_13621# a_4699_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16867 a_14369_21807# a_5351_19913# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16868 VSS a_4768_16055# a_4215_15797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16869 a_30610_18496# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1687 VSS a_13575_68743# a_13279_68841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X16870 a_30514_24918# VSS a_30118_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16871 a_20787_30199# clk_ena a_20961_30305# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16872 a_24186_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16873 a_34553_42658# a_33489_43131# a_34552_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16874 a_8891_66964# a_9405_66627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X16875 a_22178_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16876 a_6334_69679# a_5779_71285# a_6524_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16877 vcm a_18162_55166# a_44266_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16878 a_19470_62194# pmat.rowon_n[6] a_19074_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16879 a_2080_59165# a_1643_58773# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1688 VDD pmat.rowon_n[0] a_22086_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16880 a_44174_59142# pmat.row_n[3] a_44666_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16881 VDD a_11921_37462# a_10985_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X16882 a_39193_42043# a_38737_41814# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X16883 nmat.rowon_n[10] a_14458_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16884 a_2882_31965# a_2163_31741# a_2319_31836# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16885 a_20474_16886# nmat.rowon_n[7] a_20078_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16886 VSS pmat.row_n[9] a_29510_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16887 a_35630_70548# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16888 a_33526_15882# pmat.rowoff_n[7] a_33130_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16889 VSS pmat.row_n[7] a_42562_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1689 a_8507_20175# a_8256_20291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X16890 VDD a_14943_26703# a_17136_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16891 vcm a_18162_67214# a_21174_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16892 a_39246_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16893 VDD a_24719_38517# a_14773_39394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16894 a_21174_55126# a_18546_55168# a_21082_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16895 vcm a_18162_24552# a_35230_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16896 a_3262_59343# a_3175_59585# a_2858_59475# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X16897 vcm a_18162_66210# a_34226_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16898 a_45270_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16899 a_11965_42583# a_12061_42325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X169 a_46339_31029# a_47011_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u M=3
X1690 a_44570_70226# pmat.rowon_n[14] a_44174_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16900 a_21574_59504# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16901 a_20179_40719# a_19925_41046# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16902 a_37960_42693# a_36801_42405# a_37864_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16903 VDD a_6895_48981# a_6882_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16904 a_38242_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16905 a_34626_58500# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16906 VSS a_16311_28327# a_26329_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16907 a_2847_50069# a_2672_50095# a_3026_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16908 VSS pmat.row_n[3] a_34530_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16909 a_4853_28335# a_4809_28577# a_4687_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1691 a_29114_62154# pmat.row_n[6] a_29606_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16910 VSS a_2100_44343# a_2051_44111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16911 a_4520_60975# a_4041_61225# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X16912 a_55578_39250# comp.adc_nor_latch_0.R ndecision_finish VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16913 a_23707_40693# a_12228_40693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16914 a_12967_12863# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16915 VDD VDD a_43170_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16916 VSS a_15667_27239# a_45556_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16917 a_8333_24847# a_6829_26703# a_8861_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16918 a_49590_67214# pmat.rowon_n[11] a_49194_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16919 VSS pmat.row_n[8] a_46578_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1692 a_33622_60508# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16920 a_22628_30485# a_22871_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16921 a_33685_48437# a_33957_48437# a_34356_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X16922 VDD VDD a_19074_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16923 a_44666_21508# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16924 VSS a_13837_39069# a_13529_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16925 a_44266_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16926 a_31122_7890# VDD a_31614_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16927 a_47186_65166# a_18162_65206# a_47278_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16928 VSS a_31539_51946# pmat.col[0] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X16929 a_51294_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1693 VDD a_13641_23439# a_33870_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X16930 a_20474_9858# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16931 VSS a_3325_20175# a_4811_22351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X16932 a_39550_59182# pmat.rowon_n[3] a_39154_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16933 a_14461_48463# a_12044_49641# a_13688_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16934 VSS pmat.row_n[0] a_36538_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16935 a_25494_7850# VDD a_25098_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16936 a_28442_29199# a_27794_28879# a_28273_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16937 a_20170_16520# a_18546_16518# a_20078_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16938 a_21371_50087# a_45238_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16939 VDD nmat.rowon_n[7] a_37146_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1694 a_9367_50871# a_8385_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X16940 a_34552_36391# a_33489_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16941 VSS pmat.row_n[10] a_19470_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16942 a_51598_70226# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16943 vcm a_18162_17524# a_29206_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16944 a_12585_40443# a_15549_39867# a_16612_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16945 a_23486_64202# pmat.rowon_n[8] a_23090_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16946 a_33222_15516# a_18546_15514# a_33130_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16947 vcm a_18162_12504# a_30210_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16948 VDD a_2163_58941# a_2124_59067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X16949 a_10139_32117# a_9944_32259# a_10449_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X1695 VSS a_20439_27247# a_33925_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16950 a_47678_12472# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16951 VDD nmat.rowon_n[2] a_21082_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16952 VSS a_10839_11989# a_12253_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16953 a_45178_13914# a_18162_13508# a_45270_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16954 VDD nmat.rowon_n[13] a_51202_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16955 a_24186_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16956 VSS a_9103_56383# a_9037_56457# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X16957 a_41558_62194# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16958 VDD a_19459_35279# a_19565_35279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16959 a_8452_65149# a_5307_67655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1696 a_27198_68178# a_18546_68220# a_27106_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16960 a_24490_72234# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16961 a_11697_56775# a_6787_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X16962 a_9749_19061# a_3688_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X16963 vcm a_18162_71230# a_42258_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16964 vcm a_18162_11500# a_34226_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16965 vcm a_18162_61190# a_38242_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16966 a_22178_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16967 a_35138_24958# a_18162_24552# a_35230_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16968 VDD pmat.rowon_n[10] a_45178_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16969 a_42658_63520# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1697 a_48190_21946# a_18162_21540# a_48282_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16970 a_8121_49257# a_8267_49159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16971 a_27198_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16972 VSS a_27498_32117# a_27976_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16973 a_45270_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16974 a_41699_52521# a_18243_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16975 VSS pmat.row_n[5] a_31518_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16976 a_28202_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16977 vcm a_18162_9492# a_45270_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16978 a_26515_38007# a_25393_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X16979 a_12013_47919# a_11634_48285# a_11941_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1698 a_18235_42359# a_18272_42693# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X16980 vcm a_18162_70226# a_46274_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16981 a_10515_75895# a_11014_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16982 VDD a_8919_71615# a_8906_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16983 VDD nmat.rowon_n[12] a_28110_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16984 VDD ANTENNA__1197__A.DIODE a_45747_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16985 a_13144_65149# a_5462_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16986 a_33049_27497# a_25879_31591# nmat.col_n[11] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X16987 a_50690_72556# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16988 VDD pmat.rowon_n[9] a_49194_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16989 a_46674_62516# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1699 pmat.row_n[2] a_23815_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16990 a_9766_8207# a_9731_8439# a_9463_8439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X16991 a_35277_30333# a_35242_30099# a_35039_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16992 result_out[9] a_1644_66933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16993 VDD pmat.rowon_n[4] a_50198_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16994 vcm a_18162_59182# a_32218_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16995 VDD a_11067_27239# a_37927_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16996 a_5699_32687# a_5253_32687# a_5603_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16997 a_26552_43781# a_25393_43493# a_26515_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16998 a_5134_41909# a_4984_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.21e+06u as=0p ps=0u w=840000u l=150000u
X16999 vcm a_18162_72234# a_19166_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_51598_55166# VSS a_51202_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X170 a_26456_43781# a_26552_43781# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X1700 a_8851_12533# a_8656_12675# a_9161_12925# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X17000 VDD a_1769_47919# a_3707_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X17001 a_32522_16886# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17002 VSS a_29220_37253# a_29183_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X17003 a_4498_15101# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17004 a_9873_74031# a_9831_74183# a_7099_74313# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X17005 a_23182_70186# a_18546_70228# a_23090_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17006 VDD pmat.rowon_n[1] a_39154_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17007 a_3763_6409# a_3413_6037# a_3668_6397# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X17008 a_30118_10902# a_18162_10496# a_30210_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17009 a_10139_32117# a_9983_32385# a_10284_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X1701 a_34530_62194# pmat.rowon_n[6] a_34134_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17010 a_20078_71190# pmat.row_n[15] a_20570_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17011 a_19166_60146# a_18546_60188# a_19074_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17012 vcm a_18162_22544# a_37238_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17013 a_49590_20902# pmat.rowoff_n[12] a_49194_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17014 a_20570_20504# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17015 a_19566_64524# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17016 a_20170_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17017 a_41254_20536# a_18546_20534# a_41162_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17018 a_28705_39141# a_28116_38567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17019 a_2557_69679# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1702 a_12257_8527# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17020 VDD pmat.rowon_n[6] a_23090_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17021 a_37238_10496# a_18546_10494# a_37146_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17022 a_44570_69222# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17023 a_5185_10089# a_2972_9991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17024 VDD nmat.rowon_n[14] a_47186_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17025 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17026 a_10287_24759# a_5351_19913# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17027 VSS a_44976_47349# a_44870_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X17028 a_39550_12870# pmat.rowoff_n[4] a_39154_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17029 a_4601_35727# a_4267_35407# a_4517_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X1703 a_7605_63401# a_7563_63303# a_7509_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X17030 a_1770_35015# a_2467_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17031 a_45064_44807# a_44966_43255# a_45295_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17032 a_29493_31375# a_29635_31029# a_28803_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17033 a_24094_70186# pmat.row_n[14] a_24586_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17034 a_45178_58138# a_18162_58178# a_45270_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17035 a_26456_43781# a_25393_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17036 a_21082_12910# a_18162_12504# a_21174_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17037 a_28110_68178# a_18162_68218# a_28202_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17038 VSS pmat.row_n[13] a_21478_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17039 a_6641_47375# a_5566_44905# a_6553_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1704 VSS a_24921_27221# nmat.col_n[5] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17040 a_47893_35951# a_47207_35951# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17041 a_14471_3561# _1184_.A2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17042 a_45178_17930# pmat.row_n[9] a_45670_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17043 a_34134_11906# a_18162_11500# a_34226_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17044 a_30210_9492# a_18546_9490# a_30118_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17045 a_11347_40214# a_11389_40443# a_11347_40541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17046 nmat.col_n[3] a_12250_4175# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17047 a_2250_31965# a_2163_31741# a_1846_31851# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17048 a_79085_40202# a_79181_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17049 VDD _1179_.X a_40402_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1705 VSS _1154_.X a_47591_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X17050 a_36234_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17051 a_22178_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17052 a_38546_18894# nmat.rowon_n[5] a_38150_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17053 VSS a_5331_28309# a_3351_27249# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17054 VSS a_24719_37429# a_14773_38306# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17055 VSS pmat.row_n[12] a_25494_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17056 a_22482_65206# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17057 a_10363_53153# a_6559_33767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17058 a_4259_24643# a_3305_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17059 VSS a_5423_67191# a_4421_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1706 VDD a_84028_9615# nmat.col_n[30] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X17060 a_45178_9898# a_18162_9492# a_45270_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17061 a_22578_17492# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17062 vcm a_18162_69222# a_39246_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17063 a_6914_57167# a_3866_57399# a_6611_57399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17064 a_49194_16926# pmat.row_n[8] a_49686_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17065 a_41699_52521# _1187_.A2 a_41481_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17066 a_4252_9839# a_4167_9615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17067 a_10677_44007# a_10985_44220# a_10651_44211# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X17068 a_20078_18934# a_18162_18528# a_20170_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17069 a_7072_26311# a_7186_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X1707 vcm a_18162_20536# a_24186_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17070 a_43262_67174# a_18546_67216# a_43170_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17071 a_50198_11906# pmat.row_n[3] a_50690_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17072 vcm a_18162_64202# a_40250_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17073 VSS ANTENNA__1196__A2.DIODE a_22280_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17074 a_6883_51335# a_4259_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X17075 a_36142_19938# pmat.row_n[11] a_36634_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17076 a_10305_19881# a_8305_20871# a_10233_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17077 a_35534_64202# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17078 a_40158_68178# pmat.row_n[12] a_40650_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17079 a_39246_57134# a_18546_57176# a_39154_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1708 a_47582_61190# pmat.rowon_n[5] a_47186_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17080 a_33130_21946# pmat.row_n[13] a_33622_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17081 a_22085_36374# a_21621_35515# a_22684_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X17082 a_33130_17930# a_18162_17524# a_33222_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17083 VDD pmat.rowon_n[3] a_43170_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17084 a_7521_47081# a_2215_47375# a_6747_46831# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X17085 VSS pmat.row_n[6] a_39550_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17086 VSS pmat.row_n[3] a_28506_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17087 a_20107_41046# a_19925_41046# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17088 a_25494_56170# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17089 VSS a_2007_42644# a_1895_43194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1709 VSS pmat.row_n[9] a_44570_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17090 a_6641_25731# a_4068_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17091 VSS a_2319_65564# a_2250_65693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17092 a_30210_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17093 a_32522_57174# pmat.rowon_n[1] a_32126_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17094 a_26594_16488# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17095 a_23090_13914# pmat.row_n[5] a_23582_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17096 a_2557_61885# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17097 a_23604_36391# a_22541_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17098 vcm a_18162_63198# a_44266_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17099 a_31371_29673# a_19405_28853# a_31299_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X171 VDD a_2319_59036# a_2250_59165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X1710 a_31518_67214# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17100 a_44174_67174# pmat.row_n[11] a_44666_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17101 a_2325_40821# a_2107_41225# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X17102 VSS comp.adc_comp_circuit_0.adc_comp_buffer_0.in comp.adc_comp_circuit_0.adc_comp_buffer_1.in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X17103 a_5329_54965# a_4075_68583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17104 a_29510_55166# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17105 VSS a_14773_38306# a_13837_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X17106 a_13139_54599# a_11202_55687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17107 VSS a_3956_59317# a_3894_59343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X17108 a_44570_22910# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17109 a_22377_49667# a_21371_50087# a_22281_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1711 VDD a_4863_13077# a_4379_13818# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X17110 a_21174_63158# a_18546_63200# a_21082_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17111 VSS a_8325_10901# a_8259_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17112 a_21574_67536# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17113 a_38242_18528# a_18546_18526# a_38150_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17114 a_51694_56492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17115 a_31122_24958# VDD a_31614_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17116 a_34226_62154# a_18546_62196# a_34134_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17117 a_21082_57134# a_18162_57174# a_21174_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17118 a_34626_66532# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17119 VDD a_6975_34538# a_6127_35076# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1712 a_10785_12015# a_2648_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17120 a_7477_31029# a_7259_31433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X17121 a_30210_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17122 VSS a_16083_50069# a_18429_51189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17123 VSS a_16745_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17124 VSS VDD a_48586_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17125 VDD a_38552_32521# a_38727_32447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17126 a_34134_56130# a_18162_56170# a_34226_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17127 VSS pmat.row_n[14] a_21478_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17128 a_17900_40743# a_16837_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17129 vcm a_18162_14512# a_39246_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1713 VDD a_30111_47911# a_35786_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X17130 VDD a_1781_9308# a_2193_11254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17131 VSS VDD a_46578_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17132 a_15107_44535# a_13985_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17133 a_8717_7485# a_8673_7093# a_8551_7497# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17134 VDD a_8385_51727# a_9995_52299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17135 a_50594_70226# pmat.rowon_n[14] a_50198_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17136 a_35138_62154# pmat.row_n[6] a_35630_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17137 a_29510_9858# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17138 a_12341_57141# a_6927_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17139 VDD a_6283_31591# a_28455_47381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1714 VSS a_23395_53135# a_27708_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X17140 a_37813_39867# a_36227_38771# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17141 VSS pmat.row_n[13] a_25494_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17142 a_20170_24552# a_18546_24550# a_20078_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17143 a_33281_49551# a_28915_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X17144 VSS a_30155_36893# a_30095_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X17145 a_40554_62194# pmat.rowon_n[6] a_40158_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17146 a_28602_57496# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17147 a_3211_77129# a_2695_76757# a_3116_77117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X17148 VDD a_5687_71829# a_5626_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X17149 a_6763_13103# a_5173_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1715 VDD a_6833_37281# a_6723_37405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X17150 VDD a_13091_18535# a_14839_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X17151 a_25590_51433# a_17139_30503# a_25287_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17152 VDD VSS a_32126_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17153 VDD a_11927_27399# a_17323_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17154 a_23486_72234# VDD a_23090_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17155 a_7063_57711# a_6835_51183# a_6700_57863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17156 vcm a_18162_20536# a_30210_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17157 a_33222_23548# a_18546_23546# a_33130_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17158 a_33839_46805# a_39647_48767# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17159 a_29206_13508# a_18546_13506# a_29114_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1716 a_48282_59142# a_18546_59184# a_48190_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17160 a_47211_50069# _1154_.A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17161 a_2215_17999# a_1591_18005# a_2107_18377# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17162 a_8703_6202# a_9459_5461# a_9417_5737# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17163 a_23815_28023# a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17164 VSS pmat.row_n[4] a_28506_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17165 a_37542_60186# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17166 a_40554_9858# nmat.rowon_n[14] a_40158_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17167 a_35171_50095# a_30663_50087# a_35077_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X17168 a_37542_19898# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17169 VDD a_41237_28585# a_41878_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1717 vcm a_18162_56170# a_45270_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17170 VDD a_46817_27221# nmat.col[27] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17171 a_22817_41317# a_22361_41479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17172 a_32522_10862# nmat.rowon_n[13] a_32126_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17173 a_7895_16694# a_7644_16341# a_7436_16519# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17174 VSS a_4319_15039# a_4253_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X17175 a_9552_67191# a_9545_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17176 a_38642_22512# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17177 a_42658_71552# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17178 VSS a_14261_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17179 VDD pmat.rowoff_n[12] a_42166_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1718 a_29933_52521# _1187_.A2 pmat.col_n[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X17180 a_6523_42479# a_6007_42479# a_6428_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17181 a_8612_63695# a_8175_63669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17182 VSS a_9337_15033# a_9271_15101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17183 nmat.rowon_n[13] a_14839_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17184 VSS a_4068_25615# a_5547_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17185 a_45270_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17186 a_42166_61150# a_18162_61190# a_42258_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17187 a_40256_42919# a_39193_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17188 a_2944_52789# a_2419_53351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17189 a_24214_29967# a_23043_28335# a_24214_30287# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X1719 a_23055_41781# a_10781_42364# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17190 a_25098_71190# a_18162_71230# a_25190_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17191 a_22522_50247# a_21371_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X17192 a_23815_50069# a_23971_50228# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X17193 VSS a_10569_64489# a_11713_64899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X17194 VSS pmat.row_n[10] a_27502_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17195 a_31518_58178# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17196 a_31518_16886# nmat.rowon_n[7] a_31122_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17197 VDD a_2411_33749# a_5132_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17198 VSS a_31701_37462# a_30765_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X17199 a_38083_32521# a_37637_32149# a_37987_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X172 a_2203_64073# a_1757_63701# a_2107_64073# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X1720 a_24833_34191# a_24667_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X17200 VDD a_36753_46805# a_36783_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17201 a_46674_70548# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17202 a_39154_14918# a_18162_14512# a_39246_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17203 VSS a_2163_74173# a_2124_74299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17204 a_19083_28879# a_14365_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17205 a_36663_34191# a_36486_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17206 a_1846_72107# a_2163_71997# a_2121_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17207 cgen.dlycontrol2_in[0] a_1591_37039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17208 a_16291_43805# a_12237_38772# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X17209 vcm a_18162_67214# a_32218_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1721 a_21478_59182# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17210 a_43262_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17211 a_5713_48463# a_4719_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17212 a_43566_69222# pmat.rowon_n[13] a_43170_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17213 a_46182_60146# a_18162_60186# a_46274_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17214 vcm a_18162_57174# a_28202_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17215 a_32218_55126# a_18546_55168# a_32126_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17216 vcm a_18162_17524# a_50290_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17217 a_29114_70186# a_18162_70226# a_29206_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17218 a_32618_59504# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17219 a_28506_14878# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1722 a_13354_2223# _1196_.B1 a_13185_2473# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X17220 VSS a_10985_42044# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17221 VDD a_10927_41245# a_10953_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X17222 a_19566_72556# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17223 a_20170_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17224 VDD a_37960_42693# a_37864_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X17225 a_41791_51727# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17226 VDD nmat.rowon_n[2] a_19074_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17227 VDD a_7160_33927# a_7067_34293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17228 VDD pmat.rowon_n[14] a_23090_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17229 VDD a_10995_76207# a_11397_76457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1723 VDD a_13160_31433# a_13335_31359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17230 VDD nmat.rowon_n[13] a_49194_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17231 VDD nmat.rowon_n[15] a_23090_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17232 cgen.dlycontrol3_in[1] a_1591_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17233 VDD a_32411_49559# a_28915_50959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X17234 a_19074_62154# a_18162_62194# a_19166_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17235 a_24861_29673# a_22307_27791# a_24861_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17236 a_23182_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17237 a_47582_68218# pmat.rowon_n[12] a_47186_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17238 VSS pmat.row_n[9] a_44570_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17239 VSS a_22527_27221# nmat.col[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1724 VDD a_13091_28327# a_26609_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X17240 a_33309_41479# a_33489_42043# a_34552_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X17241 VSS a_5266_17143# a_5271_17271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17242 a_6909_31061# a_6743_31061# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17243 VDD a_21970_48071# a_21923_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17244 a_42258_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17245 a_4255_69135# a_4396_69109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17246 VSS a_13432_62581# a_3923_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17247 a_45212_30761# a_30663_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17248 a_5445_62927# a_5462_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17249 a_21082_20942# a_18162_20536# a_21174_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1725 a_21478_17890# nmat.rowon_n[6] a_21082_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17250 a_83007_26703# ANTENNA__1395__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17251 vcm a_18162_18528# a_27198_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17252 a_21478_65206# pmat.rowon_n[9] a_21082_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17253 VSS pmat.row_n[0] a_47582_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17254 VDD pmat.rowon_n[5] a_44174_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17255 a_31214_16520# a_18546_16518# a_31122_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17256 VDD a_77245_40202# a_77058_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17257 VDD nmat.rowon_n[7] a_48190_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17258 a_14457_15823# a_14103_15936# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17259 a_6520_37039# a_6403_37252# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1726 VSS pmat.row_n[8] a_48586_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17260 VSS cgen.dlycontrol4_in[0] a_1945_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17261 a_26498_17890# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17262 VDD nmat.rowon_n[4] a_35138_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17263 VDD a_1923_69823# a_1643_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17264 VSS pmat.row_n[7] a_30514_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17265 a_7079_34837# a_6904_34863# a_7258_34863# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17266 VSS a_7865_16341# a_7799_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17267 a_8399_18115# a_7644_16341# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17268 a_36142_68178# a_18162_68218# a_36234_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17269 VDD a_16863_52815# pmat.rowon_n[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1727 a_2781_8585# a_1591_8213# a_2672_8585# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17270 VSS a_41297_27221# nmat.col[22] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17271 VDD nmat.sample a_18546_9490# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X17272 VSS a_4613_19087# a_5179_20175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17273 VSS a_10515_13967# a_16926_46261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17274 a_43261_48783# a_43315_48437# a_43273_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17275 a_7803_67655# a_5363_70543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X17276 a_49194_67174# a_18162_67214# a_49286_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17277 a_13443_43447# a_13837_43421# a_13503_43421# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X17278 vcm a_18162_72234# a_40250_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17279 a_35534_72234# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1728 a_45574_13874# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17280 comp.adc_comp_circuit_0.adc_comp_buffer_1.in comp.adc_inverter_1.in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17281 a_39246_65166# a_18546_65208# a_39154_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17282 a_44266_8488# a_18546_8486# a_44174_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17283 a_31122_58138# pmat.row_n[2] a_31614_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17284 a_39646_69544# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17285 VSS a_40105_47375# a_46763_44431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17286 VDD pmat.rowon_n[11] a_43170_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17287 a_31518_11866# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17288 VSS a_2648_29397# a_10388_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17289 a_39154_59142# a_18162_59182# a_39246_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1729 a_1857_5059# a_1761_7119# a_1775_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17290 nmat.col[7] a_10883_3303# a_14558_5263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17291 VSS a_79368_39738# a_79181_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17292 a_43262_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17293 VDD a_11067_27239# a_27249_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17294 a_13896_74953# a_12981_74581# a_13549_74549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X17295 VSS a_13837_37981# a_13529_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17296 a_31425_37218# a_30913_36603# a_31976_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X17297 a_9581_71855# a_9375_72007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X17298 a_26194_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17299 a_28506_55166# VSS a_28110_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X173 a_19074_56130# pmat.row_n[0] a_19566_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1730 VSS a_15144_36165# a_15107_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X17300 VDD a_12792_58633# a_12967_58559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17301 a_6914_9117# a_6548_8751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17302 a_43566_22910# nmat.rowon_n[1] a_43170_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17303 VDD a_37827_30793# a_37945_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X17304 a_41162_21946# pmat.row_n[13] a_41654_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17305 a_29711_47679# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17306 a_41162_17930# a_18162_17524# a_41254_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17307 a_7165_47081# a_4979_38127# a_6743_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X17308 a_11793_71311# a_9279_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17309 VDD a_12309_38659# a_39473_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1731 a_46274_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17310 VDD VSS a_30118_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17311 a_27411_46805# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17312 a_29510_63198# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17313 VSS a_28915_50959# a_46211_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17314 VSS pmat.row_n[8] a_20474_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17315 a_44174_12910# pmat.row_n[4] a_44666_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17316 a_47582_21906# nmat.rowon_n[2] a_47186_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17317 a_26659_34967# a_26767_34967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17318 a_34226_70186# a_18546_70228# a_34134_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17319 a_21082_65166# a_18162_65206# a_21174_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1732 a_36634_71552# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17320 a_27106_22950# pmat.row_n[14] a_27598_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17321 vcm a_18162_22544# a_48282_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17322 a_44320_32259# a_42791_32375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17323 a_3319_76751# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17324 VSS a_9827_53379# a_9639_53339# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17325 a_31614_20504# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17326 a_31214_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17327 VDD a_39472_48841# a_39647_48767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17328 a_4165_71017# a_2791_57703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17329 VSS a_8539_76181# a_6292_69831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1733 a_28506_23914# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17330 a_34134_64162# a_18162_64202# a_34226_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X17331 a_37542_13874# nmat.rowon_n[10] a_37146_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17332 a_23395_53135# a_38851_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17333 vcm a_18162_7484# a_23182_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17334 VDD a_25129_31751# a_25084_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X17335 a_3871_6031# a_3247_6037# a_3763_6409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17336 VDD pmat.rowoff_n[7] a_24094_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17337 a_21574_12472# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17338 VSS a_19928_37253# a_19817_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X17339 a_35242_30099# a_35520_30083# a_35476_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1734 a_11634_48285# a_11547_48061# a_11230_48171# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X17340 VSS a_43561_47893# a_43495_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17341 a_16890_36911# a_16713_36911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17342 a_40628_39429# a_39469_39141# a_40591_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17343 VSS a_4680_63669# a_3751_64757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X17344 a_35138_70186# pmat.row_n[14] a_35630_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17345 a_8453_46287# a_8079_46519# a_8381_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17346 a_43170_18934# pmat.row_n[10] a_43662_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17347 a_2672_33775# a_1591_33775# a_2325_34017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17348 a_32126_12910# a_18162_12504# a_32218_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17349 a_2369_23805# a_2325_23413# a_2203_23817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1735 a_32126_15922# pmat.row_n[7] a_32618_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17350 VSS pmat.row_n[13] a_32522_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17351 a_47839_30761# a_35244_32411# a_47767_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17352 a_9869_69921# a_9651_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X17353 result_out[8] a_1644_65845# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17354 VSS a_1674_68047# a_8031_76757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17355 a_36538_60186# pmat.rowon_n[4] a_36142_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17356 a_25590_11468# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17357 a_36538_19898# nmat.rowon_n[4] a_36142_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17358 a_1757_36501# a_1591_36501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17359 a_10677_37479# a_10985_37692# a_10651_37683# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1736 vcm a_18162_8488# a_27198_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17360 a_29206_21540# a_18546_21538# a_29114_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17361 a_47278_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17362 a_8267_49159# a_8907_48437# a_8853_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17363 a_20078_9898# pmat.row_n[1] a_20570_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17364 a_49590_9858# nmat.rowon_n[14] a_49194_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17365 a_83092_15055# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17366 a_34887_38007# a_33765_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17367 a_41254_68178# a_18546_68220# a_41162_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17368 a_33526_65206# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17369 VSS comp_latch a_7419_14379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1737 VSS pmat.row_n[13] a_32522_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17370 a_5510_9615# a_4865_8181# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17371 a_37238_58138# a_18546_58180# a_37146_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17372 VSS a_36419_28023# nmat.col_n[16] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17373 a_5553_73487# a_5497_73719# a_5363_73807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17374 a_19405_28853# a_7415_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17375 a_37987_32521# a_37471_32149# a_37892_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17376 a_47186_19938# pmat.row_n[11] a_47678_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17377 a_23663_39913# a_23700_39655# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X17378 VSS a_2319_59036# a_2250_59165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17379 VDD a_1925_26935# a_1738_26677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1738 a_1846_67755# a_2163_67645# a_2121_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X17380 a_23486_57174# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17381 a_20570_62516# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17382 a_7907_52031# a_7732_52105# a_8086_52093# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17383 a_22787_42325# a_10949_43124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17384 a_4523_21276# a_5179_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X17385 a_30514_58178# pmat.rowon_n[2] a_30118_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17386 a_44570_71230# pmat.rowon_n[15] a_44174_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17387 a_7407_17455# a_4976_16091# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17388 a_13769_24847# a_13367_24527# a_13683_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X17389 a_29114_63158# pmat.row_n[7] a_29606_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1739 a_29206_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17390 VDD a_24895_39605# a_24719_39605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X17391 a_33622_61512# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17392 a_27198_69182# a_18546_69224# a_27106_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17393 VSS a_1586_33927# a_3983_41941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17394 a_6803_77269# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17395 a_36142_8894# pmat.row_n[0] a_36634_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17396 a_24586_19500# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17397 a_12332_49917# a_5651_66975# a_11852_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17398 a_22684_40743# a_22269_40391# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X17399 VDD a_4866_52245# a_4259_73807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X174 a_27836_40743# a_27421_41814# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X1740 a_8439_69653# a_11391_69831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17400 VDD a_10515_61839# a_14011_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17401 a_12461_29423# a_11603_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17402 a_42562_8854# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17403 a_46674_8456# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17404 a_42562_23914# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17405 a_19675_51157# a_19831_51316# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X17406 a_39154_22950# a_18162_22544# a_39246_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17407 a_12242_51435# a_12559_51325# a_12517_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17408 a_36234_19532# a_18546_19530# a_36142_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17409 a_43262_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1741 a_36142_61150# a_18162_61190# a_36234_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17410 VSS a_31263_28309# a_30699_29397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.1275e+11p ps=3.87e+06u w=650000u l=150000u
X17411 vcm a_18162_65206# a_28202_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17412 a_28110_69182# pmat.row_n[13] a_28602_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17413 a_32218_63158# a_18546_63200# a_32126_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17414 a_32618_67536# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17415 a_49286_18528# a_18546_18526# a_49194_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17416 VSS pmat.row_n[10] a_35534_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17417 a_29864_39429# a_28705_39141# a_29768_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X17418 VSS pmat.row_n[0] a_28506_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17419 a_32126_57134# a_18162_57174# a_32218_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1742 a_12311_19783# a_9528_20407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17420 a_42795_28111# ANTENNA__1195__A1.DIODE nmat.col_n[22] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17421 VDD a_2191_27412# a_1895_27962# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X17422 a_46811_33927# a_30571_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X17423 VSS pmat.row_n[9] a_48586_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17424 cgen.dlycontrol4_in[1] a_1626_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17425 a_21124_36391# a_19965_36603# a_21028_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X17426 a_29124_37253# a_28061_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17427 VDD a_30819_40191# a_30679_40513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17428 a_1761_9839# a_1591_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17429 VSS _1184_.A2 a_38012_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1743 a_22178_56130# a_18546_56172# a_22086_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17430 a_13985_44581# a_12292_44869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17431 vcm a_18162_57174# a_36234_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17432 a_7631_15253# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17433 VSS pmat.row_n[14] a_32522_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17434 a_29206_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17435 a_45911_36815# a_43533_30761# a_45815_36815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17436 a_40250_55126# a_18546_55168# a_40158_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17437 a_40650_59504# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17438 VDD config_1_in[14] a_2235_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X17439 a_36538_14878# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1744 VSS a_4979_38127# a_6747_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5665e+12p ps=1.652e+07u w=650000u l=150000u M=4
X17440 vcm a_18162_56170# a_49286_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17441 a_29189_47349# a_28971_47753# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17442 a_19470_24918# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17443 a_25494_17890# nmat.rowon_n[6] a_25098_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17444 a_33949_39867# a_33007_38771# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X17445 a_5506_60751# a_4843_54826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17446 VSS a_10049_60663# a_11521_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17447 a_1643_61493# a_1846_61651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17448 a_49590_13874# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17449 a_46811_33927# a_44444_32233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 vcm a_18162_55166# a_49286_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17450 VSS a_30913_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17451 a_23090_55126# VDD a_23582_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17452 a_6621_16885# a_3305_17999# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17453 a_3894_59343# a_3175_59585# a_3331_59317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17454 a_31214_24552# a_18546_24550# a_31122_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17455 a_14486_47919# a_14528_48114# a_14486_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X17456 a_51598_62194# pmat.rowon_n[6] a_51202_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17457 VSS a_29217_41570# a_32035_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X17458 a_30210_66170# a_18546_66212# a_30118_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17459 a_27198_14512# a_18546_14510# a_27106_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1746 a_21621_35515# a_20848_36165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17460 VDD a_21867_34709# a_14773_37218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17461 a_26194_56130# a_18546_56172# a_26102_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17462 a_31976_36391# a_30913_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17463 a_25098_7890# VDD a_25590_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17464 a_14379_61519# a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17465 VDD pmat.rowon_n[2] a_30118_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17466 a_29510_16886# nmat.rowon_n[7] a_29114_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17467 VSS pmat.row_n[5] a_26498_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17468 a_23486_10862# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17469 VDD a_6823_58951# a_3938_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1747 a_19074_71190# a_18162_71230# a_19166_71190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17470 a_30514_11866# nmat.rowon_n[12] a_30118_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17471 a_5688_52423# a_5731_58951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17472 a_12107_62037# a_11842_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17473 a_48586_60186# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17474 VDD a_14773_38306# a_13837_37981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X17475 a_48586_19898# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17476 a_46667_46287# a_46582_46519# a_46449_46261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17477 a_50198_70186# a_18162_70226# a_50290_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17478 VSS pmat.row_n[10] a_38546_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17479 vcm a_18162_62194# a_31214_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1748 a_49194_59142# pmat.row_n[3] a_49686_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17480 a_31122_66170# pmat.row_n[10] a_31614_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17481 a_42562_64202# pmat.rowon_n[8] a_42166_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17482 a_36634_23516# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17483 a_5683_57711# a_5535_57993# a_5320_57863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17484 a_36234_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17485 a_27066_31599# a_24861_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17486 VDD nmat.rowon_n[2] a_40158_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17487 a_6093_74281# a_6051_74183# a_6009_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17488 a_43262_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17489 a_40158_62154# a_18162_62194# a_40250_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1749 VDD a_2100_44343# a_2051_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17490 a_49686_22512# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17491 a_39246_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17492 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17493 a_23090_72194# a_18162_72234# a_23182_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17494 a_28506_63198# pmat.rowon_n[7] a_28110_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17495 ctopp pmat.sw ctopp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u M=2
X17496 a_25190_17524# a_18546_17522# a_25098_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17497 a_39646_14480# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17498 a_37146_15922# a_18162_15516# a_37238_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17499 VDD pmat.rowoff_n[4] a_43170_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X175 a_1644_57141# a_1674_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1750 VSS pmat.row_n[5] a_22482_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17500 a_8031_26703# a_2683_22089# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17501 vcm a_18162_68218# a_30210_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17502 a_41254_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17503 a_25042_31055# a_24160_30199# a_24959_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X17504 VDD nmat.rowon_n[1] a_26102_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17505 a_2893_72765# a_2858_72531# a_2655_72373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17506 a_35390_47081# a_33957_48437# a_35306_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17507 a_31323_29967# a_31072_30083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X17508 VDD a_2683_22089# a_9385_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17509 VSS VDD a_20474_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1751 a_25494_16886# nmat.rowon_n[7] a_25098_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17510 a_1644_60949# a_1823_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17511 a_12242_51435# a_12520_51451# a_12476_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17512 a_3208_33597# a_3091_33402# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17513 a_19470_65206# pmat.rowon_n[9] a_19074_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17514 VSS pmat.row_n[5] a_50594_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17515 VSS a_79368_40202# a_79181_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17516 vcm a_18162_13508# a_26194_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17517 a_4341_7119# a_4254_7351# a_3551_6202# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17518 a_7118_32182# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17519 VSS pmat.row_n[15] a_33526_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1752 VDD a_2659_35015# a_2617_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17520 a_30210_11500# a_18546_11498# a_30118_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17521 a_6747_46831# a_4955_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X17522 VDD nmat.rowon_n[12] a_47186_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17523 a_4525_44655# a_2659_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X17524 VDD pmat.rowon_n[12] a_37146_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17525 a_4306_14735# a_3229_14741# a_4144_15113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17526 a_38546_68218# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17527 a_39219_52271# ANTENNA__1184__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17528 a_5227_15862# a_4976_16091# a_4768_16055# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17529 a_31214_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1753 a_48282_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17530 VSS a_5320_57863# a_3770_57399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17531 a_27198_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17532 VSS a_45370_48169# a_45428_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17533 a_18203_48981# a_18359_49140# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X17534 a_8360_7485# a_8243_7290# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X17535 vcm a_18162_59182# a_51294_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17536 a_3331_72373# a_3136_72515# a_3641_72765# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X17537 a_15048_41605# a_13985_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17538 a_34226_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17539 a_16911_52423# a_17183_52251# a_17141_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1754 a_11372_50461# a_10703_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17540 a_51598_16886# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17541 VSS a_5417_11445# a_5223_11079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17542 a_7808_61493# a_8193_61493# a_7937_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X17543 a_34949_52245# a_34705_51959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17544 VSS a_11057_35836# a_23883_34165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17545 a_40256_41831# a_39193_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17546 a_11327_39087# a_11339_39319# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17547 a_38242_60146# a_18546_60188# a_38150_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17548 a_38642_64524# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17549 vcm a_18162_19532# a_25190_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1755 a_83656_2767# ANTENNA__1196__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.955e+12p pd=1.791e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X17550 a_32126_20942# a_18162_20536# a_32218_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17551 a_16593_31849# a_1781_9308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17552 a_43170_69182# a_18162_69222# a_43262_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17553 VDD pmat.rowon_n[6] a_42166_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17554 VSS a_5654_9527# a_5721_8527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17555 VDD a_1923_61759# a_1643_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17556 a_24490_18894# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17557 VDD a_14287_70543# a_14839_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X17558 a_4719_69929# a_2419_69455# a_4801_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17559 a_11525_14433# a_11307_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1756 a_6541_15279# a_6375_15279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17560 VDD a_13605_71017# a_13158_71285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17561 a_29114_9898# pmat.row_n[1] a_29606_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17562 a_4253_15113# a_3063_14741# a_4144_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17563 VDD nmat.rowon_n[4] a_46182_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17564 a_4518_41935# a_3983_41941# a_4432_42313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17565 a_14749_47197# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X17566 a_2099_25236# a_2191_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17567 a_28202_71190# a_18546_71232# a_28110_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17568 a_50594_63198# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17569 a_39154_60146# pmat.row_n[4] a_39646_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1757 a_9063_24527# a_6829_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17570 vcm a_18162_7484# a_31214_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17571 a_47186_68178# a_18162_68218# a_47278_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17572 VSS pmat.row_n[13] a_40554_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17573 a_38907_48841# a_38391_48469# a_38812_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X17574 VDD pmat.rowon_n[7] a_28110_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17575 a_24186_9492# a_18546_9490# a_24094_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17576 VSS a_2375_63316# a_1895_63866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17577 VDD a_12309_36483# a_23420_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X17578 a_27794_28879# a_27355_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X17579 a_8084_71677# a_5779_71285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1758 a_12905_17973# a_12687_18377# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X17580 a_10839_11989# a_12967_12863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17581 VDD a_3622_29967# pmat.sw VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8e+11p ps=7.6e+06u w=1e+06u l=150000u M=5
X17582 a_5565_19605# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17583 a_12196_34215# a_11133_34427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17584 a_20570_70548# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17585 a_41254_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17586 VSS a_4025_54965# a_3970_55311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X17587 a_29114_71190# pmat.row_n[15] a_29606_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17588 a_24186_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17589 a_14738_59663# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X1759 a_23395_53135# a_26891_28327# a_44023_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X17590 VDD a_3866_57399# a_3431_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17591 VDD nmat.rowon_n[14] a_40158_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17592 a_41558_65206# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17593 pmat.rowon_n[14] a_14839_69135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17594 nmat.rowon_n[2] a_14747_7663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17595 a_41654_17492# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17596 a_41558_23914# pmat.rowoff_n[15] a_41162_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17597 a_3331_72373# a_3175_72641# a_3476_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X17598 a_30210_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17599 a_11501_10927# a_11207_11079# a_11417_10927# VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X176 VDD a_31879_34191# a_31985_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1760 vcm a_18162_67214# a_26194_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17600 VSS a_9405_66627# a_10249_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17601 a_21028_36391# a_19965_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17602 a_32969_29967# a_32865_30199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17603 a_12270_32509# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17604 a_26425_52521# _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17605 a_6343_18517# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17606 VSS a_2411_16101# a_10097_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17607 a_27198_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17608 a_4167_9615# a_2021_11043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X17609 a_6833_37281# a_6615_37039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1761 VSS pmat.row_n[7] a_47582_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17610 VSS a_6800_22869# a_6830_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17611 a_44570_56170# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17612 a_38546_21906# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17613 VDD a_11261_43421# a_10867_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17614 a_28543_27497# a_27763_27221# a_28325_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17615 a_45670_16488# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17616 a_35230_69182# a_18546_69224# a_35138_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17617 a_42166_13914# pmat.row_n[5] a_42658_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17618 a_27502_66210# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17619 a_14471_4943# ANTENNA__1190__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X1762 a_30210_65166# a_18546_65208# a_30118_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17620 VSS pmat.row_n[8] a_31518_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17621 a_25098_23954# pmat.row_n[15] a_25590_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17622 a_10205_51433# a_10245_51335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X17623 a_14830_3087# ANTENNA__1183__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X17624 a_25098_19938# a_18162_19532# a_25190_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17625 VDD a_7431_71829# a_7255_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X17626 a_83166_10703# ANTENNA__1190__A1.DIODE a_82788_10357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17627 a_7888_27907# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17628 VSS a_7099_74313# a_5403_67655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17629 VDD cgen.dlycontrol3_in[2] a_28975_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1763 a_8851_12533# a_8695_12801# a_8996_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X17630 a_32126_65166# a_18162_65206# a_32218_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17631 a_35534_14878# nmat.rowon_n[9] a_35138_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17632 a_12651_35823# a_12474_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17633 a_28110_55126# a_18162_55166# a_28202_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17634 a_24490_59182# pmat.rowon_n[3] a_24094_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17635 VSS pmat.row_n[0] a_21478_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17636 VSS config_2_in[13] a_2235_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17637 a_41703_27791# _1154_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17638 a_34611_36649# a_33489_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17639 a_48586_13874# nmat.rowon_n[10] a_48190_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1764 VDD a_33957_48437# a_33685_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X17640 VDD nmat.rowon_n[7] a_22086_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17641 vcm a_18162_65206# a_36234_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17642 a_36142_69182# pmat.row_n[13] a_36634_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17643 a_40250_63158# a_18546_63200# a_40158_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17644 a_28110_14918# pmat.row_n[6] a_28602_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17645 VDD a_35752_43781# a_35656_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X17646 a_40650_67536# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17647 a_29114_18934# a_18162_18528# a_29206_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17648 a_32618_12472# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17649 vcm a_18162_64202# a_49286_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1765 a_37542_69222# pmat.rowon_n[13] a_37146_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17650 a_49194_68178# pmat.row_n[12] a_49686_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17651 a_30118_13914# a_18162_13508# a_30210_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17652 a_24186_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17653 a_11469_35862# a_11297_36091# a_11255_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17654 a_50198_63158# pmat.row_n[7] a_50690_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17655 a_11021_43011# a_19689_42405# a_20811_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17656 VDD a_17619_43439# a_17725_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17657 VSS VDD a_25494_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17658 a_46752_46607# a_46027_44905# a_46449_46261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17659 a_32371_50247# a_32514_50141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1766 a_30610_69544# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17660 VSS pmat.row_n[14] a_40554_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17661 a_7072_52093# a_6835_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17662 a_4241_13653# a_4075_13653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17663 VSS a_32367_51946# pmat.col[12] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17664 a_26194_64162# a_18546_64204# a_26102_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17665 vcm a_18162_61190# a_23182_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17666 a_26594_68540# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17667 VDD pmat.rowon_n[10] a_30118_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17668 a_22830_27497# ANTENNA__1395__B1.DIODE a_22527_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17669 a_20173_30753# a_19955_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1767 vcm a_18162_17524# a_44266_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17670 VDD a_8307_23439# a_8417_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17671 a_30210_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17672 a_8481_10396# a_9195_7423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17673 a_4837_54447# a_4259_73807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17674 a_35630_7452# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17675 a_6953_5487# a_6574_5853# a_6881_5487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17676 VSS a_11339_39319# a_12764_40541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17677 vcm a_18162_70226# a_31214_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17678 a_35230_14512# a_18546_14510# a_35138_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17679 a_11533_64489# a_5651_66975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1768 a_26194_55126# a_18546_55168# a_26102_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17680 a_46765_51727# ANTENNA__1197__A.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17681 a_4871_17429# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X17682 a_20316_47607# a_18547_51565# a_20547_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17683 a_42562_72234# VDD a_42166_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17684 vcm a_18162_60186# a_27198_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17685 a_27106_64162# pmat.row_n[8] a_27598_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17686 a_2129_10383# a_1959_10383# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17687 VDD VDD a_45178_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17688 VSS VDD a_41558_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17689 a_31614_62516# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1769 a_26594_59504# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17690 a_48282_13508# a_18546_13506# a_48190_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17691 vcm a_18162_10496# a_45270_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17692 a_10111_30511# a_9595_30511# a_10016_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17693 a_40591_43447# a_39469_43493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17694 a_39246_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17695 a_32367_51946# a_32319_50345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17696 a_9375_72007# a_8919_71615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17697 a_51598_7850# VDD a_51202_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17698 a_3565_33597# a_3521_33205# a_3399_33609# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17699 a_7109_29423# a_7415_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X177 VDD a_30527_31573# a_30485_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1770 ANTENNA__1197__B.DIODE a_25695_28111# a_44389_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=8
X17700 a_9213_53903# a_8735_54207# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17701 VDD pmat.rowon_n[1] a_24094_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17702 a_39550_70226# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17703 vcm a_18162_22544# a_22178_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17704 a_22482_9858# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17705 VDD ANTENNA__1395__A1.DIODE a_41515_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17706 VSS a_13801_34427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17707 a_10499_67503# a_10226_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17708 a_40554_24918# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17709 a_25647_37607# a_21981_34191# a_25821_37483# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1771 a_10867_41271# a_11261_41245# a_10927_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X17710 VSS a_22541_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17711 VSS a_17478_46805# a_12079_9615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17712 a_27502_7850# VDD a_27106_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17713 a_37146_23954# a_18162_23548# a_37238_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17714 VDD cgen.dlycontrol1_in[1] a_25755_34343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X17715 a_22178_10496# a_18546_10494# a_22086_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17716 a_22056_27907# a_12061_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17717 VSS pmat.row_n[1] a_32522_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17718 VSS a_5731_58799# a_3866_57399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17719 a_24490_12870# pmat.rowoff_n[4] a_24094_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1772 VSS a_6369_39465# a_6619_41909# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17720 a_47278_19532# a_18546_19530# a_47186_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17721 VDD config_1_in[3] a_1591_13103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X17722 a_30118_58138# a_18162_58178# a_30210_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17723 vcm a_18162_21540# a_26194_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17724 a_44174_71190# a_18162_71230# a_44266_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17725 a_49590_62194# pmat.rowon_n[6] a_49194_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17726 a_43170_7890# a_18162_7484# a_43262_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17727 VSS pmat.row_n[10] a_46578_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17728 VSS a_10851_30485# a_10785_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17729 a_43566_15882# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1773 VDD a_11681_35823# a_11317_36924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X17730 a_13966_64783# a_12889_64789# a_13804_65161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17731 a_12075_24527# a_11897_21263# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.1e+11p pd=2.82e+06u as=0p ps=0u w=1e+06u l=150000u
X17732 a_24404_30287# a_24374_29941# a_24214_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17733 a_50594_16886# nmat.rowon_n[7] a_50198_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17734 a_5687_38279# a_5671_40097# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17735 a_4266_18038# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X17736 a_5131_16189# a_3688_17179# a_4768_16055# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X17737 VDD nmat.rowon_n[1] a_34134_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17738 a_10045_51727# a_9427_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17739 a_30118_17930# pmat.row_n[9] a_30610_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1774 a_11145_6575# a_9668_10651# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X17740 a_27198_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17741 a_19074_7890# a_18162_7484# a_19166_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17742 vcm a_18162_67214# a_51294_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17743 a_9135_23983# a_8291_23983# a_9217_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17744 vcm a_18162_57174# a_47278_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17745 VSS pmat.row_n[5] a_19470_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17746 a_6445_5487# a_5967_5461# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17747 a_12167_21263# a_5899_21807# a_11949_21237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17748 a_51294_55126# a_18546_55168# a_51202_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17749 a_21174_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1775 a_29036_41831# a_27877_42043# a_28999_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X17750 a_29206_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17751 a_51694_59504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17752 a_23486_18894# nmat.rowon_n[5] a_23090_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17753 a_7533_19087# a_7131_19407# a_7369_19407# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X17754 a_47582_14878# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17755 a_8568_26703# a_8031_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X17756 a_38642_72556# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17757 VDD pmat.rowon_n[14] a_42166_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17758 vcm a_18162_69222# a_24186_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17759 a_34134_16926# pmat.row_n[8] a_34626_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1776 VSS a_14719_37737# a_15651_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X17760 a_35230_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17761 vcm a_18162_9492# a_47278_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17762 a_11249_11177# a_11207_11079# a_11167_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17763 VDD pmat.rowon_n[4] a_38150_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17764 a_21082_19938# pmat.row_n[11] a_21574_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17765 a_18546_14510# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X17766 a_26957_38779# a_26276_39429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17767 a_17902_43439# a_17725_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17768 a_24186_57134# a_18546_57176# a_24094_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17769 a_10541_53387# a_9213_53903# a_10455_53387# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1777 a_19965_39867# a_19509_39638# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X17770 VSS a_33957_48437# a_33715_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17771 a_46705_38671# a_46427_39009# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17772 a_9463_8439# a_2648_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17773 a_8289_46607# a_3746_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17774 VSS a_7419_14379# a_7295_14441# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17775 VDD a_9375_72007# a_9333_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X17776 a_25190_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17777 VDD a_11693_70767# a_11893_71427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17778 VSS pmat.row_n[6] a_24490_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17779 a_45277_32687# a_44923_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1778 a_15844_52277# a_15657_52317# a_15757_52535# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X17780 a_13643_29415# a_34030_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17781 a_8197_76757# a_8031_76757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17782 a_33765_41317# a_33309_41479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X17783 a_3960_19465# a_2879_19093# a_3613_19061# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17784 a_3911_44431# a_2659_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X17785 a_27795_38007# a_28189_37981# a_12585_39355# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X17786 a_9963_54447# a_9213_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17787 VDD a_9460_10615# a_8111_11209# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17788 a_43267_47081# a_35186_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17789 a_6579_29199# a_4068_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1779 VSS pmat.row_n[9] a_38546_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17790 VDD pmat.rowon_n[15] a_28110_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17791 VSS pmat.row_n[11] a_36538_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17792 vcm a_18162_18528# a_46274_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17793 a_40554_65206# pmat.rowon_n[9] a_40158_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17794 VSS _1183_.A2 a_38996_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8675e+11p ps=3.79e+06u w=650000u l=150000u
X17795 a_50290_16520# a_18546_16518# a_50198_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17796 a_28202_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17797 VSS a_2787_55535# a_2882_54991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17798 a_40317_52271# ANTENNA__1187__B1.DIODE a_40099_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17799 VSS pmat.row_n[10] a_49590_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X178 vcm a_18162_22544# a_24186_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1780 a_14641_57167# a_14287_57280# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17800 a_4509_62037# a_4583_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X17801 a_2325_15797# a_2107_16201# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17802 VSS a_30543_40721# a_30489_40747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17803 VDD a_37709_52245# pmat.col[18] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17804 VDD nmat.rowon_n[14] a_49194_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17805 a_47678_23516# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17806 a_47278_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17807 VDD nmat.rowon_n[2] a_51202_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17808 a_26102_21946# a_18162_21540# a_26194_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17809 vcm a_18162_15516# a_20170_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1781 VDD a_6763_13103# a_7165_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X17810 a_23182_18528# a_18546_18526# a_23090_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17811 a_43566_56170# pmat.rowon_n[0] a_43170_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17812 a_37638_15484# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17813 VSS a_30913_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X17814 VDD nmat.rowon_n[10] a_41162_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17815 a_26498_66210# pmat.rowon_n[10] a_26102_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17816 a_4149_41941# a_3983_41941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17817 VDD a_2325_34017# a_2215_34141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17818 a_14486_46831# a_14379_46287# a_14486_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X17819 a_48190_15922# a_18162_15516# a_48282_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1782 VDD a_10569_64489# a_10957_64899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.197e+11p ps=1.41e+06u w=420000u l=150000u
X17820 a_14365_68743# a_13327_70741# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17821 a_20439_27247# a_10223_26703# a_20354_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X17822 vcm a_18162_14512# a_24186_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17823 a_45270_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17824 a_47582_55166# VSS a_47186_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17825 a_20499_31274# a_20591_31029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17826 a_29023_38571# a_23821_35279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17827 a_38150_11906# pmat.row_n[3] a_38642_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17828 VSS VDD a_31518_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17829 a_3514_57487# a_1591_56623# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X1783 a_21174_17524# a_18546_17522# a_21082_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17830 a_47186_9898# a_18162_9492# a_47278_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17831 a_11337_25071# a_9075_28023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17832 VDD pmat.rowon_n[13] a_35138_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17833 a_22111_36950# a_20605_40719# a_22039_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17834 VSS ANTENNA__1197__B.DIODE pmat.col[30] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17835 VSS a_40837_46261# a_45884_38377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17836 a_3173_25045# a_2648_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17837 a_35230_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17838 VDD pmat.rowon_n[12] a_48190_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17839 a_28110_63158# a_18162_63198# a_28202_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1784 a_31122_65166# pmat.row_n[9] a_31614_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17840 a_6277_18543# a_5087_18543# a_6168_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17841 a_12429_62607# a_12081_62723# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17842 a_10953_34951# a_11133_34427# a_12255_34473# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17843 a_36167_38825# a_36561_38780# a_36227_38771# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X17844 VDD a_13549_74549# a_13439_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17845 vcm a_18162_72234# a_49286_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17846 a_36634_65528# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17847 a_46182_22950# pmat.row_n[14] a_46674_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17848 VDD a_16163_43413# a_15921_38550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17849 a_50198_71190# pmat.row_n[15] a_50690_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1785 VDD nmat.rowon_n[6] a_38150_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17850 a_49286_60146# a_18546_60188# a_49194_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17851 a_36142_55126# a_18162_55166# a_36234_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17852 a_50690_20504# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17853 a_49686_64524# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17854 a_50290_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17855 VSS pmat.row_n[7] a_25494_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17856 a_22482_60186# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17857 a_22482_19898# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17858 result_out[11] a_1644_70197# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X17859 VSS a_30571_50959# a_45648_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1786 a_36234_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17860 a_39550_23914# pmat.rowoff_n[15] a_39154_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17861 a_36142_14918# pmat.row_n[6] a_36634_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17862 VSS pmat.row_n[12] a_36538_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17863 a_3026_28157# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17864 a_35534_18894# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17865 a_40650_12472# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17866 VSS a_26552_43781# a_26515_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X17867 a_26194_72194# a_18546_72236# a_26102_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17868 a_39646_56492# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17869 a_13801_38779# a_10927_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1787 a_16837_35515# a_16381_35286# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X17870 a_19074_24958# VDD a_19566_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17871 VSS a_11149_40188# a_11568_40541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17872 a_23582_22512# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17873 a_8031_13353# a_7165_13353# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17874 a_44266_22544# a_18546_22542# a_44174_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17875 a_6281_77537# a_6063_77295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X17876 VDD pmat.rowon_n[8] a_26102_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17877 a_51202_12910# a_18162_12504# a_51294_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17878 a_30561_52521# a_24867_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17879 a_30210_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1788 a_6554_43255# a_6619_41909# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=0p ps=0u w=650000u l=150000u
X17880 VSS pmat.row_n[13] a_51598_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17881 a_4535_38377# a_3325_36495# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17882 a_33684_32143# a_33205_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X17883 pmat.col_n[2] _1194_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17884 a_10691_28995# a_9395_27791# a_10609_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17885 a_7313_74005# a_2407_49289# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17886 a_27106_72194# VDD a_27598_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17887 a_38546_70226# pmat.rowon_n[14] a_38150_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17888 a_31614_70548# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17889 a_2163_65469# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1789 a_13259_41001# a_13653_40956# a_12235_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X17890 a_24094_14918# a_18162_14512# a_24186_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17891 a_48282_21540# a_18546_21538# a_48190_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17892 a_27598_60508# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17893 a_7900_54269# a_5211_57172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17894 a_23981_41835# a_10767_39087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17895 VSS a_1674_57711# a_9135_62613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17896 a_31122_60146# a_18162_60186# a_31214_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17897 a_28867_40871# a_28975_40871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17898 a_2107_26159# a_1757_26159# a_2012_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X17899 a_12061_26703# a_11713_26819# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X179 a_13977_23439# a_12463_22351# a_13559_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X1790 VDD a_33684_32143# a_34895_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X17900 a_10339_21263# a_10498_19631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17901 a_50198_18934# a_18162_18528# a_50290_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17902 a_19582_46983# a_19678_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17903 VSS a_24407_31375# a_40771_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17904 VSS a_14335_16519# a_14195_7351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17905 VDD a_1586_18231# a_2603_22357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X17906 a_42562_57174# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17907 a_9595_28879# a_4339_27804# a_9511_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X17908 VSS a_7521_19631# a_5351_19913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X17909 a_16552_46805# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X1791 VSS config_1_in[6] a_1591_2767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17910 VSS a_13091_52047# a_19759_48987# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17911 a_25494_67214# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17912 a_8013_25615# a_7665_25731# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X17913 a_32522_68218# pmat.rowon_n[12] a_32126_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17914 a_46274_69182# a_18546_69224# a_46182_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17915 vcm a_18162_66210# a_43262_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17916 a_2215_40847# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17917 a_43662_19500# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17918 VDD a_2847_43327# a_2834_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17919 VDD a_14471_27247# a_9963_28111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1792 a_12237_36596# a_12543_36950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17920 a_42562_9858# nmat.rowon_n[14] a_42166_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17921 VDD _1194_.B1 pmat.col_n[27] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X17922 VDD a_13275_48783# a_14461_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17923 VSS a_21032_44007# a_20995_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X17924 cgen.dlycontrol3_in[1] a_1591_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17925 a_4259_24643# a_3325_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17926 a_46578_14878# nmat.rowon_n[9] a_46182_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17927 a_25590_63520# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17928 VSS a_7295_14441# a_7085_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17929 VSS pmat.row_n[0] a_32522_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1793 a_49686_21508# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17930 a_10967_77532# a_10772_77563# a_11277_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X17931 a_5402_56079# a_5211_57172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17932 a_23935_52047# ANTENNA__1195__A1.DIODE pmat.col_n[4] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X17933 a_29606_18496# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17934 a_39497_29967# a_39127_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17935 VDD nmat.rowon_n[7] a_33130_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17936 VDD a_3351_27249# a_3123_27399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17937 vcm a_18162_65206# a_47278_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17938 a_47186_69182# pmat.row_n[13] a_47678_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17939 VDD a_18107_53034# pmat.rowoff_n[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1794 a_49286_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17940 a_51294_63158# a_18546_63200# a_51202_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17941 VDD nmat.rowon_n[4] a_20078_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17942 a_38205_32117# a_37987_32521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X17943 a_51694_67536# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17944 a_19470_58178# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17945 a_21082_68178# a_18162_68218# a_21174_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17946 a_13974_10749# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17947 a_51202_57134# a_18162_57174# a_51294_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17948 a_38996_50959# a_38770_50755# a_38627_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17949 VDD a_2199_13887# a_2740_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X1795 a_18953_43493# a_17996_41831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X17950 a_1644_71285# a_1591_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17951 a_35230_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17952 a_34134_67174# a_18162_67214# a_34226_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17953 VSS a_12934_35823# a_16147_36911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17954 a_2879_57487# a_4535_56623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17955 a_6428_42479# a_6311_42692# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17956 a_82787_13077# ANTENNA__1187__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17957 a_9313_22057# a_4703_24527# a_9217_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17958 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17959 a_51202_7890# a_18162_7484# a_51294_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1796 a_21082_57134# pmat.row_n[1] a_21574_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17960 a_24186_65166# a_18546_65208# a_24094_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17961 a_5138_65479# a_5267_65479# a_5275_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17962 VSS pmat.row_n[14] a_51598_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17963 a_5166_13353# a_5131_13255# a_4863_13077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17964 a_48282_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17965 a_24586_69544# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17966 vcm a_18162_17524# a_38242_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17967 a_42258_15516# a_18546_15514# a_42166_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17968 a_24094_59142# a_18162_59182# a_24186_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17969 VSS a_6979_51157# a_6925_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1797 a_42462_48071# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17970 a_4333_30511# a_4167_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17971 a_12152_66415# a_3923_68021# a_12049_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X17972 a_44570_17890# nmat.rowon_n[6] a_44174_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17973 cgen.dlycontrol2_in[4] a_2603_42479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17974 a_1757_63701# a_1591_63701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17975 a_40979_46287# a_40741_46565# a_40467_46261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17976 a_42166_55126# VDD a_42658_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17977 a_9339_28335# a_4339_27804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17978 VDD a_2046_30184# a_19439_32149# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X17979 a_25098_65166# pmat.row_n[9] a_25590_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1798 VSS a_42307_31756# a_25695_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.7375e+11p ps=3.75e+06u w=650000u l=150000u M=4
X17980 a_11848_48285# a_11634_48285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17981 a_23849_51727# _1192_.A2 pmat.col_n[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X17982 VSS pmat.row_n[0] a_21478_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17983 VDD nmat.rowon_n[15] a_25098_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17984 a_9871_53903# a_4128_64391# a_9953_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17985 a_46274_14512# a_18546_14510# a_46182_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17986 vcm a_18162_11500# a_43262_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17987 VDD a_12197_38306# a_11261_37981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X17988 a_45270_56130# a_18546_56172# a_45178_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17989 a_7865_16341# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1799 a_10055_31591# a_18947_49811# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X17990 a_37649_46607# a_33423_47695# a_37553_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17991 VSS pmat.row_n[5] a_45574_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17992 a_42562_10862# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17993 a_31518_8854# nmat.rowon_n[15] a_31122_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17994 VSS pmat.row_n[15] a_28506_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17995 VSS a_9655_6335# a_9589_6409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17996 a_25494_20902# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17997 a_3868_33609# a_2787_33237# a_3521_33205# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17998 vcm a_18162_23548# a_20170_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17999 a_28626_29423# a_15667_28111# a_28545_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.6575e+11p ps=1.81e+06u w=650000u l=150000u
X18 a_30210_59142# a_18546_59184# a_30118_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X180 VSS a_11116_18695# a_10975_18231# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1800 a_7343_16042# a_7387_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18000 a_20848_41605# a_19689_41317# a_20811_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18001 VDD a_36288_44527# a_36394_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18002 a_2121_67503# a_1643_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18003 a_12993_66415# a_12217_66389# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18004 a_32522_21906# nmat.rowon_n[2] a_32126_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18005 a_19166_16520# a_18546_16518# a_19074_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18006 a_5278_19631# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18007 a_28110_56130# pmat.row_n[0] a_28602_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18008 VSS a_38905_28853# a_37827_30793# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18009 a_37238_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1801 VSS a_3859_23699# a_2411_16101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X18010 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18011 VSS a_4037_69109# a_2944_69928# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18012 vcm a_18162_22544# a_33222_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18013 VSS a_10286_60405# a_10227_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18014 VDD a_9983_32385# a_9944_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18015 a_48190_23954# a_18162_23548# a_48282_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18016 a_4124_18231# a_3305_17999# a_4266_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X18017 a_4122_19087# a_3045_19093# a_3960_19465# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18018 a_5173_9839# a_3663_9269# a_5185_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18019 a_22482_13874# nmat.rowon_n[10] a_22086_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1802 a_10391_69653# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18020 a_42029_48169# a_42292_47893# a_41663_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X18021 a_7405_32441# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18022 a_47582_63198# pmat.rowon_n[7] a_47186_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18023 VSS a_19283_49783# a_24270_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18024 a_42166_72194# a_18162_72234# a_42258_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18025 VSS pmat.row_n[4] a_44570_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18026 a_23090_8894# a_18162_8488# a_23182_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18027 VSS pmat.row_n[11] a_44570_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18028 VDD a_12585_39355# a_27881_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X18029 a_18511_51433# a_12263_50959# a_18429_51189# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1803 a_31518_20902# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18030 VSS a_3583_11775# a_3517_11849# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X18031 a_34530_66210# pmat.rowon_n[10] a_34134_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18032 vcm a_18162_8488# a_36234_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18033 VSS pmat.row_n[14] a_27502_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18034 a_19074_58138# pmat.row_n[2] a_19566_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18035 a_5257_19087# a_5087_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18036 a_18546_55168# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X18037 a_47965_35951# a_38851_28327# a_47893_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18038 VSS a_2847_28095# a_2781_28169# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X18039 a_83827_26159# ANTENNA__1195__A1.DIODE nmat.col_n[29] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1804 a_9681_8527# a_9827_8181# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X18040 a_19470_11866# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18041 a_2882_67869# a_2163_67645# a_2319_67740# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18042 VSS a_4396_66933# a_4340_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18043 a_46274_8488# a_18546_8486# a_46182_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18044 VDD nmat.rowon_n[1] a_45178_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18045 _0467_ a_14371_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18046 vcm a_18162_58178# a_45270_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18047 VDD a_28915_50959# a_46487_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18048 a_21478_60186# pmat.rowon_n[4] a_21082_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18049 a_21478_19898# nmat.rowon_n[4] a_21082_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1805 a_34134_56130# pmat.row_n[0] a_34626_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18050 VDD a_39781_41245# a_39387_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18051 a_7665_25731# a_7779_22583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18052 a_3859_23699# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X18053 a_24747_29967# a_24214_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18054 a_32218_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18055 VDD nmat.rowon_n[9] a_35138_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18056 result_out[15] a_1644_76181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18057 a_36142_63158# a_18162_63198# a_36234_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18058 a_49686_72556# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18059 a_7429_52093# a_7385_51701# a_7263_52105# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1806 vcm a_18162_13508# a_22178_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18060 a_22178_58138# a_18546_58180# a_22086_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18061 VDD nmat.rowon_n[2] a_49194_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18062 a_20525_27247# a_10223_26703# a_20439_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X18063 a_21995_35101# a_12513_36924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18064 vcm a_18162_69222# a_35230_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18065 a_46274_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18066 a_43170_11906# a_18162_11500# a_43262_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18067 a_4036_67477# a_4421_67477# a_4165_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X18068 a_9177_6397# a_9133_6005# a_9011_6409# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18069 a_49194_62154# a_18162_62194# a_49286_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1807 a_25190_16520# a_18546_16518# a_25098_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18070 a_32126_19938# pmat.row_n[11] a_32618_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18071 a_1644_53877# a_1591_52815# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18072 a_20179_41046# a_14533_39631# a_20107_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X18073 VDD nmat.rowon_n[10] a_39154_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18074 a_36634_10464# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18075 VDD a_7109_29423# a_46857_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18076 a_7865_16341# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18077 a_19566_20504# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18078 VDD VDD a_26102_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18079 a_19166_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1808 a_43262_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18080 cgen.dlycontrol1_in[2] a_1591_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18081 a_13641_54965# a_13423_55369# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18082 a_4866_52245# a_2315_44124# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18083 a_51202_20942# a_18162_20536# a_51294_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18084 vcm a_18162_19532# a_44266_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18085 a_26194_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18086 a_77245_39738# a_77341_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18087 VSS pmat.row_n[11] a_47582_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18088 a_3160_29967# a_2217_29973# a_3052_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18089 VSS config_2_in[0] a_1591_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1809 VDD a_41731_49525# a_43971_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18090 a_51598_65206# pmat.rowon_n[9] a_51202_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18091 VDD a_13091_28327# a_34797_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18092 a_35730_47919# a_30111_47911# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X18093 vcm a_18162_7484# a_25190_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18094 a_24094_22950# a_18162_22544# a_24186_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18095 a_22449_49667# a_19584_52423# a_22377_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18096 a_1761_7119# a_1591_7119# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18097 VSS a_1586_33927# a_5823_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18098 VSS pmat.row_n[3] a_37542_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18099 VDD a_5415_71543# a_4409_74183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X181 a_42562_9858# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1810 a_39646_13476# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18100 VDD pmat.rowon_n[8] a_34134_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18101 a_21174_19532# a_18546_19530# a_21082_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18102 pmat.col_n[15] a_28915_50959# a_34497_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X18103 a_41558_57174# pmat.rowon_n[1] a_41162_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18104 VDD pmat.rowon_n[7] a_47186_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18105 a_35752_43781# a_34593_43493# a_35715_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18106 a_34226_18528# a_18546_18526# a_34134_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18107 VSS pmat.row_n[10] a_20474_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18108 a_12002_49667# a_11948_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18109 VDD a_4523_21276# a_13367_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.68e+11p ps=1.64e+06u w=420000u l=150000u
X1811 a_6334_65327# a_6292_65479# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X18110 a_6904_40303# a_5823_40303# a_6557_40545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X18111 a_5445_62927# a_5357_62779# a_5065_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18112 a_25393_43493# a_24937_43655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18113 a_36571_44527# a_36394_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18114 a_26957_37691# a_26501_37462# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18115 VSS pmat.row_n[9] a_33526_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18116 a_13273_10357# a_13055_10761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X18117 a_35630_60508# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18118 a_38546_55166# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18119 a_43262_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1812 a_4043_33535# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18120 vcm a_18162_57174# a_21174_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18121 a_8612_12559# a_8175_12533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18122 vcm a_18162_14512# a_35230_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18123 a_21478_14878# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18124 a_22086_9898# pmat.row_n[1] a_22578_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18125 vcm a_18162_56170# a_34226_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18126 a_40158_24958# VDD a_40650_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18127 a_7444_8751# a_7176_8751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18128 a_13345_40743# a_13653_40956# a_12235_39913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X18129 VDD pmat.rowon_n[13] a_46182_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1813 VDD nmat.rowon_n[12] a_43170_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18130 a_34530_13874# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18131 VDD a_5871_32362# a_5391_32900# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X18132 a_35656_43781# a_34593_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18133 a_32618_9460# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18134 a_1775_35113# a_1770_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18135 VSS a_5257_69679# a_5232_72373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18136 a_25590_71552# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18137 a_46274_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18138 a_43170_56130# a_18162_56170# a_43262_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18139 a_2433_52093# a_2398_51859# a_2195_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1814 a_25301_40229# a_23884_40517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18140 a_20752_44869# a_19689_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18141 a_29206_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18142 VSS config_1_in[14] a_2235_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18143 a_46578_66210# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18144 VSS pmat.row_n[8] a_50594_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18145 a_44174_23954# pmat.row_n[15] a_44666_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18146 a_35953_30333# a_2007_25597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18147 VDD a_8765_76725# a_8655_76751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18148 VSS a_13140_50247# a_13091_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18149 a_44174_19938# a_18162_19532# a_44266_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1815 a_28506_64202# pmat.rowon_n[8] a_28110_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18150 VSS a_4227_34293# a_4257_34319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18151 a_14458_5487# a_9411_2215# a_14372_5487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X18152 a_47678_65528# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18153 a_33489_36603# a_30155_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18154 a_51202_65166# a_18162_65206# a_51294_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18155 VSS a_19615_41959# a_19428_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18156 a_47186_55126# a_18162_55166# a_47278_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18157 VSS pmat.row_n[0] a_40554_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18158 a_2865_4943# a_2695_4943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18159 a_37542_24918# VSS a_37146_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1816 a_46578_9858# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18160 a_33526_60186# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18161 VDD a_6904_34863# a_7079_34837# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18162 VDD a_7865_16341# a_7895_16694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18163 a_33526_19898# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18164 VDD a_11067_16359# a_16679_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18165 VSS pmat.row_n[10] a_23486_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18166 a_37638_57496# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18167 VDD a_4339_27804# a_10765_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18168 VSS a_3727_66113# a_3688_65987# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18169 a_8695_12801# a_3571_13627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1817 a_11969_8751# a_9583_10121# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X18170 a_44570_8854# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18171 a_48682_8456# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18172 VDD a_10751_72917# a_10699_72943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18173 a_43072_50095# ANTENNA__1197__A.DIODE a_42769_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18174 VDD VSS a_41162_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18175 a_47186_14918# pmat.row_n[6] a_47678_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18176 VSS pmat.row_n[12] a_47582_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18177 a_21574_23516# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18178 a_21174_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18179 a_10513_24135# a_10239_20291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1818 a_37795_29111# a_37827_30793# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18180 a_42258_23548# a_18546_23546# a_42166_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18181 a_51694_12472# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18182 a_13328_55357# a_5682_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18183 VDD a_42683_32375# a_40903_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X18184 VSS a_5197_16121# a_5131_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18185 a_34626_22512# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18186 a_24186_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18187 VSS pmat.row_n[4] a_37542_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18188 a_27708_52271# ANTENNA__1190__A1.DIODE a_27405_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18189 a_38569_46831# a_1781_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1819 VDD a_33436_44527# a_33542_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18190 a_41558_10862# nmat.rowon_n[13] a_41162_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18191 VDD a_12431_69367# a_11487_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X18192 a_27995_30287# a_28715_28879# a_29282_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X18193 VDD nmat.rowon_n[6] a_27106_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18194 a_24586_14480# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18195 a_22086_15922# a_18162_15516# a_22178_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18196 a_25190_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18197 a_83196_3561# ANTENNA__1184__B1.DIODE nmat.col[19] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X18198 a_45270_64162# a_18546_64204# a_45178_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18199 vcm a_18162_61190# a_42258_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X182 a_42562_24918# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1820 a_2107_64073# a_1757_63701# a_2012_64061# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X18200 a_9441_20189# a_13427_18303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X18201 a_14264_72777# a_13183_72405# a_13917_72373# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18202 a_45670_68540# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18203 a_26609_51433# a_16311_28327# pmat.col[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18204 a_5785_48463# a_5411_48695# a_5713_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18205 a_35138_14918# a_18162_14512# a_35230_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18206 a_8455_7497# a_8105_7125# a_8360_7485# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18207 a_27877_42043# a_27421_41814# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18208 a_11230_48171# a_11508_48187# a_11464_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18209 VSS a_25681_28879# a_27355_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 vcm a_18162_12504# a_35230_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18210 a_19166_24552# a_18546_24550# a_19074_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18211 a_12237_36596# a_12543_36950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18212 a_28602_13476# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18213 a_25098_10902# pmat.row_n[2] a_25590_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18214 a_40554_58178# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18215 VDD nmat.rowon_n[12] a_32126_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18216 vcm a_18162_60186# a_46274_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18217 VDD pmat.rowon_n[12] a_22086_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18218 a_23486_68218# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18219 a_46182_64162# pmat.row_n[8] a_46674_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1822 a_10595_53361# a_10205_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X18220 VSS a_35068_46805# a_12263_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u M=2
X18221 a_19647_48052# a_19441_47491# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X18222 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18223 a_50690_62516# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18224 VDD a_11116_18695# a_10975_18231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18225 a_28079_37737# a_26957_37691# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18226 VDD a_2847_36799# a_2834_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18227 a_32957_30287# a_32865_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18228 a_27106_7890# VDD a_27598_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18229 a_26933_46831# a_26889_47073# a_26767_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1823 a_21478_12870# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18230 a_38193_29199# a_37827_30793# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X18231 a_36142_56130# pmat.row_n[0] a_36634_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18232 a_38150_70186# a_18162_70226# a_38242_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18233 vcm a_18162_62194# a_19166_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18234 a_26329_28111# a_15667_27239# nmat.col_n[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18235 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18236 a_19074_66170# pmat.row_n[10] a_19566_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18237 vcm a_18162_22544# a_41254_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18238 a_23182_60146# a_18546_60188# a_23090_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18239 a_33526_7850# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1824 VSS a_13327_70741# a_13575_68743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X18240 a_23582_64524# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18241 a_20078_61150# pmat.row_n[5] a_20570_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18242 vcm a_18162_12504# a_37238_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18243 a_4895_12559# a_4865_12533# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18244 a_41254_10496# a_18546_10494# a_41162_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18245 VDD a_38851_28327# a_45396_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X18246 a_34356_48783# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X18247 VSS pmat.row_n[14] a_35534_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18248 VDD nmat.rowon_n[4] a_31122_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18249 a_28061_36965# a_27605_37127# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X1825 VDD nmat.rowon_n[2] a_26102_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18250 a_24094_60146# pmat.row_n[4] a_24586_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18251 VDD a_21371_50087# a_24775_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18252 a_78802_40202# a_78898_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18253 a_32126_68178# a_18162_68218# a_32218_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18254 a_31122_8894# a_18162_8488# a_31214_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18255 a_22193_28995# a_21365_27247# a_22097_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18256 a_46274_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18257 VDD a_45019_38645# a_46949_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18258 a_21341_28585# a_8583_29199# a_21187_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18259 a_15101_29423# a_14829_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1826 a_27890_32143# a_27498_32117# a_26479_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X18260 VSS comp.adc_nor_latch_0.R comp_latch VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18261 nmat.col_n[31] ANTENNA__1197__B.DIODE a_82833_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18262 a_8355_11254# comp_latch a_7896_11079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18263 VSS pmat.row_n[5] a_38546_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18264 a_20474_7850# VDD a_20078_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18265 a_29772_40517# a_28613_40229# a_29735_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18266 a_40250_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18267 a_42562_18894# nmat.rowon_n[5] a_42166_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18268 a_25301_40229# a_23884_40517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18269 a_9685_74281# a_9655_74216# a_7099_74313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X1827 VSS a_1644_54421# result_out[1] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18270 a_3883_65845# a_3727_66113# a_4028_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18271 a_35138_59142# a_18162_59182# a_35230_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X18272 a_9183_72007# a_9279_71829# a_9581_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18273 a_49590_24918# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18274 a_19166_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18275 a_6823_58951# a_5081_53135# a_6990_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X18276 VSS a_16911_52423# a_14287_70543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18277 VDD a_13653_35516# a_13259_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18278 VSS a_23541_52245# pmat.col[4] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18279 vcm a_18162_59182# a_39246_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1828 VDD a_41731_49525# a_43191_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X18280 a_43262_57134# a_18546_57176# a_43170_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18281 VSS a_39193_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X18282 a_40158_58138# pmat.row_n[2] a_40650_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18283 a_7012_23145# a_3351_27249# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18284 a_37776_37479# a_36617_37691# a_37680_37479# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X18285 a_39550_16886# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18286 VSS a_7163_53333# a_7109_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18287 VDD config_1_in[4] a_1591_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18288 a_22541_36603# a_22085_36374# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18289 VSS pmat.row_n[6] a_43566_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1829 a_29206_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18290 a_40554_11866# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18291 a_37146_10902# a_18162_10496# a_37238_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18292 a_12217_66389# a_13973_66933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18293 a_10873_38517# a_30771_39425# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X18294 VDD VDD a_34134_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18295 a_26102_18934# pmat.row_n[10] a_26594_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18296 a_23486_21906# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18297 VSS VDD a_26498_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18298 a_5046_67655# a_3866_57399# a_5183_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X18299 a_35099_34191# a_34922_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X183 a_47582_7850# VDD a_47186_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1830 a_46578_62194# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18300 a_2882_56989# a_2124_56891# a_2319_56860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18301 a_30610_16488# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18302 a_20170_69182# a_18546_69224# a_20078_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18303 a_13606_18365# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18304 VDD pmat.rowon_n[15] a_47186_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18305 a_2905_14013# a_2526_13647# a_2833_14013# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X18306 a_22178_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18307 a_1644_70197# a_1591_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18308 a_8906_71311# a_7829_71317# a_8744_71689# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18309 a_19470_60186# pmat.rowon_n[4] a_19074_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1831 VDD a_11455_50237# a_11416_50363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18310 a_35230_7484# a_18546_7482# a_35138_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18311 a_19470_19898# nmat.rowon_n[4] a_19074_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18312 VDD a_29455_31293# a_28803_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X18313 a_20474_14878# nmat.rowon_n[9] a_20078_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18314 a_2861_76757# a_2695_76757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18315 a_1674_57711# a_1644_57685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18316 vcm a_18162_9492# a_40250_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18317 a_8937_15823# a_8767_15823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18318 VSS pmat.row_n[7] a_29510_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18319 a_38546_63198# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1832 VSS a_1761_4399# a_1775_5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X18320 a_33526_13874# nmat.rowon_n[10] a_33130_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18321 a_12124_47197# a_11910_47197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X18322 vcm a_18162_65206# a_21174_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18323 VSS a_14195_7351# a_14195_7119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18324 a_21082_69182# pmat.row_n[13] a_21574_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18325 VSS ANTENNA__1197__A.DIODE pmat.col_n[0] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X18326 vcm a_18162_64202# a_34226_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18327 a_34134_68178# pmat.row_n[12] a_34626_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18328 a_45574_66210# pmat.rowon_n[10] a_45178_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18329 VSS ANTENNA__1184__B1.DIODE a_12066_3087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1833 a_4831_34561# a_1586_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18330 a_26194_9492# a_18546_9490# a_26102_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18331 VDD pmat.rowoff_n[15] a_43170_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18332 a_15722_31599# a_1858_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18333 a_13091_7655# a_16552_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18334 a_13620_10761# a_12705_10389# a_13273_10357# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X18335 a_43170_64162# a_18162_64202# a_43262_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18336 VSS a_9441_20189# a_10287_24759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18337 a_5621_48783# a_4719_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18338 VSS a_28915_50959# a_47591_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18339 a_8481_18115# a_7809_17705# a_8399_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1834 VSS pmat.row_n[4] a_50594_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18340 VSS VDD a_50594_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18341 VDD nmat.rowon_n[14] a_42166_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18342 a_49590_65206# pmat.rowon_n[9] a_49194_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18343 a_37519_46983# a_33423_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18344 VDD nmat.rowon_n[9] a_46182_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18345 VDD a_3571_13627# a_9319_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18346 a_44266_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18347 a_14372_58799# a_10239_14183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18348 a_31596_34191# a_31419_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18349 a_45396_31849# a_45019_38645# a_45589_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1835 a_18973_29199# a_8583_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18350 a_47186_63158# a_18162_63198# a_47278_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18351 a_39550_57174# pmat.rowon_n[1] a_39154_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18352 a_17203_48579# a_16800_47213# a_17131_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18353 a_20170_14512# a_18546_14510# a_20078_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18354 a_20474_71230# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18355 a_20787_30199# a_20895_30199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18356 VSS pmat.row_n[8] a_19470_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18357 a_1644_56053# a_1591_56623# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18358 VDD ANTENNA__1196__A2.DIODE a_83839_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18359 vcm a_18162_15516# a_29206_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1836 VSS pmat.row_n[11] a_50594_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18360 a_33222_13508# a_18546_13506# a_33130_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18361 vcm a_18162_10496# a_30210_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18362 a_47678_10464# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18363 VSS a_45805_32661# a_45119_32661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18364 a_24186_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18365 VDD a_2046_30184# a_5823_34863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18366 a_41558_60186# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18367 a_41558_19898# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18368 VDD a_8197_20871# a_10333_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X18369 a_2325_17973# a_2107_18377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X1837 a_29510_72234# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18370 a_24490_70226# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18371 a_7894_51727# a_6817_51733# a_7732_52105# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18372 a_40158_9898# a_18162_9492# a_40250_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18373 a_2595_13621# a_2400_13763# a_2905_14013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18374 a_22086_23954# a_18162_23548# a_22178_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18375 a_45270_72194# a_18546_72236# a_45178_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18376 a_33719_44527# a_33542_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18377 a_10513_24643# a_9441_20189# a_10422_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18378 a_38150_63158# pmat.row_n[7] a_38642_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18379 a_35138_22950# a_18162_22544# a_35230_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1838 VDD a_1586_18231# a_4075_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18380 VDD pmat.rowon_n[8] a_45178_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18381 a_42658_61512# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18382 a_32218_19532# a_18546_19530# a_32126_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18383 a_2325_42997# a_2107_43401# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18384 a_26194_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18385 a_27502_61190# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18386 VSS _1154_.A a_40415_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18387 VSS pmat.row_n[10] a_31518_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18388 VSS a_28915_50959# a_47724_47081# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18389 VDD a_17012_47349# a_14379_6567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1839 VSS pmat.row_n[14] a_33526_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18390 a_2781_28169# a_1591_27797# a_2672_28169# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18391 a_22541_39867# a_21124_39655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18392 VDD pmat.rowon_n[0] a_35138_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18393 VSS a_3207_65845# a_1823_68565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18394 VDD a_10515_15055# a_14646_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18395 a_46182_72194# VDD a_46674_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18396 a_14174_51859# a_14452_51843# a_14408_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18397 a_47035_37289# a_43776_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18398 VDD a_3325_20175# a_8338_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18399 a_50690_70548# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X184 a_39154_23954# a_18162_23548# a_39246_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1840 a_3325_20175# a_2847_20479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18400 a_12491_32509# a_7939_31591# a_12128_32375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18401 a_46674_60508# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18402 vcm a_18162_57174# a_32218_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18403 a_7841_52105# a_6651_51733# a_7732_52105# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18404 a_11759_10615# comp_latch VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18405 a_4144_15113# a_3229_14741# a_3797_14709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X18406 vcm a_18162_70226# a_19166_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18407 a_32522_14878# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18408 VDD VSS a_39154_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18409 a_13620_10761# a_12539_10389# a_13273_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1841 VDD a_34816_34191# a_34922_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18410 a_23582_72556# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18411 vcm a_18162_20536# a_37238_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18412 a_38727_32447# a_2007_25597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18413 a_19566_62516# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18414 a_20170_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18415 a_28116_39655# a_26957_39867# a_28020_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X18416 VDD pmat.rowon_n[4] a_23090_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18417 a_44570_67214# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18418 a_20811_38007# a_19689_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18419 VDD a_25839_49783# a_25743_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1842 vcm a_18162_71230# a_47278_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18420 VDD VDD a_47186_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18421 VSS VDD a_43566_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18422 a_39550_10862# nmat.rowon_n[13] a_39154_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18423 a_2499_13077# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18424 a_36538_9858# nmat.rowon_n[14] a_36142_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18425 a_40954_29423# a_38905_28853# a_40785_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18426 a_4266_27830# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X18427 VSS a_30155_42583# a_12116_40871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X18428 a_23083_47753# a_22567_47381# a_22988_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18429 VDD a_3521_33205# a_3411_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1843 VDD pmat.rowon_n[11] a_37146_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18430 VSS pmat.row_n[11] a_21478_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18431 VDD a_4991_69831# a_11559_68619# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18432 a_24490_9858# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18433 ANTENNA__1395__A1.DIODE a_47591_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X18434 vcm a_18162_18528# a_31214_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18435 VSS pmat.row_n[0] a_51598_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18436 a_48682_18496# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18437 a_48586_24918# VSS a_48190_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18438 a_45178_15922# pmat.row_n[7] a_45670_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18439 a_29510_7850# VDD a_29114_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1844 a_31214_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18440 a_8452_65149# a_5307_67655# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18441 VSS a_13427_18303# a_13361_18377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X18442 VSS pmat.row_n[10] a_34530_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18443 a_42709_27791# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18444 a_22493_31353# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18445 VSS pmat.row_n[1] a_34530_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18446 a_32618_23516# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18447 a_22111_37277# a_21857_36950# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18448 VSS a_6612_15797# a_1586_8439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18449 VDD a_2375_16532# a_1895_15994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1845 a_7355_37013# a_7180_37039# a_7534_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18450 a_32218_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18451 a_5271_17271# a_5266_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18452 a_83092_27023# ANTENNA__1395__A1.DIODE a_82789_26677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18453 VSS a_14287_69455# a_14839_68047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18454 a_3303_33609# a_2787_33237# a_3208_33597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18455 a_38546_16886# nmat.rowon_n[7] a_38150_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18456 VSS a_39079_40947# a_39321_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X18457 a_10245_51335# a_9995_52299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X18458 a_45178_7890# a_18162_7484# a_45270_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18459 a_22578_15484# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1846 a_18235_39095# a_17113_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X18460 VDD nmat.rowon_n[5] a_25098_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18461 vcm a_18162_67214# a_39246_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18462 a_43262_65166# a_18546_65208# a_43170_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18463 vcm a_18162_62194# a_40250_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18464 a_43662_69544# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18465 a_40158_66170# pmat.row_n[10] a_40650_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18466 a_39246_55126# a_18546_55168# a_39154_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18467 a_39646_59504# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18468 a_12003_52815# a_11752_52931# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18469 a_33130_15922# a_18162_15516# a_33222_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1847 a_27198_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18470 a_2610_21807# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18471 a_43591_48246# a_43267_47081# a_43132_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18472 a_13144_65149# a_5462_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18473 a_14943_26703# a_14725_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X18474 a_26102_69182# a_18162_69222# a_26194_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18475 VDD a_5232_72373# a_3956_72373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18476 VSS pmat.row_n[1] a_28506_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18477 pmat.rowon_n[7] a_21647_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X18478 a_30210_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18479 a_32522_55166# VSS a_32126_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1848 VDD a_10873_39605# a_10817_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18480 VSS a_15543_31573# a_15477_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18481 VDD a_34277_38550# a_33341_38780# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X18482 a_2319_69916# a_2163_69821# a_2464_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X18483 a_23090_11906# pmat.row_n[3] a_23582_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18484 VSS a_6559_8527# a_7648_9117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=640000u l=150000u
X18485 VDD a_12047_14165# a_12034_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18486 a_4597_44655# a_2315_44124# a_4525_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18487 a_17322_49667# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18488 VDD pmat.rowon_n[13] a_20078_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18489 pmat.rowon_n[13] a_14839_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1849 a_2405_19087# a_2228_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18490 a_44174_65166# pmat.row_n[9] a_44666_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18491 vcm a_18162_9492# a_49286_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18492 VDD a_5197_16121# a_5227_15862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18493 a_29206_66170# a_18546_66212# a_29114_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18494 a_8563_7119# a_7939_7125# a_8455_7497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18495 a_20170_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18496 VDD nmat.rowon_n[4] a_29114_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18497 VSS a_18795_28882# a_19083_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18498 a_33299_32143# a_32771_31599# a_33205_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X18499 VDD pmat.rowon_n[12] a_33130_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X185 a_24186_10496# a_18546_10494# a_24094_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1850 vcm a_18162_58178# a_51294_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18500 a_11116_18695# a_9441_20189# a_11258_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X18501 a_12513_39100# a_13555_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18502 a_13985_35877# a_13319_35507# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18503 a_11023_76359# a_10699_75119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18504 VDD a_2672_16201# a_2847_16127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18505 VSS a_19268_34191# a_19374_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18506 a_6732_44111# a_4399_51157# a_6641_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X18507 a_35178_32509# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18508 a_44570_20902# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18509 a_10589_22351# a_10209_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1851 a_47678_63520# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18510 VSS a_29772_40517# a_29735_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18511 a_82787_14709# ANTENNA__1183__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18512 vcm a_18162_72234# a_34226_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18513 a_21574_65528# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18514 a_47186_56130# pmat.row_n[0] a_47678_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18515 a_3054_54223# a_2791_57703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18516 a_38242_16520# a_18546_16518# a_38150_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18517 a_4707_32156# a_16635_31573# a_16593_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18518 VSS pmat.row_n[15] a_42562_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18519 a_31122_22950# pmat.row_n[14] a_31614_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1852 a_6579_21583# a_3351_27249# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18520 VSS a_5038_28853# a_4679_28853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18521 a_34226_60146# a_18546_60188# a_34134_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18522 a_21082_55126# a_18162_55166# a_21174_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18523 a_34626_64524# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18524 vcm a_18162_12504# a_48282_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18525 a_4123_16042# a_4215_15797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18526 a_2012_23805# a_1895_23610# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18527 VDD a_2315_44124# a_4257_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18528 a_11977_66665# a_11883_62063# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18529 a_30210_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1853 VSS pmat.row_n[6] a_23486_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18530 VDD a_2935_38279# a_4351_39872# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18531 a_24490_23914# pmat.rowoff_n[15] a_24094_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18532 a_21082_14918# pmat.row_n[6] a_21574_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18533 VSS pmat.row_n[12] a_21478_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18534 a_22871_29967# a_22459_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18535 a_9090_56079# a_8013_56085# a_8928_56457# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18536 a_5805_49007# a_5639_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18537 a_24586_56492# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18538 VSS a_2389_45859# a_4837_45519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X18539 VSS pmat.row_n[14] a_46578_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1854 a_20474_18894# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18540 a_3026_8573# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X18541 a_11507_39087# a_11327_39087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18542 a_12061_9001# a_9583_10121# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X18543 VSS a_36571_44527# a_36677_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18544 a_35138_60146# pmat.row_n[4] a_35630_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18545 a_44266_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18546 a_8587_23555# a_7779_22583# a_8491_23555# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18547 a_34942_51701# a_26891_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18548 VSS a_11427_73180# a_11358_73309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18549 a_4503_6335# a_4328_6409# a_4682_6397# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1855 VDD a_14641_57711# a_14839_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X18550 a_13555_37782# a_13597_37571# a_13555_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18551 a_30913_38053# a_29220_37253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18552 VSS pmat.row_n[6] a_36538_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18553 VSS a_8439_69653# a_7730_69109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X18554 a_40554_60186# pmat.rowon_n[4] a_40158_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18555 a_40554_19898# nmat.rowon_n[4] a_40158_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18556 VSS VDD a_19470_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18557 a_28602_55488# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18558 a_1643_71829# a_1846_72107# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18559 VDD a_2935_38279# a_4399_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1856 a_5043_37191# a_2659_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X18560 vcm a_18162_23548# a_29206_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18561 VSS a_8305_20871# a_8399_18115# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18562 a_23486_70226# pmat.rowon_n[14] a_23090_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18563 a_3727_66113# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18564 VSS pmat.row_n[5] a_49590_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18565 VSS a_31675_47695# a_44665_45519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18566 a_33222_21540# a_18546_21538# a_33130_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18567 a_4705_39759# a_4351_39872# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18568 a_51294_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18569 VDD a_4339_27804# a_11867_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1857 VDD pmat.rowon_n[5] a_51202_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18570 VSS a_4339_27804# a_11713_26819# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18571 a_37238_71190# a_18546_71232# a_37146_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18572 a_7044_62607# a_5081_53135# a_6583_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18573 VSS a_4979_38127# a_5455_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18574 a_29206_11500# a_18546_11498# a_29114_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18575 a_11881_16911# a_11711_16911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18576 a_10284_32143# a_10070_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18577 VDD VSS a_37146_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18578 a_49194_9898# a_18162_9492# a_49286_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18579 a_55418_40254# comp.adc_nor_latch_0.R comp_latch VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1858 a_12212_22467# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18580 a_41254_58138# a_18546_58180# a_41162_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18581 VSS pmat.row_n[2] a_28506_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18582 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18583 a_4809_63695# a_4583_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18584 a_10319_50959# a_9427_50095# a_9457_51163# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18585 a_11969_8751# a_11051_8903# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18586 a_51202_19938# pmat.row_n[11] a_51694_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18587 a_19689_39141# a_18272_39429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18588 VSS a_12263_50959# a_17049_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18589 a_26498_61190# pmat.rowon_n[5] a_26102_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1859 VDD a_2944_65576# a_2882_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X18590 VDD _1179_.X a_45554_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X18591 a_7415_29397# a_10097_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X18592 a_6634_26133# a_4068_25615# a_6657_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18593 a_48190_10902# a_18162_10496# a_48282_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18594 a_38150_71190# pmat.row_n[15] a_38642_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18595 VSS a_9375_72007# a_9225_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18596 a_38642_20504# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18597 VDD VDD a_45178_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18598 a_12967_58559# a_1957_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18599 a_12277_51183# a_12242_51435# a_11807_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X186 a_31518_69222# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1860 a_37542_22910# nmat.rowon_n[1] a_37146_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18600 a_38242_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18601 a_31214_69182# a_18546_69224# a_31122_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18602 a_45270_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18603 a_27198_59142# a_18546_59184# a_27106_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18604 VSS a_9368_9991# a_8472_11739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18605 a_28202_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18606 VSS pmat.row_n[8] a_27502_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18607 VSS a_40969_30287# a_41795_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X18608 a_6681_62927# a_4025_54965# a_6583_62607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X18609 a_31518_14878# nmat.rowon_n[9] a_31122_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1861 a_32514_50141# a_25879_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18610 VSS a_5558_9527# a_6017_6575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18611 conversion_finished_out a_1644_77813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18612 VDD a_12235_39913# a_13345_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X18613 a_8789_60431# a_8841_60405# a_6175_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18614 a_39154_12910# a_18162_12504# a_39246_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18615 a_40250_19532# a_18546_19530# a_40158_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18616 a_33719_34191# a_33542_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18617 VSS a_14113_36604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X18618 a_25667_35253# a_11317_36924# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18619 vcm a_18162_65206# a_32218_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1862 a_39473_41605# a_31793_41570# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X18620 VSS pmat.row_n[13] a_39550_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18621 a_32126_69182# pmat.row_n[13] a_32618_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18622 vcm a_18162_55166# a_28202_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18623 a_43566_67214# pmat.rowon_n[11] a_43170_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18624 a_28110_59142# pmat.row_n[3] a_28602_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18625 vcm a_18162_15516# a_50290_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18626 a_39647_48767# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18627 a_22715_32521# a_22199_32149# a_22620_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X18628 VSS a_39193_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X18629 a_1849_45205# a_1683_45205# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1863 a_33526_17890# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18630 a_22043_35041# a_12345_36924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18631 a_37129_36130# a_36617_36603# a_37680_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X18632 a_19566_70548# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18633 a_20170_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18634 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18635 a_19074_60146# a_18162_60186# a_19166_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18636 VDD a_39939_29967# a_40509_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18637 a_33222_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18638 vcm a_18162_17524# a_23182_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18639 VSS a_22537_36911# a_40399_36911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1864 a_39387_40183# a_39781_40157# a_12309_38659# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X18640 a_35476_29967# a_35039_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18641 a_29206_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18642 a_13167_42359# a_13561_42333# a_13227_42333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X18643 VDD a_1591_61519# a_4135_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18644 a_38150_18934# a_18162_18528# a_38242_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18645 a_18487_50069# a_18823_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X18646 VSS a_9668_10651# a_10789_6575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18647 VSS a_19487_49159# a_18359_49140# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18648 a_7929_24233# a_6173_22895# a_7847_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18649 VSS a_13768_22325# a_14642_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1865 VSS a_12531_42583# a_12344_42325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18650 a_37542_58178# pmat.rowon_n[2] a_37146_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18651 pmat.col_n[30] a_46934_53135# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18652 a_2012_50095# a_1895_50308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18653 a_30913_36603# a_29404_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18654 pmat.col_n[12] a_31535_49525# a_31307_49871# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18655 vcm a_18162_16520# a_27198_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18656 a_48282_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18657 a_45178_66170# a_18162_66210# a_45270_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18658 nmat.rowoff_n[10] a_9963_13967# a_14011_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X18659 a_31214_14512# a_18546_14510# a_31122_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1866 VSS a_43659_28853# a_44463_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X18660 a_30210_56130# a_18546_56172# a_30118_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18661 a_26498_15882# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18662 VSS pmat.row_n[5] a_30514_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18663 VSS a_1923_31743# a_3565_33597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18664 VSS a_12604_47080# a_12542_47197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18665 VSS a_9731_8439# a_9681_8527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18666 VDD nmat.sample a_18546_7482# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X18667 a_44570_9858# nmat.rowon_n[14] a_44174_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18668 a_38546_8854# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18669 a_46522_34293# a_32405_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X1867 a_24186_71190# a_18546_71232# a_24094_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18670 a_22178_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18671 VSS a_9583_10121# a_11813_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18672 a_6997_25731# a_3305_27791# a_6924_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X18673 a_12981_8213# a_12815_8213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18674 vcm a_18162_70226# a_40250_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18675 a_35534_70226# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18676 a_6833_17027# a_3305_17999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18677 a_39246_63158# a_18546_63200# a_39154_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18678 a_45866_38279# a_45625_36495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X18679 a_9831_74183# a_10697_75218# a_10693_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1868 a_83677_3855# _1194_.A2 nmat.col[28] VDD sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u M=4
X18680 a_40650_23516# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18681 a_39646_67536# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18682 a_40250_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18683 a_6168_18543# a_5253_18543# a_5821_18785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18684 a_33130_23954# a_18162_23548# a_33222_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18685 VDD pmat.rowon_n[9] a_43170_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18686 a_49194_24958# VDD a_49686_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18687 VSS a_5871_32362# a_5391_32900# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18688 VSS a_1643_56597# a_1591_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18689 a_22620_32509# a_6007_33767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X1869 _1196_.B1 a_44533_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u M=16
X18690 a_25280_46831# a_13275_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18691 a_39154_57134# a_18162_57174# a_39246_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18692 a_2250_54991# a_2124_55107# a_1846_55123# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18693 pmat.rowon_n[2] a_12447_16143# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X18694 VDD a_24643_51959# pmat.col_n[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X18695 a_10967_77532# a_10811_77437# a_11112_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18696 a_25494_62194# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18697 a_6451_67655# a_13102_71311# a_13966_71631# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X18698 a_43262_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18699 VSS a_4976_16091# a_6621_16885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X187 VDD a_6559_8527# a_7648_9117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.499e+11p ps=2.35e+06u w=840000u l=150000u
X1870 VSS nmat.sample a_18546_17522# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X18700 a_37743_27497# a_24591_28327# a_37525_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18701 a_32522_63198# pmat.rowon_n[7] a_32126_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18702 a_27616_52047# ANTENNA__1190__A1.DIODE a_27313_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18703 a_11852_49783# a_12002_49917# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18704 a_2715_51969# a_1586_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18705 VSS pmat.row_n[14] a_39550_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18706 a_11897_2767# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18707 a_43662_14480# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18708 a_43566_20902# pmat.rowoff_n[12] a_43170_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18709 VDD a_22522_50247# a_22475_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1871 a_43170_68178# a_18162_68218# a_43262_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18710 a_41162_15922# a_18162_15516# a_41254_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18711 VDD pmat.rowon_n[0] a_46182_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18712 a_26594_24520# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18713 a_14011_60431# a_10515_61839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18714 VDD nmat.rowon_n[1] a_30118_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18715 vcm a_18162_58178# a_30210_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18716 a_30699_29397# a_13641_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18717 a_6699_76983# a_6975_76823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18718 a_9337_15033# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18719 a_41654_8456# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1872 VDD VSS a_24094_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18720 a_29206_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18721 a_8928_73865# a_7847_73493# a_8581_73461# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18722 a_38242_24552# a_18546_24550# a_38150_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18723 VDD nmat.rowon_n[9] a_20078_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18724 a_44174_10902# pmat.row_n[2] a_44666_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18725 a_17187_49783# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18726 VDD nmat.rowon_n[15] a_51202_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18727 a_4124_28023# a_4339_27804# a_4266_27830# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X18728 a_21082_63158# a_18162_63198# a_21174_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18729 a_27106_20942# pmat.row_n[12] a_27598_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1873 a_45152_48783# a_44870_48437# a_21279_48999# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18730 a_34626_72556# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18731 a_42562_68218# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18732 a_27106_16926# a_18162_16520# a_27198_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18733 vcm a_18162_20536# a_48282_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18734 VDD config_2_in[12] a_1591_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X18735 a_10873_39605# a_30679_40513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X18736 VDD pmat.rowon_n[2] a_37146_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18737 a_31214_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18738 VSS pmat.row_n[0] a_23486_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18739 VDD nmat.rowon_n[15] a_27106_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1874 a_19268_34191# a_19091_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18740 a_34134_62154# a_18162_62194# a_34226_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X18741 a_37542_11866# nmat.rowon_n[12] a_37146_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18742 VSS a_15899_47939# a_15711_47899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18743 a_10575_15253# a_10400_15279# a_10754_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18744 VDD a_1591_31599# a_1683_46295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18745 a_6037_59887# a_4025_54965# a_5939_60137# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X18746 VDD nmat.rowon_n[10] a_24094_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18747 a_21574_10464# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18748 a_33526_8854# nmat.rowon_n[15] a_33130_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18749 a_12543_39453# a_12289_39126# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1875 VSS pmat.row_n[0] a_37542_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18750 a_13054_16367# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18751 a_45574_59182# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18752 pmat.rowoff_n[10] pmat.rowon_n[7] a_14747_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X18753 a_18107_53034# a_18199_52789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18754 a_43170_16926# pmat.row_n[8] a_43662_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18755 a_28506_69222# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18756 VSS pmat.row_n[11] a_32522_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18757 a_19928_37253# a_18769_36965# a_19891_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18758 a_14923_38825# a_13801_38779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18759 a_5747_44655# a_4257_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1876 VDD a_44976_47349# a_44870_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18760 a_19049_41959# a_19145_41781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18761 VDD nmat.rowon_n[4] a_50198_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18762 VSS pmat.row_n[3] a_22482_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18763 a_49590_58178# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18764 VSS a_5785_48463# a_5688_52423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18765 a_28202_61150# a_18546_61192# a_28110_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18766 a_25098_8894# a_18162_8488# a_25190_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18767 a_51202_68178# a_18162_68218# a_51294_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18768 vcm a_18162_68218# a_37238_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18769 a_20078_7890# VDD a_20570_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1877 a_10055_22671# a_8197_20871# a_10209_22351# VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X18770 a_30913_39867# a_29772_40517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X18771 VDD pmat.rowon_n[7] a_32126_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18772 VDD a_1643_74005# a_1591_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18773 a_2163_65469# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18774 a_16966_29673# a_17306_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X18775 VDD a_40837_46261# a_44923_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X18776 a_37238_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18777 a_48282_8488# a_18546_8486# a_48190_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18778 a_12270_30511# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18779 VSS a_31015_29111# a_30603_29575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X1878 a_6975_76823# a_9287_77055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18780 VDD a_19399_48437# a_16800_47213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X18781 a_5205_57533# a_4075_68583# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18782 VSS a_5257_62215# a_4413_62037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18783 VSS pmat.row_n[2] a_26498_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18784 a_20570_60508# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18785 a_23486_55166# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18786 VSS a_6853_14967# a_7253_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18787 a_29114_61150# pmat.row_n[5] a_29606_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18788 a_3514_57167# a_2419_69455# a_3514_57487# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X18789 a_38242_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1879 a_12225_74575# a_10515_75895# a_12153_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X18790 VDD a_23815_50069# pmat.row_n[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X18791 a_26041_36374# a_25209_36965# a_26272_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X18792 a_27198_67174# a_18546_67216# a_27106_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18793 a_13414_17999# a_12337_18005# a_13252_18377# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18794 a_5821_32929# a_5603_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X18795 VDD pmat.rowon_n[13] a_31122_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18796 a_34530_61190# pmat.rowon_n[5] a_34134_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18797 VSS a_4383_7093# a_11987_10089# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18798 VSS a_5363_33551# a_12079_31061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18799 a_5499_19631# a_5351_19913# a_5136_19783# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X188 VSS a_15549_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X1880 VSS a_31701_37462# a_32035_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X18800 a_31214_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18801 a_5541_71855# a_2879_57487# a_5323_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18802 a_35306_47081# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18803 a_8928_56457# a_8013_56085# a_8581_56053# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X18804 VSS VDD a_45574_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18805 a_42562_21906# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18806 a_39154_20942# a_18162_20536# a_39246_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18807 a_12476_51549# a_11807_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18808 VSS a_46811_33927# a_45908_33749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18809 VSS a_31425_37218# a_32035_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X1881 a_6998_8751# a_6956_8965# a_6412_8725# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18810 a_31518_66210# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18811 a_45178_57134# pmat.row_n[1] a_45670_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18812 a_35230_59142# a_18546_59184# a_35138_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18813 vcm a_18162_63198# a_28202_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18814 VSS a_17113_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X18815 a_28110_67174# pmat.row_n[11] a_28602_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18816 vcm a_18162_23548# a_50290_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18817 a_18751_53034# a_18777_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18818 a_49286_16520# a_18546_16518# a_49194_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18819 a_32618_65528# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1882 a_46940_45519# a_7109_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X18820 VDD a_2847_63999# a_2834_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18821 VSS pmat.row_n[8] a_35534_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18822 a_12155_20719# a_11903_20969# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18823 a_24781_52521# ANTENNA__1395__B1.DIODE pmat.col[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X18824 a_4165_71017# a_1591_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18825 a_32126_55126# a_18162_55166# a_32218_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18826 VSS pmat.row_n[7] a_48586_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18827 a_45574_12870# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18828 a_22482_24918# VSS a_22086_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18829 a_22578_57496# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1883 VSS a_10383_13077# a_1781_9308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X18830 a_28506_22910# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18831 a_13361_18377# a_12171_18005# a_13252_18377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18832 vcm a_18162_55166# a_36234_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18833 VSS a_11297_36091# a_35799_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18834 a_7092_74005# a_6795_76989# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18835 a_32126_14918# pmat.row_n[6] a_32618_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18836 vcm a_18162_7484# a_27198_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18837 VSS pmat.row_n[12] a_32522_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18838 a_3661_74941# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18839 a_11773_39087# a_11507_39087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1884 VSS a_13653_40956# a_13345_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X18840 a_36142_59142# pmat.row_n[3] a_36634_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18841 a_5445_73807# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18842 result_out[0] a_1644_53877# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18843 VDD a_34277_37462# a_33341_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X18844 a_13328_55357# a_5682_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18845 pmat.col_n[11] ANTENNA__1184__B1.DIODE a_30561_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18846 a_49194_58138# pmat.row_n[2] a_49686_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18847 a_25494_15882# pmat.rowoff_n[7] a_25098_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18848 VSS pmat.row_n[4] a_22482_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18849 a_1643_65301# a_1846_65579# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1885 a_29114_8894# pmat.row_n[0] a_29606_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18850 a_49590_11866# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18851 VSS a_13837_39069# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X18852 VSS a_5136_19783# a_5087_19319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18853 a_10763_28995# a_9741_28585# a_10691_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18854 vcm a_18162_24552# a_27198_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18855 vcm a_18162_66210# a_26194_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18856 VSS pmat.row_n[6] a_47582_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18857 VDD nmat.rowon_n[14] a_36142_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18858 VDD a_6637_69367# a_5497_62839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X18859 a_51598_60186# pmat.rowon_n[4] a_51202_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1886 a_8919_71615# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18860 a_30210_64162# a_18546_64204# a_30118_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18861 a_51598_19898# nmat.rowon_n[4] a_51202_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18862 VSS a_18272_35077# a_18235_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18863 a_9556_69679# a_9139_68841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18864 a_30610_68540# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18865 VSS a_28591_36519# a_11149_36924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X18866 a_26594_58500# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18867 a_29510_14878# nmat.rowon_n[9] a_29114_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18868 VSS pmat.row_n[3] a_26498_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18869 a_24094_9898# pmat.row_n[1] a_24586_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1887 a_28202_70186# a_18546_70228# a_28110_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18870 VDD VSS a_48190_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18871 VSS a_20475_49783# a_20267_50345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X18872 a_5411_12167# a_4865_12533# a_5645_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18873 VDD a_19928_37253# a_19817_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X18874 VDD a_13273_10357# a_13163_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18875 a_13173_68597# a_10991_68591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18876 a_34626_9460# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18877 vcm a_18162_60186# a_31214_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18878 VSS pmat.row_n[8] a_38546_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18879 a_31122_64162# pmat.row_n[8] a_31614_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1888 a_16926_46261# a_16083_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X18880 a_5351_60663# a_4025_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18881 a_36634_21508# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18882 a_36234_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18883 a_7355_37013# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18884 VDD a_34924_41605# a_34828_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X18885 a_39154_65166# a_18162_65206# a_39246_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18886 a_11417_10927# a_9675_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18887 VSS _1192_.A2 a_82817_25935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18888 a_43262_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18889 a_40158_60146# a_18162_60186# a_40250_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1889 a_35138_10902# a_18162_10496# a_35230_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X18890 a_49686_20504# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18891 a_49286_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18892 a_21082_56130# pmat.row_n[0] a_21574_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18893 a_23090_70186# a_18162_70226# a_23182_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18894 VDD a_9184_51335# a_6979_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X18895 a_24847_39631# a_12228_39605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18896 a_25190_15516# a_18546_15514# a_25098_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18897 vcm a_18162_12504# a_22178_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18898 a_6637_46348# a_4955_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18899 a_39646_12472# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X189 a_14471_3561# a_10883_3303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X1890 a_25098_71190# pmat.row_n[15] a_25590_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18900 a_41162_23954# a_18162_23548# a_41254_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18901 VSS a_5462_62215# a_5257_62215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18902 a_37146_13914# a_18162_13508# a_37238_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18903 VDD nmat.rowon_n[13] a_43170_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18904 a_46578_8854# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18905 a_6063_77295# a_5713_77295# a_5968_77295# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18906 VDD pmat.rowoff_n[12] a_26102_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18907 VSS a_5351_19913# a_13467_21263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X18908 a_41558_68218# pmat.rowon_n[12] a_41162_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18909 a_51294_19532# a_18546_19530# a_51202_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1891 a_25590_20504# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18910 a_29206_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18911 VSS pmat.row_n[14] a_20474_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18912 a_46578_61190# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18913 VSS a_7717_14735# a_21279_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X18914 a_5403_67655# a_6787_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18915 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18916 VSS pmat.row_n[10] a_50594_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18917 a_29510_71230# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18918 vcm a_18162_11500# a_26194_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18919 a_33785_30287# a_31339_31787# a_33567_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1892 a_23648_47753# a_22567_47381# a_23301_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X18920 a_18176_36165# a_17113_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18921 VSS a_5809_51335# a_5731_58951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18922 a_9385_22057# a_5899_21807# a_9313_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18923 VSS a_8356_23671# a_8307_23439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X18924 a_27106_24958# a_18162_24552# a_27198_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18925 a_15660_31029# nmat.en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18926 VDD pmat.rowon_n[10] a_37146_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18927 a_13763_67191# a_13973_66933# a_13909_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X18928 a_11444_55535# a_10815_55785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X18929 a_31214_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1893 VSS a_10378_7637# a_10789_6575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X18930 VSS a_44447_45431# a_42024_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X18931 a_27198_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18932 vcm a_18162_57174# a_51294_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18933 VSS pmat.row_n[5] a_23486_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18934 a_5173_45993# a_4313_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18935 a_20474_17890# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18936 VDD a_7068_11703# a_6853_14967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18937 a_34030_47893# _1154_.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18938 a_51598_14878# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18939 a_38642_62516# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1894 VDD VDD a_32126_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18940 a_43170_67174# a_18162_67214# a_43262_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18941 a_48586_58178# pmat.rowon_n[2] a_48190_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18942 VDD pmat.rowon_n[4] a_42166_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18943 vcm a_18162_59182# a_24186_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18944 VDD a_3571_13627# a_4075_13653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18945 VSS VDD a_37542_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18946 VSS a_12368_35823# a_12474_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18947 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18948 a_24490_16886# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18949 a_33436_44527# a_33259_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1895 VSS pmat.row_n[12] a_40554_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18950 nmat.en_bit_n[0] pmat.en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18951 a_38727_32447# a_38552_32521# a_38906_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18952 a_22086_10902# a_18162_10496# a_22178_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18953 a_82863_64213# _1154_.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X18954 a_19948_51959# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X18955 a_29114_7890# VDD a_29606_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18956 VDD a_10751_71543# a_9279_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X18957 VDD ANTENNA__1395__A1.DIODE a_23759_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18958 a_36538_69222# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18959 a_10569_64489# a_10167_64239# a_10405_64239# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X1896 pmat.rowoff_n[13] a_14839_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X18960 VDD pmat.rowon_n[15] a_32126_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18961 VSS pmat.row_n[11] a_40554_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18962 a_35534_7850# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18963 a_15435_29111# a_15543_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18964 VDD pmat.rowon_n[5] a_28110_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18965 VSS a_2319_69916# a_2250_70045# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18966 a_35230_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18967 VDD a_30255_49783# pmat.col[11] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X18968 a_11990_73309# a_11232_73211# a_11427_73180# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18969 a_37146_58138# a_18162_58178# a_37238_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1897 VDD a_3408_11849# a_3583_11775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18970 a_51694_23516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18971 a_51294_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18972 a_23486_63198# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18973 a_21621_40955# a_19409_40719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X18974 VDD a_2407_49289# a_6877_64822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18975 a_18583_51433# a_18547_51565# a_18511_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18976 VDD VDD a_40158_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18977 a_37146_17930# pmat.row_n[9] a_37638_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18978 VSS pmat.row_n[15] a_37542_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18979 a_26102_11906# a_18162_11500# a_26194_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1898 a_25190_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18980 a_36466_46831# a_30111_47911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18981 a_29036_41831# a_27877_42043# a_28940_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X18982 VDD nmat.rowon_n[5] a_44174_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18983 a_41654_15484# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18984 a_41558_21906# nmat.rowon_n[2] a_41162_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18985 a_7263_42453# a_7088_42479# a_7442_42479# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18986 a_30514_66210# pmat.rowon_n[10] a_30118_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18987 a_8385_51727# a_7907_52031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18988 VSS a_10975_18231# a_10975_17999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18989 VDD a_24374_29941# a_24959_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1899 a_46274_20536# a_18546_20534# a_46182_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18990 a_27198_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18991 a_40467_46261# a_40741_46565# a_40676_46653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18992 a_22482_7850# VDD a_22086_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18993 a_9827_10166# comp_latch a_9368_9991# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18994 a_35230_67174# a_18546_67216# a_35138_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18995 a_42166_11906# pmat.row_n[3] a_42658_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18996 a_27502_64202# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18997 VSS a_35108_39655# a_35071_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18998 a_12353_54223# a_12311_54135# a_11902_56775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X18999 a_13446_14191# a_10515_13967# a_13360_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_10943_8903# a_11051_8903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X190 VSS a_9528_20407# a_9227_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X1900 a_4995_52815# a_5123_52423# a_5081_53135# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.36e+12p pd=1.272e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X19000 a_25098_21946# pmat.row_n[13] a_25590_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19001 a_10070_32143# a_9983_32385# a_9666_32275# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19002 a_49286_24552# a_18546_24550# a_49194_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19003 VDD nmat.rowon_n[9] a_31122_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19004 a_25098_17930# a_18162_17524# a_25190_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19005 a_48282_66170# a_18546_66212# a_48190_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19006 VDD pmat.rowon_n[3] a_35138_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19007 a_82783_53524# _1519_.A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19008 VDD a_27001_30511# a_30085_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19009 VDD a_25647_34343# a_12345_36924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X1901 a_35534_8854# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19010 VDD a_23741_42567# a_23880_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X19011 VSS a_8568_26703# a_20525_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19012 a_28171_35561# a_27049_35515# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19013 a_32126_63158# a_18162_63198# a_32218_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19014 VSS a_11949_21237# a_11897_21263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19015 a_17536_38567# a_16377_38779# a_17440_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19016 a_8459_73865# a_8013_73493# a_8363_73865# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X19017 VDD pmat.rowon_n[2] a_48190_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19018 a_24490_57174# pmat.rowon_n[1] a_24094_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19019 a_48586_11866# nmat.rowon_n[12] a_48190_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1902 a_19417_43990# a_19689_44581# a_20752_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X19020 a_27560_36391# a_26497_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19021 vcm a_18162_63198# a_36234_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19022 a_7369_19407# a_4976_16091# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19023 a_14729_5263# a_10883_3303# nmat.col[7] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19024 a_36142_67174# pmat.row_n[11] a_36634_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19025 a_19488_52423# a_16800_47213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19026 a_28110_12910# pmat.row_n[4] a_28602_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19027 a_7561_22467# a_6817_21807# a_7479_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19028 a_40650_65528# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19029 a_32618_10464# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1903 a_9184_51335# a_7521_47081# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19030 vcm a_18162_62194# a_49286_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19031 a_6829_26703# a_6634_26133# a_6829_27023# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19032 a_49194_66170# pmat.row_n[10] a_49686_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19033 VDD a_5749_30265# a_5779_30006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19034 a_24186_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19035 VSS a_14365_22351# a_14919_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19036 a_50198_61150# pmat.row_n[5] a_50690_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19037 VDD a_3202_29941# a_3160_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19038 a_15048_35077# a_13985_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19039 a_36538_22910# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1904 VDD pmat.rowon_n[6] a_28110_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19040 a_7295_14441# a_5266_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19041 VDD a_3480_17143# a_2467_16341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19042 vcm a_18162_9492# a_42258_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19043 VSS pmat.row_n[12] a_40554_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19044 a_19605_30511# a_19439_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19045 a_30210_72194# a_18546_72236# a_30118_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19046 a_43662_56492# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19047 a_26194_62154# a_18546_62196# a_26102_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19048 a_2163_58941# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19049 VDD pmat.rowon_n[13] a_29114_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1905 a_49590_69222# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19050 a_26594_66532# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19051 a_23090_63158# pmat.row_n[7] a_23582_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19052 VDD a_28915_50959# a_32836_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19053 VDD pmat.rowon_n[8] a_30118_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19054 a_44266_12504# a_18546_12502# a_44174_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19055 a_26102_56130# a_18162_56170# a_26194_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19056 VDD a_12568_35077# a_12472_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X19057 vcm a_18162_68218# a_48282_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19058 a_28202_9492# a_18546_9490# a_28110_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19059 a_4135_61225# a_2727_58470# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1906 VDD a_45589_31599# a_18243_28327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X19060 VSS a_31425_37218# a_30489_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X19061 a_4043_22869# a_2007_25597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X19062 a_30489_40747# a_24833_40719# a_30403_40747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X19063 VDD pmat.rowon_n[0] a_20078_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19064 a_12195_36694# a_12013_36694# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19065 VSS VDD a_38546_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19066 VSS a_13091_18535# a_14839_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X19067 a_6800_22869# a_6651_22895# a_7096_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19068 a_4266_28157# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19069 a_31122_72194# VDD a_31614_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1907 a_50594_64202# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19070 a_42562_70226# pmat.rowon_n[14] a_42166_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19071 a_27106_62154# pmat.row_n[6] a_27598_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19072 a_2319_52789# a_2163_53057# a_2464_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X19073 a_17113_39141# a_13503_39069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X19074 a_48282_11500# a_18546_11498# a_48190_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19075 a_31614_60508# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19076 a_13719_36649# a_14113_36604# a_13779_36595# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X19077 VDD nmat.rowon_n[14] a_44174_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19078 a_49286_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19079 VDD VSS a_24094_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1908 a_22280_52271# ANTENNA__1395__A1.DIODE a_21977_52245# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X19080 VDD a_10985_42044# a_10591_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19081 VDD a_34002_34191# a_34639_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19082 vcm a_18162_20536# a_22178_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19083 a_25190_23548# a_18546_23546# a_25098_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19084 VDD a_10515_75895# a_10699_75119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19085 a_45574_61190# pmat.rowon_n[5] a_45178_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19086 a_5331_13951# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19087 VSS pmat.row_n[9] a_42562_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19088 a_12162_40719# a_12116_40871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19089 a_28506_71230# pmat.rowon_n[15] a_28110_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1909 a_38812_47741# a_38569_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X19090 a_2122_19087# a_1945_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19091 a_2215_27791# a_1591_27797# a_2107_28169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19092 VSS a_20848_38341# a_20811_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19093 a_50290_69182# a_18546_69224# a_50198_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19094 a_24490_10862# nmat.rowon_n[13] a_24094_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19095 a_35036_32375# a_34243_32143# a_35178_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X19096 a_3229_14741# a_3063_14741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19097 nmat.rowon_n[13] a_14839_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19098 a_46274_59142# a_18546_59184# a_46182_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19099 a_6929_17027# a_3305_15823# a_6833_17027# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X191 a_32687_46607# a_7415_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1910 a_7521_19631# a_6821_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19100 vcm a_18162_56170# a_43262_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19101 a_30205_31849# a_27155_31599# a_30121_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.9e+11p pd=2.98e+06u as=0p ps=0u w=1e+06u l=150000u
X19102 a_26459_42657# a_10873_40693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19103 a_49590_60186# pmat.rowon_n[4] a_49194_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19104 a_6842_57711# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19105 VSS pmat.row_n[8] a_46578_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19106 a_49590_19898# nmat.rowon_n[4] a_49194_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19107 a_43566_13874# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19108 a_5325_9269# a_4611_9839# a_5829_9615# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19109 a_50594_14878# nmat.rowon_n[9] a_50198_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1911 a_26773_40955# a_26317_40726# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X19110 a_6435_40303# a_5989_40303# a_6339_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19111 a_42166_9898# a_18162_9492# a_42258_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19112 a_54136_39932# comp.adc_comp_circuit_0.adc_comp_buffer_1.in VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X19113 a_44266_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19114 VDD a_30663_50087# a_45563_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19115 VDD pmat.rowoff_n[12] a_34134_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19116 a_33622_18496# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19117 a_33526_24918# VSS a_33130_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19118 a_30118_15922# pmat.row_n[7] a_30610_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19119 a_27198_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1912 a_19166_22544# a_18546_22542# a_19074_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19120 VSS a_3175_59585# a_3136_59459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19121 a_2748_11837# a_2129_10383# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19122 vcm a_18162_65206# a_51294_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19123 a_51202_69182# pmat.row_n[13] a_51694_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19124 vcm a_18162_55166# a_47278_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19125 a_3476_72399# a_3262_72399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19126 VSS a_36561_38780# a_36253_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19127 VDD a_8491_47911# a_8079_46519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19128 a_47186_59142# pmat.row_n[3] a_47678_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19129 VSS pmat.row_n[10] a_19470_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1913 VDD a_35244_32411# a_44647_35520# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19130 a_23486_16886# nmat.rowon_n[7] a_23090_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19131 a_28442_29199# a_15667_28111# a_28356_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19132 a_28202_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19133 a_30561_29673# a_28812_29575# a_29455_31293# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19134 a_10137_22351# a_9303_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19135 a_15651_37737# a_16045_37692# a_14719_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X19136 a_38642_70548# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19137 vcm a_18162_67214# a_24186_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19138 a_35230_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19139 VDD a_18975_40871# a_18963_41085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1914 VDD a_10216_62985# a_10391_62911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19140 a_35534_69222# pmat.rowon_n[13] a_35138_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19141 a_18546_12502# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X19142 vcm a_18162_17524# a_42258_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19143 VSS a_1643_31573# a_1591_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19144 a_24186_55126# a_18546_55168# a_24094_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19145 a_48282_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19146 a_39647_48767# a_39472_48841# a_39826_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19147 a_24586_59504# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19148 a_83656_2767# _1154_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X19149 a_28336_29967# a_18563_27791# a_28946_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1915 a_29114_70186# pmat.row_n[14] a_29606_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19150 a_9103_73791# a_8928_73865# a_9282_73853# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19151 a_9227_20291# a_4613_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19152 a_2405_17455# a_2228_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19153 VDD a_8581_73461# a_8471_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X19154 a_11829_53359# a_4128_64391# a_11737_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X19155 VDD clk_dig a_12171_18005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19156 VDD a_11435_58791# a_14289_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19157 a_33596_47081# a_32687_46607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19158 a_39550_68218# pmat.rowon_n[12] a_39154_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19159 VSS pmat.row_n[9] a_36538_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1916 VSS pmat.row_n[3] a_43566_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19160 VSS a_9831_74183# a_9655_74216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19161 vcm a_18162_16520# a_46274_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19162 VDD nmat.rowon_n[6] a_36142_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19163 a_50290_14512# a_18546_14510# a_50198_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19164 a_50594_71230# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19165 a_45287_33231# a_45019_38645# a_44888_33205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19166 a_34593_43493# a_33283_42333# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X19167 VSS pmat.row_n[8] a_49590_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19168 VSS pmat.sw a_10147_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X19169 VDD VDD a_49194_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1917 VDD nmat.rowon_n[15] a_40158_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19170 VSS VDD a_45574_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19171 a_47678_21508# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19172 a_47278_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19173 a_33436_34191# a_33259_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19174 a_8121_49257# a_8091_49192# a_7578_48553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X19175 a_37795_29111# a_18563_27791# a_38193_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19176 a_36341_39141# a_35108_39655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X19177 a_6200_70919# a_11397_76457# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19178 VDD a_16478_29423# a_28273_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19179 a_26889_47073# a_26671_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X1918 a_40554_56170# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19180 pmat.col[5] a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X19181 a_38546_9858# nmat.rowon_n[14] a_38150_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19182 a_11427_73180# a_11232_73211# a_11737_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19183 a_50594_9858# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19184 vcm a_18162_18528# a_19166_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19185 a_2215_17999# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19186 VSS pmat.row_n[0] a_39550_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19187 a_32126_56130# pmat.row_n[0] a_32618_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19188 a_23182_16520# a_18546_16518# a_23090_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19189 VSS a_13837_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X1919 a_37146_18934# pmat.row_n[10] a_37638_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19190 a_41254_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19191 vcm a_18162_13508# a_20170_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19192 a_37638_13476# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19193 VDD nmat.rowon_n[12] a_41162_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19194 a_26498_64202# pmat.rowon_n[8] a_26102_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19195 a_26498_9858# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19196 a_29225_37483# a_29159_37607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19197 vcm a_18162_12504# a_33222_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19198 a_41237_28585# a_18563_27791# a_41237_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19199 a_3814_65871# a_3688_65987# a_3410_66003# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X192 VSS pmat.row_n[4] a_35534_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1920 VSS VDD a_37542_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19200 VSS ANTENNA__1184__B1.DIODE a_30473_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19201 VSS a_37820_30485# a_45489_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19202 a_48190_13914# a_18162_13508# a_48282_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19203 a_27198_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19204 VSS a_3305_17999# a_5455_22057# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X19205 VSS a_45253_27221# nmat.col[25] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19206 a_11041_40948# a_11071_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19207 a_44570_62194# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19208 VSS cgen.enable_dlycontrol_in a_24667_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19209 a_26149_27247# a_11067_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1921 a_26102_12910# a_18162_12504# a_26194_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19210 a_12445_12533# a_12227_12937# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X19211 a_27502_72234# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19212 a_1644_54421# a_1591_54991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19213 VSS a_10764_32117# a_10702_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X19214 VSS pmat.row_n[14] a_31518_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19215 a_12375_42895# a_12198_42895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19216 a_22265_28995# a_19405_28853# a_22193_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19217 vcm a_18162_71230# a_45270_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19218 VDD pmat.rowon_n[11] a_35138_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19219 VSS a_1643_52789# a_1591_52815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1922 a_34850_47695# a_33986_47375# a_35186_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X19220 a_47186_7890# a_18162_7484# a_47278_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19221 a_24955_30761# a_20616_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19222 VSS cgen.dlycontrol3_in[0] a_10767_39087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19223 a_45670_24520# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19224 a_35230_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19225 a_3123_27399# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19226 VDD pmat.rowon_n[10] a_48190_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19227 VSS pmat.row_n[6] a_21478_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19228 a_4987_34293# a_4831_34561# a_5132_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X19229 VSS a_3571_13627# a_9319_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1923 a_9826_47375# a_8749_47381# a_9664_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X19230 a_7072_62037# a_7457_62037# a_7201_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X19231 VDD a_4307_35639# a_4517_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19232 a_48282_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19233 VSS pmat.row_n[5] a_34530_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19234 a_35534_22910# nmat.rowon_n[1] a_35138_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19235 VDD a_4533_38279# a_6369_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19236 a_3663_9269# a_5558_9527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19237 VDD a_12604_47080# a_12542_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19238 a_14439_72703# a_14264_72777# a_14618_72765# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19239 VSS a_82971_11989# nmat.col_n[28] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u M=2
X1924 a_41654_16488# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19240 a_22178_71190# a_18546_71232# a_22086_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19241 a_11173_50095# a_11138_50347# a_10703_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19242 vcm a_18162_70226# a_49286_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19243 a_4809_13621# a_4591_14025# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19244 VDD VSS a_22086_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19245 a_46182_20942# pmat.row_n[12] a_46674_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19246 a_46182_16926# a_18162_16520# a_46274_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19247 a_17046_51843# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19248 a_33130_8894# pmat.row_n[0] a_33622_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19249 a_49686_62516# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1925 VSS pmat.row_n[13] a_26498_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19250 a_50290_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19251 vcm a_18162_59182# a_35230_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19252 a_2672_28169# a_1757_27797# a_2325_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19253 a_2217_29973# a_2051_29973# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19254 a_11071_39958# a_11113_39747# a_11071_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19255 VSS a_30489_36893# a_30181_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19256 a_18084_38341# a_17021_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19257 a_39550_21906# nmat.rowon_n[2] a_39154_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19258 a_36142_12910# pmat.row_n[4] a_36634_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19259 a_7009_10927# a_2021_9563# a_5746_11703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1926 a_23486_66210# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19260 a_7164_31421# a_7047_31226# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X19261 a_35534_16886# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19262 a_32405_32463# a_9963_28111# a_32319_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19263 a_40650_10464# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19264 a_26194_70186# a_18546_70228# a_26102_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19265 VSS a_2046_30184# a_4167_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19266 a_19074_22950# pmat.row_n[14] a_19566_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19267 a_33130_10902# a_18162_10496# a_33222_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19268 a_46934_35951# a_43776_30287# a_46848_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19269 a_23090_71190# pmat.row_n[15] a_23582_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1927 a_1644_68021# a_1674_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19270 a_8091_49192# a_8267_49159# a_8477_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19271 a_23582_20504# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19272 VSS a_2244_26935# a_2021_26677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19273 VDD VDD a_30118_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19274 a_7732_52105# a_6817_51733# a_7385_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X19275 a_23182_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19276 a_44266_20536# a_18546_20534# a_44174_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19277 VDD pmat.rowon_n[6] a_26102_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19278 a_26102_64162# a_18162_64202# a_26194_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19279 VDD a_41481_52245# pmat.col[22] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1928 a_30514_67214# pmat.rowon_n[11] a_30118_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19280 a_10591_42089# a_10985_42044# a_10651_42035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X19281 a_3417_47919# a_3151_48285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19282 a_47582_69222# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19283 a_30210_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19284 VSS pmat.row_n[11] a_51598_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19285 a_29282_30287# a_18563_27791# a_28336_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19286 VDD a_13357_37429# a_13769_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X19287 a_4591_14025# a_4075_13653# a_4496_14013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X19288 pmat.rowoff_n[12] a_10055_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X19289 VSS a_12987_26159# a_13013_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1929 VDD a_1923_31743# a_3052_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X19290 a_2007_21482# a_2099_21237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19291 a_3133_72765# a_2655_72373# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19292 a_9463_53511# a_10455_53387# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X19293 a_27106_70186# pmat.row_n[14] a_27598_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19294 a_48190_58138# a_18162_58178# a_48282_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19295 a_16911_51959# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19296 VDD nmat.rowon_n[9] a_29114_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19297 a_22493_31353# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19298 VSS pmat.row_n[3] a_41558_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19299 VDD nmat.rowon_n[15] a_20078_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X193 a_49286_19532# a_18546_19530# a_49194_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1930 VSS a_9411_15831# a_3571_13627# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19300 a_24094_12910# a_18162_12504# a_24186_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19301 VDD a_14497_42658# a_13561_42333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X19302 VSS comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.84e+07u l=3.9e+06u
X19303 a_33986_47375# a_14887_46377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X19304 VSS pmat.row_n[13] a_24490_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19305 a_48190_17930# pmat.row_n[9] a_48682_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19306 VSS a_35499_28023# nmat.col_n[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19307 a_9225_76207# a_9183_76359# a_8539_76181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X19308 a_5713_77295# a_5547_77295# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19309 a_36459_29673# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X1931 VSS a_14371_25071# a_13641_23439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u M=4
X19310 a_39246_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19311 a_11603_28335# a_11159_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19312 VSS pmat.row_n[2] a_45574_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19313 a_42562_55166# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19314 nmat.rowoff_n[9] a_9963_13967# a_12907_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X19315 pmat.rowoff_n[9] a_14460_61225# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X19316 VSS pmat.row_n[12] a_28506_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19317 a_25494_65206# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19318 VSS a_1586_8439# a_1591_15829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19319 a_11525_14433# a_11307_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1932 a_9405_66627# a_9287_65087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19320 VDD a_35186_47375# a_43315_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19321 a_23090_18934# a_18162_18528# a_23182_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19322 a_3704_57487# a_2879_57487# a_3514_57167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19323 a_46274_67174# a_18546_67216# a_46182_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19324 vcm a_18162_64202# a_43262_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19325 a_39154_19938# pmat.row_n[11] a_39646_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19326 a_43170_68178# pmat.row_n[12] a_43662_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19327 a_35399_32509# a_34243_32143# a_35036_32375# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X19328 VDD pmat.rowon_n[13] a_50198_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19329 VDD pmat.rowon_n[3] a_46182_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1933 a_22105_48169# a_20475_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19330 a_22482_58178# pmat.rowon_n[2] a_22086_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19331 VSS a_31339_31787# a_30412_31751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19332 a_50290_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19333 a_25590_61512# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19334 a_28506_56170# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19335 a_33222_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19336 a_30118_66170# a_18162_66210# a_30210_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19337 VSS a_1923_53055# a_1881_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19338 a_2847_20479# a_2672_20553# a_3026_20541# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19339 VSS a_7186_25615# a_7665_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1934 a_27198_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19340 VDD a_31793_41570# a_30857_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X19341 a_19166_69182# a_18546_69224# a_19074_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19342 a_29606_16488# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19343 a_41254_8488# a_18546_8486# a_41162_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19344 VSS a_2468_21959# a_2099_21237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19345 vcm a_18162_63198# a_47278_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19346 a_47186_67174# pmat.row_n[11] a_47678_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19347 a_32827_46805# a_14887_46377# a_33322_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19348 a_51694_65528# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19349 a_51202_55126# a_18162_55166# a_51294_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1935 a_46027_52047# _1194_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X19350 VSS a_2191_27412# a_1895_27962# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X19351 a_20848_36165# a_19689_35877# a_20811_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X19352 a_22459_48463# a_22015_48579# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19353 a_35230_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19354 VDD a_12447_16143# a_14287_57280# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19355 a_41654_57496# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19356 a_47582_22910# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19357 VDD a_27947_41245# a_27913_42333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X19358 a_24186_63158# a_18546_63200# a_24094_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19359 a_51202_14918# pmat.row_n[6] a_51694_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1936 a_22482_8854# nmat.rowon_n[15] a_22086_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19360 VSS pmat.row_n[12] a_51598_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19361 a_24586_67536# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19362 vcm a_18162_15516# a_38242_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19363 VSS a_13357_37429# a_13776_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19364 VSS a_12219_63303# a_12076_62839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19365 a_42258_13508# a_18546_13506# a_42166_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19366 VSS a_11202_55687# a_13181_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19367 a_34134_24958# nmat.en_bit_n[1] a_34626_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19368 VSS a_2411_33749# a_2369_41213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19369 a_2740_13647# a_2526_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1937 a_20474_59182# pmat.rowon_n[3] a_20078_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19370 a_13915_47375# a_13688_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19371 a_2651_29098# a_2743_28853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19372 a_3248_30333# a_2051_29973# a_3052_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19373 a_24094_57134# a_18162_57174# a_24186_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19374 a_16213_29673# a_16025_29469# a_16131_29429# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19375 a_44447_45431# a_44573_45173# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19376 VDD comp.adc_comp_circuit_0.adc_comp_buffer_1.in a_54790_39198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X19377 a_44570_15882# pmat.rowoff_n[7] a_44174_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19378 VSS pmat.row_n[4] a_41558_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19379 VSS pmat.row_n[14] a_24490_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1938 a_9963_13967# a_15747_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X19380 vcm a_18162_24552# a_46274_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19381 a_17397_48463# a_17049_48579# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X19382 VDD a_20695_32447# a_20682_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19383 VSS a_14113_36604# a_13805_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19384 VDD a_79085_39738# a_78898_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19385 VDD pmat.rowon_n[0] a_31122_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19386 a_7479_22467# a_7693_22365# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19387 VSS a_28247_34191# a_29477_36395# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19388 VDD a_16505_40157# a_16111_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19389 VDD a_2563_34837# a_2467_35015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1939 a_44570_55166# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19390 VSS a_28281_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X19391 VSS VDD a_49590_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19392 VSS a_28969_27765# nmat.col[9] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19393 a_13439_74575# a_12815_74581# a_13331_74953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19394 a_12075_24847# a_10959_23983# a_12075_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19395 VSS a_43720_32143# a_46896_44905# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19396 a_1985_76001# a_1674_68047# a_1899_76001# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X19397 a_45670_58500# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19398 VDD a_12003_52815# a_12311_54135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19399 a_3944_28853# clk_dig VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X194 VDD a_12851_28853# a_17702_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X1940 a_12066_3087# ANTENNA__1184__B1.DIODE a_11897_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X19400 VSS pmat.row_n[3] a_45574_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19401 vcm a_18162_7484# a_20170_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19402 a_28631_44265# a_27509_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19403 VDD a_24867_53135# a_29933_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19404 VSS pmat.row_n[13] a_28506_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19405 a_23182_24552# a_18546_24550# a_23090_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19406 vcm a_18162_21540# a_20170_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19407 a_43566_62194# pmat.rowon_n[6] a_43170_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19408 a_4437_6409# a_3247_6037# a_4328_6409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19409 a_26321_46831# a_26155_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1941 a_18546_61192# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X19410 VSS a_6487_5629# a_6448_5755# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19411 VDD a_45064_44807# a_44628_45717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X19412 a_19166_14512# a_18546_14510# a_19074_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19413 a_26498_72234# VDD a_26102_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19414 VDD a_4719_30287# a_9258_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19415 vcm a_18162_20536# a_33222_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19416 a_31097_44581# a_30641_44743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X19417 VDD pmat.rowon_n[2] a_22086_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19418 VDD a_24602_48169# a_25802_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X19419 VSS a_1925_20871# a_1738_20693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1942 a_35230_68178# a_18546_68220# a_35138_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19420 a_22482_11866# nmat.rowon_n[12] a_22086_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19421 a_15747_50069# a_16083_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19422 a_44695_31393# a_43533_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19423 a_8789_60431# a_5651_66975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X19424 VDD a_1643_58773# a_1591_58799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19425 VSS ANTENNA__1190__B1.DIODE a_14458_4399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19426 a_42166_70186# a_18162_70226# a_42258_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19427 a_34530_64202# pmat.rowon_n[8] a_34134_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19428 VDD a_7808_61493# a_7563_63303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X19429 a_30514_59182# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1943 a_27502_65206# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19430 vcm a_18162_12504# a_41254_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19431 a_5805_49007# a_5639_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19432 a_35230_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19433 VSS a_20855_36885# a_19233_38215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19434 a_9761_30511# a_9595_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19435 a_30543_40721# cgen.dlycontrol4_in[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19436 VDD pmat.rowoff_n[12] a_45178_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19437 VSS a_11113_38659# a_14923_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19438 a_12561_57167# a_12613_57141# a_5682_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X19439 VDD a_4533_38279# a_5659_38127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1944 a_4671_23983# a_4516_21531# a_4308_24135# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X19440 a_48282_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19441 a_45178_61150# a_18162_61190# a_45270_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19442 VDD ANTENNA__1190__A1.DIODE a_31303_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19443 VSS a_23395_53135# a_44084_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19444 a_11505_47919# a_10795_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19445 a_28110_71190# a_18162_71230# a_28202_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19446 VSS a_16800_47213# a_17739_50871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19447 a_34530_58178# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19448 VDD pmat.rowoff_n[4] a_35138_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19449 a_8097_24233# a_7779_22583# a_8025_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1945 a_18162_15516# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X19450 a_31695_43439# a_31518_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19451 a_2655_59317# a_2858_59475# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19452 vcm a_18162_68218# a_22178_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19453 a_45432_46983# a_43315_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19454 a_14005_8585# a_12815_8213# a_13896_8585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19455 a_7079_34837# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19456 a_46182_24958# a_18162_24552# a_46274_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19457 a_15916_52277# a_14653_53458# a_15844_52277# VSS sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X19458 a_49686_70548# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19459 a_50290_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1946 a_27598_17492# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19460 vcm a_18162_18528# a_40250_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19461 a_25821_39659# a_25671_40719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19462 vcm a_18162_67214# a_35230_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19463 a_46274_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19464 a_3026_39037# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19465 a_22178_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19466 a_46578_69222# pmat.rowon_n[13] a_46182_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19467 a_49194_60146# a_18162_60186# a_49286_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19468 a_16671_39913# a_12585_40443# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19469 VDD a_43561_47893# a_43591_48246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1947 VSS a_7415_29397# a_33423_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u M=8
X19470 VSS a_6553_53047# a_6559_53903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X19471 VSS pmat.row_n[15] a_25494_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19472 a_43662_8456# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19473 a_27903_50345# a_13091_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19474 VDD nmat.rowon_n[12] a_39154_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19475 a_23182_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19476 a_20078_21946# a_18162_21540# a_20170_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19477 a_13563_24527# a_12463_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19478 a_2882_54991# a_2124_55107# a_2319_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19479 VDD a_1923_53055# a_2464_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1948 a_37739_37737# a_37776_37479# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X19480 VSS a_2747_74549# a_1823_76181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19481 VDD pmat.rowon_n[14] a_26102_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19482 a_19166_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19483 a_20605_40719# a_20179_41046# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19484 a_12449_39605# a_12116_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19485 a_26194_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19486 pmat.row_n[11] a_9963_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X19487 VSS pmat.row_n[9] a_47582_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19488 a_4255_69135# a_3508_69135# a_4037_69109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19489 VSS a_17635_39605# a_17441_40482# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1949 a_13091_28327# a_40415_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X19490 VDD nmat.rowon_n[15] a_29114_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19491 a_19865_46983# nmat.rowon_n[12] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19492 VSS pmat.row_n[0] a_25494_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19493 pmat.col_n[15] a_26891_28327# a_34425_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19494 a_41162_10902# a_18162_10496# a_41254_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19495 VSS VDD a_30514_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19496 a_24094_20942# a_18162_20536# a_24186_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19497 a_4675_54599# a_4259_73807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19498 VDD pmat.rowon_n[6] a_34134_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19499 VSS pmat.row_n[1] a_37542_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X195 VSS pmat.row_n[11] a_35534_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1950 a_4809_13621# a_4591_14025# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X19500 a_2651_8916# config_1_in[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19501 a_19165_28879# a_18973_29199# a_19083_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.57925e+11p ps=2.52e+06u w=1e+06u l=150000u
X19502 a_30118_57134# pmat.row_n[1] a_30610_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19503 a_41558_55166# VSS a_41162_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19504 VDD a_6628_77295# a_6803_77269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19505 a_20170_59142# a_18546_59184# a_20078_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19506 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19507 VDD a_4128_64391# a_10241_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19508 a_45321_30511# a_37820_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19509 VDD pmat.rowon_n[5] a_47186_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1951 a_25098_18934# a_18162_18528# a_25190_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19510 a_39125_47349# a_38907_47753# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X19511 a_34226_16520# a_18546_16518# a_34134_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19512 VSS pmat.row_n[8] a_20474_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19513 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19514 a_12162_64015# a_11883_62063# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19515 VDD a_41573_51701# pmat.col_n[21] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19516 VDD a_6872_8725# a_6956_8965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19517 a_29510_17890# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19518 VDD nmat.rowon_n[4] a_38150_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19519 a_39647_47679# a_39472_47753# a_39826_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1952 VDD pmat.rowoff_n[7] a_31122_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19520 VSS pmat.row_n[7] a_33526_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19521 a_30514_12870# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19522 a_42562_63198# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19523 a_39154_68178# a_18162_68218# a_39246_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19524 VSS a_37827_30793# a_37837_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19525 a_10333_22351# a_10071_17999# a_10209_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19526 vcm a_18162_55166# a_21174_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19527 a_44268_27247# ANTENNA__1190__A1.DIODE a_43965_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X19528 a_21082_59142# pmat.row_n[3] a_21574_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19529 nmat.rowon_n[2] a_14747_7663# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1953 a_48282_67174# a_18546_67216# a_48190_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19530 a_20179_41046# a_20221_40835# a_20179_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19531 a_27106_8894# a_18162_8488# a_27198_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19532 vcm a_18162_72234# a_43262_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19533 a_5410_30877# a_4333_30511# a_5248_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19534 a_22086_7890# VDD a_22578_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19535 a_2557_71855# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19536 a_8356_23671# a_4703_24527# a_8587_23555# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19537 a_40158_22950# pmat.row_n[14] a_40650_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19538 a_34134_58138# pmat.row_n[2] a_34626_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19539 a_7001_13103# a_5579_12394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1954 vcm a_18162_64202# a_45270_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19540 VDD pmat.rowon_n[11] a_46182_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19541 VSS _1184_.A2 a_14729_3311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19542 a_34530_11866# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19543 a_12175_55535# a_6927_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19544 VDD comp.adc_nor_latch_0.NOR_1/A a_55578_39250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19545 a_32618_7452# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19546 a_46274_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19547 VSS pmat.row_n[6] a_32522_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19548 VSS a_16324_36911# a_16430_36911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19549 a_29206_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1955 a_45178_68178# pmat.row_n[12] a_45670_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19550 a_46578_64202# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19551 a_2834_15823# a_1757_15829# a_2672_16201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19552 a_12219_63303# a_12217_66389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X19553 a_26511_52271# ANTENNA__1195__A1.DIODE pmat.col_n[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19554 a_46578_22910# nmat.rowon_n[1] a_46182_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19555 a_1846_55123# a_2163_55233# a_2121_55357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19556 VDD a_2879_57487# a_3859_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19557 a_44174_21946# pmat.row_n[13] a_44666_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19558 VDD a_4403_51701# a_1923_53055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19559 a_44174_17930# a_18162_17524# a_44266_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1956 a_5253_18543# a_5087_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19560 VDD nmat.rowon_n[9] a_50198_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19561 a_27443_32143# a_27498_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19562 VDD a_41926_46983# a_41883_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19563 VSS a_35244_32411# a_44082_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X19564 a_19166_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19565 VDD VSS a_33130_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19566 a_51202_63158# a_18162_63198# a_51294_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19567 a_34611_42089# a_33309_41479# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19568 a_12764_39453# a_12513_39100# a_12543_39126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19569 a_36538_56170# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1957 VDD a_2163_71997# a_2124_72123# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19570 a_25352_31375# a_22628_30485# a_25232_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X19571 a_19470_66210# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19572 a_24638_49159# a_21371_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19573 VSS pmat.row_n[8] a_23486_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19574 a_37638_55488# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19575 vcm a_18162_23548# a_38242_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19576 a_47186_12910# pmat.row_n[4] a_47678_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19577 a_21574_21508# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19578 a_11711_27907# a_5991_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19579 a_10702_32143# a_9983_32385# a_10139_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1958 VSS a_9279_71829# a_9225_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X19580 a_21174_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19581 a_42258_21540# a_18546_21538# a_42166_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19582 a_51694_10464# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19583 a_24094_65166# a_18162_65206# a_24186_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19584 a_4837_45519# a_4700_44655# a_4745_45519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X19585 a_41786_29673# a_28704_29568# a_41703_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X19586 a_34626_20504# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19587 a_34226_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19588 VSS _1224_.X a_45475_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19589 a_6619_56311# a_6175_60039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1959 VDD pmat.rowon_n[3] a_48190_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19590 VSS pmat.row_n[2] a_37542_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19591 a_3484_15101# a_3367_14906# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19592 a_2121_53181# a_1643_52789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19593 a_7109_53359# a_7067_53511# a_5211_57172# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X19594 VDD pmat.rowoff_n[7] a_27106_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19595 a_24586_12472# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19596 a_1927_43541# a_2263_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X19597 a_22086_13914# a_18162_13508# a_22178_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19598 a_45270_62154# a_18546_62196# a_45178_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19599 a_5157_58575# a_4719_30287# a_4719_58255# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X196 VSS a_2046_30184# a_5823_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1960 VSS a_11807_51157# a_4991_69831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X19600 a_45670_66532# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19601 a_42166_63158# pmat.row_n[7] a_42658_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19602 vcm a_18162_7484# a_29206_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19603 a_12491_30511# a_10147_29415# a_12128_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19604 VSS a_13801_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X19605 VSS a_10478_25045# a_9075_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19606 a_4712_27023# a_2952_25045# a_4627_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19607 a_6346_69929# a_6292_69831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19608 a_35138_12910# a_18162_12504# a_35230_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19609 a_3262_72399# a_3175_72641# a_2858_72531# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X1961 a_24490_58178# pmat.rowon_n[2] a_24094_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19610 a_31518_61190# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19611 a_26501_37462# a_25393_38053# a_26515_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X19612 VDD a_1674_68047# a_2695_76757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19613 VSS a_1586_50247# a_12907_54997# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19614 a_37238_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19615 a_28602_11468# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19616 a_6566_55862# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X19617 a_32160_44869# a_31097_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19618 VDD a_23815_28023# nmat.col[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X19619 VSS a_1957_43567# a_11265_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1962 pmat.sw a_3622_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.2e+11p pd=5.5e+06u as=0p ps=0u w=650000u l=150000u M=5
X19620 VDD pmat.rowon_n[10] a_22086_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19621 a_46182_62154# pmat.row_n[6] a_46674_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19622 VDD a_24921_27221# nmat.col_n[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19623 VDD nmat.rowon_n[14] a_38150_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19624 VDD a_30189_48437# a_19283_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X19625 a_50690_60508# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19626 pmat.col_n[0] _1196_.B1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19627 a_50198_9898# pmat.row_n[1] a_50690_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19628 a_25785_49871# a_25743_49783# pmat.rowoff_n[8] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X19629 a_1757_8213# a_1591_8213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1963 VSS VDD a_21478_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19630 a_44266_68178# a_18546_68220# a_44174_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19631 VSS a_5363_33551# a_6651_33239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19632 a_3859_6409# a_3413_6037# a_3763_6409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19633 a_10471_12791# a_2648_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19634 a_26102_9898# pmat.row_n[1] a_26594_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19635 VSS a_2847_38975# a_2781_39049# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X19636 a_4617_38377# a_4533_38279# a_4535_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19637 a_34530_72234# VDD a_34134_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19638 vcm a_18162_60186# a_19166_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19639 a_19074_64162# pmat.row_n[8] a_19566_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1964 VDD a_4987_34293# a_4918_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X19640 vcm a_18162_20536# a_41254_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19641 VSS a_4319_15039# a_3688_17179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19642 a_36545_51727# a_34942_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19643 a_23582_62516# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19644 vcm a_18162_10496# a_37238_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19645 a_2610_22134# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X19646 a_5183_67503# a_4985_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19647 a_26456_38341# a_25393_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19648 a_33526_58178# pmat.rowon_n[2] a_33130_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19649 a_1775_5059# a_1761_7119# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1965 a_4253_42729# a_2419_69455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19650 a_47582_71230# pmat.rowon_n[15] a_47186_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19651 VSS a_2407_49289# a_6877_64822# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19652 a_15163_32375# a_10055_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19653 a_21174_9492# a_18546_9490# a_21082_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19654 VSS a_33436_44527# a_33542_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19655 a_36278_29967# a_35559_30209# a_35715_29941# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X19656 a_41053_29967# a_28704_29568# a_40969_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19657 VSS a_12128_30663# a_10287_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19658 a_10601_65103# a_5651_66975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19659 a_13091_54447# a_13139_54599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1966 a_10147_29415# pmat.sw a_36723_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.8e+11p pd=5.16e+06u as=5.5e+11p ps=5.1e+06u w=1e+06u l=150000u M=2
X19660 a_42258_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19661 VSS a_3571_13627# a_12539_10389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19662 a_6244_71829# a_2407_49289# a_6464_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19663 VDD a_17740_31287# a_16635_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19664 a_2012_33775# a_1775_35113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19665 a_27598_19500# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19666 a_7140_27805# a_7888_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19667 a_26552_43781# a_25393_43493# a_26456_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19668 VDD pmat.rowon_n[0] a_29114_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19669 VDD a_6975_76823# a_9333_76457# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1967 a_12152_66415# a_12217_66389# a_11977_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.95e+11p ps=5.19e+06u w=1e+06u l=150000u
X19670 a_21478_69222# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19671 a_45574_23914# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19672 a_19955_32521# a_19605_32149# a_19860_32509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19673 a_39246_19532# a_18546_19530# a_39154_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19674 a_46274_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19675 a_22086_58138# a_18162_58178# a_22178_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19676 a_36142_71190# a_18162_71230# a_36234_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19677 VSS pmat.row_n[10] a_38546_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19678 a_6785_42479# a_6741_42721# a_6619_42479# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19679 a_18568_51959# a_18547_51565# a_18799_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1968 a_32126_66170# a_18162_66210# a_32218_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19680 a_6754_8751# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19681 a_42562_16886# nmat.rowon_n[7] a_42166_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19682 a_35138_57134# a_18162_57174# a_35230_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19683 VSS a_14691_29575# a_16863_29239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19684 a_22086_17930# pmat.row_n[9] a_22578_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19685 VSS pmat.row_n[15] a_22482_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19686 a_19166_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19687 a_16837_44219# a_15420_44007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X19688 VSS a_10985_44220# a_10677_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19689 VDD a_12875_16341# a_12862_16733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1969 a_13973_66933# a_13979_65087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19690 a_47290_45717# a_47026_45519# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19691 vcm a_18162_57174# a_39246_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19692 a_39307_27791# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19693 a_43262_55126# a_18546_55168# a_43170_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19694 a_43662_59504# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19695 VSS a_16045_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X19696 a_39550_14878# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19697 a_6566_55535# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19698 a_8655_76751# a_8031_76757# a_8547_77129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19699 a_13252_18377# a_12337_18005# a_12905_17973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X197 a_41883_47081# a_42024_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X1970 a_28110_13914# pmat.row_n[5] a_28602_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19700 a_28506_17890# nmat.rowon_n[6] a_28110_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19701 VDD pmat.rowon_n[14] a_34134_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19702 a_26102_16926# pmat.row_n[8] a_26594_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19703 a_23700_36391# a_22541_36603# a_23604_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19704 a_20170_67174# a_18546_67216# a_20078_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19705 a_41558_63198# pmat.rowon_n[7] a_41162_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19706 VDD cgen.dlycontrol4_in[3] a_33395_43455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19707 a_5445_73807# a_4259_73807# a_5363_73807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19708 VSS a_12152_66415# a_12581_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19709 a_34226_24552# a_18546_24550# a_34134_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1971 a_12051_22057# a_5899_21807# a_11979_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19710 a_33222_66170# a_18546_66212# a_33130_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19711 VDD pmat.rowon_n[3] a_20078_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19712 a_14408_51727# a_13739_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19713 a_21174_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19714 a_29206_56130# a_18546_56172# a_29114_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19715 VSS VDD a_39550_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19716 a_4071_48169# a_3978_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.1e+11p pd=2.82e+06u as=0p ps=0u w=1e+06u l=150000u
X19717 a_25647_37607# a_24015_36911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19718 VDD pmat.rowon_n[2] a_33130_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19719 VDD a_7824_31433# a_7999_31359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1972 a_22178_64162# a_18546_64204# a_22086_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19720 a_10932_21959# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19721 VDD ANTENNA__1195__A1.DIODE a_34797_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19722 VSS pmat.row_n[5] a_29510_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19723 VSS a_27001_30511# a_29931_30517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19724 VDD a_36789_52245# pmat.col_n[17] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19725 a_33526_11866# nmat.rowon_n[12] a_33130_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19726 VSS a_33489_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X19727 vcm a_18162_63198# a_21174_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19728 a_21082_67174# pmat.row_n[11] a_21574_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19729 nmat.col_n[20] a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1973 a_32618_11468# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19730 a_79085_40202# a_79181_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19731 VDD a_6559_33767# a_7631_55687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19732 a_51202_56130# pmat.row_n[0] a_51694_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19733 a_17900_35303# a_16837_35515# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19734 vcm a_18162_62194# a_34226_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19735 a_12953_51183# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19736 VDD a_4127_37013# a_4031_37191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19737 a_34134_66170# pmat.row_n[10] a_34626_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19738 a_10707_64783# a_10921_64786# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.331e+11p pd=2.79e+06u as=0p ps=0u w=420000u l=150000u
X19739 a_45574_64202# pmat.rowon_n[8] a_45178_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1974 vcm a_18162_63198# a_49286_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19740 a_39646_23516# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19741 a_39246_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19742 VDD nmat.rowon_n[2] a_43170_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19743 a_21478_22910# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19744 a_46274_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19745 a_43170_62154# a_18162_62194# a_43262_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19746 a_35534_56170# pmat.rowon_n[0] a_35138_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19747 a_46578_72234# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19748 VDD a_24937_43655# a_26272_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X19749 a_13805_43990# a_13985_44581# a_15107_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1975 a_14071_8511# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19750 result_out[14] a_1644_74549# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X19751 cgen.dlycontrol1_in[1] a_1591_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19752 VSS pmat.row_n[14] a_50594_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19753 a_28202_17524# a_18546_17522# a_28110_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19754 VDD VDD a_42166_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19755 VDD pmat.rowoff_n[4] a_46182_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19756 vcm a_18162_68218# a_33222_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19757 a_44266_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19758 VSS pmat.row_n[6] a_40554_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19759 VSS a_7693_22365# a_11159_23145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1976 a_28999_42089# a_27877_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19760 a_7159_58038# a_4843_54826# a_6700_57863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19761 a_5277_57533# a_5211_57172# a_5205_57533# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19762 a_39550_55166# VSS a_39154_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19763 VSS VDD a_23486_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19764 a_12453_55785# a_11202_55687# a_12038_55687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19765 VSS a_33467_46261# a_36265_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X19766 VDD a_4523_21276# a_10651_24617# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19767 a_24490_7850# VDD a_24094_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19768 VSS config_1_in[5] a_1591_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X19769 a_50594_17890# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1977 a_22578_68540# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19770 vcm a_18162_13508# a_29206_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19771 a_47120_43567# a_40105_47375# a_46817_43541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19772 VDD a_3339_59879# a_10291_77269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19773 a_41254_71190# a_18546_71232# a_41162_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19774 a_33222_11500# a_18546_11498# a_33130_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19775 a_14250_8573# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19776 a_37238_61150# a_18546_61192# a_37146_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19777 VDD a_4308_21495# a_4123_20693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19778 VDD a_3325_26159# a_3891_25623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19779 a_6557_40545# a_6339_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1978 a_49194_67174# pmat.row_n[11] a_49686_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19780 a_34226_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19781 a_5541_12559# a_4895_12559# a_5227_13077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X19782 a_2163_69821# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19783 VDD pmat.rowon_n[7] a_41162_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19784 a_4505_40125# a_3325_40847# a_4433_40125# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19785 a_29829_51433# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19786 a_40158_7890# a_18162_7484# a_40250_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19787 VDD a_22787_42325# a_15049_42902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19788 a_30514_61190# pmat.rowon_n[5] a_30118_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19789 VDD a_13479_26935# a_14725_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1979 a_7907_52031# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19790 VDD a_1643_69653# a_1591_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19791 a_45270_70186# a_18546_70228# a_45178_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19792 VSS a_19584_52423# a_21647_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19793 a_42166_71190# pmat.row_n[15] a_42658_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19794 a_12131_71829# a_12249_71311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X19795 a_2820_30333# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19796 a_20499_31274# a_20591_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19797 VDD a_9287_65087# a_9274_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19798 a_38150_61150# pmat.row_n[5] a_38642_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19799 vcm a_18162_19532# a_28202_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X198 a_40315_42089# a_39193_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X1980 a_24186_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19800 a_35138_20942# a_18162_20536# a_35230_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19801 VSS a_78165_39738# a_77978_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19802 a_79722_40050# vcm.sky130_fd_sc_hd__buf_4_3.A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19803 a_7131_64822# a_5307_67655# a_7059_64822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19804 VDD pmat.rowon_n[6] a_45178_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19805 a_3577_70197# a_3710_70455# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19806 a_39013_43655# a_39193_43131# a_40256_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19807 a_31214_59142# a_18546_59184# a_31122_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19808 VSS a_19283_49783# a_22522_50247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19809 a_26194_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1981 a_12658_42895# a_12481_42895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19810 VDD _1224_.X a_24781_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19811 a_10417_20291# a_6821_18543# a_10321_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19812 a_27502_18894# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19813 a_25821_38571# a_25755_38695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19814 a_10707_64783# a_10601_65103# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19815 VSS a_7263_42453# a_4128_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19816 VSS a_2163_55233# a_2124_55107# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19817 a_36687_46831# a_36539_47113# a_36324_46983# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X19818 VSS pmat.row_n[8] a_31518_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19819 VSS a_1923_31743# a_1881_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1982 a_50198_62154# pmat.row_n[6] a_50690_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19820 a_36753_46805# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19821 vcm a_18162_9492# a_44266_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19822 a_36234_22544# a_18546_22542# a_36142_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19823 a_46182_70186# pmat.row_n[14] a_46674_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19824 a_3733_74941# a_3354_74575# a_3661_74941# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X19825 VSS pmat.row_n[13] a_43566_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19826 a_40554_66210# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19827 vcm a_18162_55166# a_32218_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19828 a_32126_59142# pmat.row_n[3] a_32618_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19829 a_2526_13647# a_2439_13889# a_2122_13779# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X1983 a_31072_30083# a_30603_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19830 a_27836_40743# a_26773_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19831 VSS a_23063_36885# a_16981_37462# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19832 a_10822_68841# a_4991_69831# a_10740_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19833 a_8735_54207# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19834 VSS a_4128_46983# a_6837_42255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19835 a_19074_72194# VDD a_19566_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19836 VDD a_3883_65845# a_3814_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19837 VSS a_10814_29111# a_11159_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19838 a_23582_70548# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19839 a_44266_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1984 VSS a_10515_15055# nmat.rowoff_n[13] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19840 a_19566_60508# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19841 a_20170_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19842 a_27198_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19843 a_11823_74895# a_10515_75895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19844 a_8625_73853# a_8581_73461# a_8459_73865# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19845 a_27789_44743# a_27509_44219# a_28631_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X19846 a_20474_69222# pmat.rowon_n[13] a_20078_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19847 a_44570_65206# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19848 a_18546_71232# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X19849 a_44666_17492# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1985 VSS a_4032_64391# a_3609_65015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19850 a_33222_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19851 a_42166_18934# a_18162_18528# a_42258_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19852 a_20568_38567# a_19505_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19853 a_23707_40693# a_23883_40693# a_23835_40719# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19854 VSS a_36324_46983# a_35540_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19855 VSS a_22541_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X19856 VDD a_4032_64391# a_3609_65015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19857 a_24490_68218# pmat.rowon_n[12] a_24094_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19858 VSS pmat.row_n[9] a_21478_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19859 a_47582_56170# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1986 VSS a_2021_26677# a_2879_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X19860 vcm a_18162_16520# a_31214_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19861 VDD nmat.rowon_n[6] a_21082_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19862 VSS a_24638_49159# a_23971_49140# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19863 a_48682_16488# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19864 a_38242_69182# a_18546_69224# a_38150_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19865 a_45178_13914# pmat.row_n[5] a_45670_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19866 a_6681_62927# a_6175_60039# a_6772_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19867 a_13718_68591# a_13279_68841# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X19868 VSS a_28507_52245# pmat.col[9] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19869 a_13443_38007# a_13837_37981# a_13503_37981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X1987 a_46968_45743# a_47290_45717# a_46797_45993# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.435e+12p ps=1.287e+07u w=1e+06u l=150000u M=2
X19870 VSS pmat.row_n[8] a_34530_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19871 a_35630_19500# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19872 a_11713_26819# a_5991_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19873 a_28110_23954# pmat.row_n[15] a_28602_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19874 a_3411_33231# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19875 VDD a_3325_43023# a_3911_44431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19876 a_28110_19938# a_18162_19532# a_28202_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19877 a_1761_4399# a_1591_4399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19878 a_32618_21508# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19879 a_32218_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1988 a_36538_23914# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19880 a_38546_14878# nmat.rowon_n[9] a_38150_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19881 a_35138_65166# a_18162_65206# a_35230_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X19882 a_42987_50345# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19883 nmat.rowoff_n[10] a_10515_13967# a_14094_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19884 a_10409_53903# a_9871_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19885 a_27502_59182# pmat.rowon_n[3] a_27106_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19886 VSS pmat.row_n[0] a_24490_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19887 vcm a_18162_8488# a_33222_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19888 a_35382_34191# a_35205_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19889 VDD a_13837_43421# a_13443_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1989 a_47293_36815# a_47207_35951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X19890 a_2080_61519# a_1643_61493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19891 VDD nmat.rowon_n[7] a_25098_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19892 a_22578_13476# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19893 vcm a_18162_65206# a_39246_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19894 a_44174_9898# a_18162_9492# a_44266_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19895 a_39154_69182# pmat.row_n[13] a_39646_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19896 a_43262_63158# a_18546_63200# a_43170_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19897 vcm a_18162_60186# a_40250_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19898 a_27785_43131# a_27329_42902# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X19899 a_43662_67536# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X199 VDD a_21219_36885# a_21857_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1990 VSS pmat.row_n[13] a_40554_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19900 a_40158_64162# pmat.row_n[8] a_40650_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19901 a_6424_55687# a_5211_57172# a_6566_55862# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X19902 a_33130_13914# a_18162_13508# a_33222_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19903 a_2882_67869# a_2124_67771# a_2319_67740# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19904 a_4487_28157# a_4339_27804# a_4124_28023# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X19905 a_26102_67174# a_18162_67214# a_26194_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19906 VSS VDD a_28506_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19907 VSS pmat.row_n[14] a_43566_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19908 a_42703_46831# a_41926_46983# a_42191_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19909 vcm a_18162_71230# a_30210_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1991 a_4979_38127# a_4535_38377# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X19910 VSS a_9405_66627# a_10226_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19911 VDD pmat.rowon_n[11] a_20078_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19912 a_4680_63669# a_5065_63669# a_4809_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X19913 a_2021_11043# a_3583_11775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19914 a_29206_64162# a_18546_64204# a_29114_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19915 VDD pmat.rowon_n[0] a_50198_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19916 a_30610_24520# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19917 a_29606_68540# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19918 a_6265_37039# a_6099_37039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19919 a_20170_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1992 a_5465_48783# a_5411_48695# a_5383_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19920 a_6607_10615# a_6879_10473# a_6837_10499# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19921 a_2468_21959# a_2683_22089# a_2610_22134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19922 VDD pmat.rowon_n[10] a_33130_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19923 a_21883_48981# a_21923_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X19924 a_12383_40719# a_10927_41245# a_12020_40871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19925 a_33222_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19926 a_20474_22910# nmat.rowon_n[1] a_20078_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19927 a_6621_16885# a_4976_16091# a_7001_17027# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19928 vcm a_18162_70226# a_34226_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19929 a_38242_14512# a_18546_14510# a_38150_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1993 a_2632_51727# a_2195_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19930 a_38546_71230# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19931 VSS a_1586_33927# a_1591_43029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19932 a_45574_72234# VDD a_45178_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19933 a_31122_20942# pmat.row_n[12] a_31614_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19934 a_31122_16926# a_18162_16520# a_31214_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19935 a_34626_62516# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19936 vcm a_18162_10496# a_48282_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19937 nmat.col_n[12] a_12066_3087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19938 a_21082_12910# pmat.row_n[4] a_21574_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19939 a_24490_21906# nmat.rowon_n[2] a_24094_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1994 a_43662_57496# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19940 VSS a_19834_34191# a_20711_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19941 a_25040_30511# a_24861_29673# a_24737_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19942 a_2865_4943# a_2695_4943# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19943 VDD pmat.rowon_n[1] a_27106_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19944 vcm a_18162_22544# a_25190_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19945 a_15530_31965# a_14453_31599# a_15368_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19946 a_12213_53359# a_11737_53359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X19947 a_43566_24918# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19948 VSS a_4579_47919# a_6553_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19949 VDD a_1957_43567# a_11756_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1995 a_49590_22910# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19950 nmat.rowon_n[5] pmat.rowon_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19951 a_27498_32117# a_27340_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19952 a_32522_69222# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19953 a_7321_63151# a_7364_63303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X19954 a_6613_69929# a_5779_71285# a_6179_69831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X19955 nmat.rowon_n[6] a_14460_12265# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19956 a_43971_28487# a_41731_49525# a_44145_28363# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19957 VDD a_44444_32233# a_47839_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19958 a_7259_31433# a_6743_31061# a_7164_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X19959 a_1644_66933# a_1823_66941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1996 a_26194_63158# a_18546_63200# a_26102_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19960 a_27502_12870# pmat.rowoff_n[4] a_27106_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19961 a_39550_63198# pmat.rowon_n[7] a_39154_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19962 a_6087_70919# a_5081_53135# a_6254_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19963 VSS pmat.row_n[4] a_36538_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19964 VSS pmat.row_n[11] a_36538_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19965 VSS a_12020_40871# a_10949_42364# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19966 a_6723_37405# a_6099_37039# a_6615_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19967 VSS pmat.row_n[14] a_19470_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19968 VSS a_10985_37692# a_10677_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19969 a_33130_58138# a_18162_58178# a_33222_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1997 vcm a_18162_60186# a_23182_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19970 vcm a_18162_21540# a_29206_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19971 a_47186_71190# a_18162_71230# a_47278_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19972 VSS a_5351_19913# a_6564_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19973 VSS pmat.row_n[10] a_49590_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19974 a_20078_18934# pmat.row_n[10] a_20570_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19975 VDD a_6830_22895# a_12605_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19976 a_34002_44527# a_33825_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19977 a_6817_51733# a_6651_51733# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19978 a_34277_37462# a_33765_38053# a_34887_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X19979 a_6447_40669# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1998 VSS a_4308_24135# a_3387_22869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19980 vcm a_18162_68218# a_41254_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19981 VDD nmat.rowon_n[1] a_37146_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19982 vcm a_18162_58178# a_37238_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19983 a_33130_17930# pmat.row_n[9] a_33622_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19984 VSS a_17842_27497# a_39209_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19985 VDD pmat.rowon_n[15] a_41162_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19986 a_49194_7890# a_18162_7484# a_49286_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19987 a_4259_67503# a_2727_58470# a_4165_67503# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X19988 VSS a_6700_57863# a_5528_57685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19989 a_41254_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1999 a_7533_19087# a_4976_16091# a_7461_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X19990 VDD a_12079_9615# a_14839_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X19991 a_37638_8456# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19992 a_24186_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19993 a_2107_16201# a_1591_15829# a_2012_16189# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X19994 a_26498_18894# nmat.rowon_n[5] a_26102_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19995 VSS pmat.row_n[2] a_30514_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19996 a_22684_35303# a_22085_36374# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X19997 VDD a_9797_9813# a_9827_10166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19998 VDD a_5271_23447# a_4516_21531# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19999 a_23807_41959# a_21981_34191# a_23981_41835# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_51202_10902# a_18162_10496# a_51294_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20 a_38249_32509# a_38205_32117# a_38083_32521# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X200 VDD a_11149_36924# a_11093_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2000 a_26594_67536# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20000 VDD a_3175_72641# a_3136_72515# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X20001 VSS a_16083_50069# a_17049_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20002 VDD pmat.rowon_n[14] a_45178_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20003 vcm a_18162_69222# a_27198_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20004 a_38242_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20005 cgen.dlycontrol1_in[2] a_1591_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20006 a_31214_67174# a_18546_67216# a_31122_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20007 a_5257_19087# a_5087_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20008 a_24094_19938# pmat.row_n[11] a_24586_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20009 a_27198_57134# a_18546_57176# a_27106_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2001 a_23090_64162# pmat.row_n[8] a_23582_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20010 a_12533_23145# a_10959_23983# a_12449_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X20011 a_2781_39049# a_1591_38677# a_2672_39049# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20012 a_45270_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20013 VSS pmat.row_n[0] a_19470_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20014 a_35138_8894# pmat.row_n[0] a_35630_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20015 a_23021_29199# a_21341_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X20016 a_11823_46973# a_5363_33551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20017 VDD pmat.rowon_n[3] a_31122_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20018 a_28202_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20019 VSS pmat.row_n[6] a_27502_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2002 VSS a_1858_25615# a_2511_25615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X20020 VDD a_20475_49783# a_32411_49559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X20021 VDD a_7797_63151# a_9414_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20022 vcm a_18162_19532# a_36234_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20023 VSS a_45645_45895# a_44635_46025# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20024 VDD a_5329_54965# a_4587_53505# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X20025 VSS pmat.row_n[11] a_39550_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20026 vcm a_18162_63198# a_32218_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20027 a_32126_67174# pmat.row_n[11] a_32618_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20028 vcm a_18162_18528# a_49286_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20029 a_43566_65206# pmat.rowon_n[9] a_43170_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2003 VSS a_16083_50069# a_19487_49159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X20030 vcm a_18162_13508# a_50290_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20031 VDD a_2419_53351# a_4801_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20032 VSS a_78165_40202# a_77978_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20033 a_12613_57141# a_8491_47911# a_13361_56399# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20034 a_28061_36965# a_27605_37127# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X20035 a_29220_37253# a_28061_36965# a_29124_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20036 a_32035_39913# a_30913_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20037 VDD a_2319_61493# a_2250_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20038 a_3894_59343# a_3136_59459# a_3331_59317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20039 a_20170_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2004 VDD pmat.rowon_n[9] a_30118_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20040 a_38737_37479# a_39045_37692# a_38711_37683# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X20041 a_32522_22910# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20042 a_29114_21946# a_18162_21540# a_29206_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20043 a_7247_74031# a_7099_74313# a_6884_74183# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20044 VDD pmat.rowon_n[7] a_39154_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20045 a_12335_12559# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20046 vcm a_18162_15516# a_23182_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20047 VDD nmat.rowon_n[15] a_22086_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20048 a_26194_18528# a_18546_18526# a_26102_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20049 a_46578_56170# pmat.rowon_n[0] a_46182_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2005 a_44266_13508# a_18546_13506# a_44174_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20050 a_2464_70045# a_2250_70045# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20051 VDD a_17996_40743# a_17900_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20052 VSS pmat.row_n[9] a_25494_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20053 VDD a_9195_58951# a_8193_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X20054 a_35230_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20055 a_13807_72399# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20056 a_12267_36694# a_12237_36596# a_12195_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X20057 VSS a_3339_70759# a_7413_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20058 a_6641_6031# a_6337_6825# a_6559_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20059 vcm a_18162_24552# a_31214_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2006 a_13782_10383# a_12705_10389# a_13620_10761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20060 VSS pmat.row_n[6] a_51598_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20061 a_4174_47158# a_4128_46983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20062 a_3300_19453# a_3183_19258# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20063 vcm a_18162_14512# a_27198_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20064 a_48282_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20065 a_3410_66003# a_3727_66113# a_3685_66237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20066 VDD a_5651_66975# a_5423_67191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20067 vcm a_18162_56170# a_26194_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20068 VSS a_33489_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20069 VSS VDD a_34530_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2007 VDD a_1923_69823# a_2655_72373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20070 a_3111_53333# a_3199_53877# a_2971_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X20071 a_21970_48071# a_21279_48999# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20072 VDD pmat.rowon_n[13] a_38150_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20073 a_30610_58500# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20074 VSS a_10873_39605# a_11292_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20075 a_26498_13874# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20076 a_6990_59049# a_5462_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20077 VSS pmat.row_n[3] a_30514_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20078 VDD a_4025_54965# a_5939_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20079 a_38242_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2008 a_51598_71230# pmat.rowon_n[15] a_51202_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20080 a_4809_63695# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20081 a_20078_8894# a_18162_8488# a_20170_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20082 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20083 VSS a_18180_38341# a_18143_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20084 VSS a_32371_50247# a_32319_50345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20085 a_21037_43658# cgen.start_conv_in VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X20086 a_5779_58038# a_5528_57685# a_5320_57863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20087 a_5779_71285# a_6787_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X20088 a_36142_23954# pmat.row_n[15] a_36634_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20089 a_40158_72194# VDD a_40650_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2009 a_26102_57134# a_18162_57174# a_26194_57134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20090 a_36142_19938# a_18162_19532# a_36234_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20091 VSS a_25117_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20092 a_40650_21508# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20093 a_39646_65528# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20094 a_40250_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20095 a_43262_8488# a_18546_8486# a_43170_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20096 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20097 a_49194_22950# pmat.row_n[14] a_49686_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20098 a_27877_42043# a_27421_41814# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20099 a_39154_55126# a_18162_55166# a_39246_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X201 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u M=325
X2010 VSS nmat.sample_n a_18162_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X20100 VSS pmat.row_n[7] a_28506_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20101 VSS a_3923_68021# a_12993_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20102 a_25494_60186# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20103 a_25494_19898# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20104 a_30527_31573# a_31263_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20105 VSS a_8175_63669# a_1823_66941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20106 VDD a_33341_38780# a_32947_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20107 a_10167_64239# a_5363_70543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20108 a_39154_14918# pmat.row_n[6] a_39646_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20109 VSS pmat.row_n[12] a_39550_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2011 a_33281_49551# a_28915_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X20110 a_43662_12472# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20111 a_29206_72194# a_18546_72236# a_29114_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20112 VDD a_12175_27221# a_12053_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.85e+11p ps=3.57e+06u w=1e+06u l=150000u
X20113 a_41162_13914# a_18162_13508# a_41254_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20114 a_20170_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20115 a_26594_22512# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20116 a_47278_22544# a_18546_22542# a_47186_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20117 VDD a_31339_31787# a_31393_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20118 VDD pmat.rowoff_n[12] a_30118_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20119 cgen.dlycontrol2_in[3] a_1591_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2012 a_30210_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20120 a_33222_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20121 a_30118_61150# a_18162_61190# a_30210_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20122 VDD nmat.rowon_n[6] a_19074_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20123 a_2629_56623# a_2250_56989# a_2557_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20124 VDD pmat.rowoff_n[4] a_20078_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20125 a_14460_11177# nmat.rowon_n[7] a_14287_10927# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20126 VSS a_9963_13967# pmat.rowon_n[3] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X20127 a_16377_38779# a_15921_38550# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20128 a_31122_24958# a_18162_24552# a_31214_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20129 VDD a_12197_41570# a_11261_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X2013 VSS pmat.row_n[4] a_43566_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20130 a_27106_14918# a_18162_14512# a_27198_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20131 a_4768_16055# a_4976_16091# a_4910_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20132 a_33047_41001# a_31925_40955# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20133 a_34626_70548# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20134 a_9109_22467# a_7779_22583# a_9037_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20135 VSS a_45345_31029# a_34204_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20136 VSS a_7109_29423# a_45645_45895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20137 a_42658_18496# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20138 a_3621_58255# a_3746_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20139 a_31214_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2014 a_22015_28995# a_10441_21263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X20140 a_3894_72399# a_3175_72641# a_3331_72373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20141 a_11021_42619# a_13985_41317# a_15048_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20142 a_31518_69222# pmat.rowon_n[13] a_31122_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20143 a_30050_30083# a_25681_28879# a_29968_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20144 a_34134_60146# a_18162_60186# a_34226_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X20145 a_12500_31421# a_5535_29980# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X20146 a_12267_36367# a_12013_36694# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20147 VSS ANTENNA__1187__B1.DIODE a_13717_5263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20148 a_4611_9839# a_4338_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20149 a_7072_26311# a_7186_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.6975e+11p pd=2.13e+06u as=0p ps=0u w=650000u l=150000u
X2015 a_9333_76457# a_6795_76989# a_8539_76181# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X20150 a_40352_41831# a_39193_42043# a_40256_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20151 VSS ANTENNA__1395__B1.DIODE a_24861_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20152 VDD nmat.rowon_n[12] a_24094_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20153 a_18869_46831# a_18521_46837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X20154 vcm a_18162_7484# a_22178_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20155 a_45574_57174# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20156 a_28506_67214# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20157 a_32218_7484# a_18546_7482# a_32126_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20158 VSS pmat.row_n[9] a_32522_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20159 a_18546_68220# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X2016 a_8413_64061# a_8378_63827# a_8175_63669# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20160 a_49286_69182# a_18546_69224# a_49194_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20161 VDD a_3339_59879# a_11572_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20162 a_46674_19500# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20163 a_10373_30511# a_10329_30753# a_10207_30511# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20164 a_25393_41317# a_24937_41479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20165 a_21087_39913# a_19965_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20166 a_7339_32509# a_5179_31591# a_6976_32375# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20167 a_20078_69182# a_18162_69222# a_20170_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20168 VSS pmat.row_n[1] a_22482_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20169 a_20267_50345# a_19584_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2017 VDD a_37827_30793# a_38299_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X20170 a_2100_44343# a_1739_47893# a_2242_44477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20171 a_39003_48841# a_38557_48469# a_38907_48841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20172 a_28602_63520# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20173 a_2882_31965# a_2124_31867# a_2319_31836# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20174 VDD pmat.rowon_n[5] a_32126_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20175 a_11793_59663# a_11007_58229# a_10190_60663# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20176 a_14261_44219# a_13805_43990# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X20177 VDD a_20184_46983# nmat.rowon_n[12] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20178 VDD nmat.rowon_n[4] a_23090_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20179 a_10953_34951# a_11133_34427# a_12196_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2018 VDD pmat.rowon_n[1] a_20078_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20180 a_41162_58138# a_18162_58178# a_41254_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20181 a_1644_74549# a_1823_74557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20182 a_82817_25935# _1192_.B1 nmat.col[26] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20183 a_24094_68178# a_18162_68218# a_24186_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20184 a_2651_8916# config_1_in[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20185 VSS a_2263_43719# a_39169_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20186 VSS a_9135_22057# a_8197_20871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20187 a_7878_62723# a_7212_62607# a_7796_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20188 VSS a_17902_43439# a_21815_42351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20189 VSS a_22085_42902# a_23571_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X2019 VSS pmat.row_n[14] a_26498_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20190 a_44811_36469# a_44647_36201# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X20191 a_41162_17930# pmat.row_n[9] a_41654_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20192 VSS pmat.row_n[15] a_41558_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20193 a_38242_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20194 VDD a_11261_37981# a_10867_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20195 a_34002_34191# a_33825_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20196 a_27198_65166# a_18546_65208# a_27106_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20197 a_27598_69544# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20198 a_12228_39605# a_17459_37143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X20199 VDD pmat.rowon_n[11] a_31122_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X202 a_35224_50613# a_26891_28327# a_35353_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X2020 a_33839_46805# a_39647_48767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20200 a_34530_18894# nmat.rowon_n[5] a_34134_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20201 VSS a_20572_40517# a_20535_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20202 a_32371_47349# a_11067_30287# a_32802_47695# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X20203 a_27106_59142# a_18162_59182# a_27198_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20204 a_13467_21263# a_4523_21276# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20205 a_17927_47349# a_18083_47593# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X20206 a_6432_67503# a_3866_57399# a_6242_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20207 VSS a_31978_43439# a_33259_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20208 VSS a_2944_65576# a_2882_65693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20209 VSS a_25931_27221# nmat.col[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2021 a_5711_18909# a_5087_18543# a_5603_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X20210 a_31214_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20211 a_30278_30511# a_29931_30517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X20212 a_47582_17890# nmat.rowon_n[6] a_47186_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20213 a_23455_32447# a_23280_32521# a_23634_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20214 a_41558_8854# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20215 a_45670_8456# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20216 a_31518_64202# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20217 a_45178_55126# VDD a_45670_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20218 a_35230_57134# a_18546_57176# a_35138_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20219 a_10395_51183# a_9427_50095# a_10205_51433# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X2022 a_30610_14480# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20220 a_3613_19061# a_3395_19465# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X20221 a_31518_22910# nmat.rowon_n[1] a_31122_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20222 VDD a_6141_44629# a_6059_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.1e+11p ps=2.82e+06u w=1e+06u l=150000u
X20223 a_28110_65166# pmat.row_n[9] a_28602_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20224 vcm a_18162_21540# a_50290_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20225 VSS pmat.row_n[0] a_51598_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20226 VDD a_5589_14967# a_5547_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X20227 VSS pmat.row_n[6] a_35534_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20228 a_49286_14512# a_18546_14510# a_49194_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20229 VSS a_18563_27791# a_40129_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2023 a_30514_20902# pmat.rowoff_n[12] a_30118_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20230 a_48282_56130# a_18546_56172# a_48190_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20231 a_26497_36603# a_26041_36374# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20232 a_21478_56170# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20233 a_7644_16341# a_10575_15253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X20234 VSS a_11167_11177# a_11501_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20235 VDD a_23807_41959# a_12116_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X20236 a_20503_48981# a_20659_49140# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X20237 VSS pmat.row_n[5] a_48586_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20238 a_5253_32687# a_5087_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20239 a_45574_10862# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2024 VSS _1192_.A2 a_83005_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20240 a_11271_73085# a_7658_71543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20241 VDD a_17187_49783# a_17139_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X20242 VDD pmat.rowon_n[15] a_39154_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20243 a_22578_55488# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20244 VDD a_4298_67191# a_4255_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20245 a_28506_20902# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20246 vcm a_18162_23548# a_23182_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20247 a_32126_12910# pmat.row_n[4] a_32618_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20248 a_10052_52047# a_9335_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20249 VDD a_6316_8903# a_5654_9527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2025 VDD a_17996_41831# a_17900_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X20250 a_8133_46607# a_8079_46519# a_8051_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20251 a_12162_41046# a_12116_40871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20252 VSS a_8727_70197# a_7658_71543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X20253 a_25494_13874# nmat.rowon_n[10] a_25098_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20254 VSS pmat.row_n[2] a_22482_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20255 a_9869_69921# a_9651_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20256 VSS a_2835_13077# a_12489_12925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20257 a_45178_72194# a_18162_72234# a_45270_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20258 VSS pmat.row_n[4] a_47582_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20259 vcm a_18162_64202# a_26194_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2026 a_10575_15253# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20260 VSS pmat.row_n[11] a_47582_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20261 VDD VDD a_36142_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20262 a_26102_68178# pmat.row_n[12] a_26594_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20263 a_30210_62154# a_18546_62196# a_30118_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20264 VSS a_7255_71829# a_6602_72007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20265 a_37542_66210# pmat.rowon_n[10] a_37146_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20266 a_6522_18543# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20267 VDD a_47211_50069# a_11067_27239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X20268 a_30610_66532# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20269 a_11041_39860# a_11347_40214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2027 VDD pmat.rowon_n[0] a_33130_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20270 a_4037_66933# a_3983_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20271 VDD pmat.rowoff_n[15] a_35138_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20272 VDD pmat.rowon_n[3] a_29114_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20273 a_29114_8894# a_18162_8488# a_29206_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20274 a_39105_40743# a_39413_40956# a_39079_40947# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X20275 a_24094_7890# VDD a_24586_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20276 VSS a_3339_59879# a_13961_72765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X20277 a_11241_28585# a_9741_28585# a_11159_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20278 VDD nmat.rowon_n[1] a_48190_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20279 vcm a_18162_58178# a_48282_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2028 VDD ANTENNA__1197__A.DIODE a_28810_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X20280 a_40591_38007# a_39469_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20281 a_22178_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20282 a_11021_43011# a_19689_42405# a_20752_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20283 pmat.row_n[11] a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X20284 a_34626_7452# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20285 a_30514_7850# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20286 VDD a_1957_43567# a_10703_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20287 a_4253_42729# a_2659_35015# a_4253_42479# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20288 a_24131_29967# a_23043_28335# a_24214_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20289 VSS a_1643_67477# a_1591_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2029 a_38150_9898# pmat.row_n[1] a_38642_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20290 a_31122_62154# pmat.row_n[6] a_31614_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20291 VDD nmat.rowon_n[9] a_38150_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20292 a_36234_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20293 a_20354_27247# a_8568_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20294 a_5897_38127# a_5687_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20295 a_39154_63158# a_18162_63198# a_39246_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20296 a_50198_21946# a_18162_21540# a_50290_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20297 a_4307_35639# a_2659_35015# a_4345_34863# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X20298 a_49286_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20299 VSS a_12568_35077# a_12531_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X203 VSS pmat.row_n[1] a_28506_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2030 a_19470_17890# nmat.rowon_n[6] a_19074_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20300 a_35138_19938# pmat.row_n[11] a_35630_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20301 a_37749_47081# a_35186_47375# a_37654_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20302 pmat.col_n[28] a_46934_52047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20303 a_9577_28335# a_4339_27804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20304 a_39301_52521# _1224_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20305 a_25190_13508# a_18546_13506# a_25098_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20306 vcm a_18162_10496# a_22178_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20307 a_39646_10464# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20308 VSS a_11965_42583# a_11910_43047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20309 a_32522_71230# pmat.rowon_n[15] a_32126_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2031 a_17536_38567# a_16377_38779# a_17499_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X20310 a_14825_50095# a_14287_50345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20311 VSS pmat.row_n[12] a_37542_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20312 vcm a_18162_19532# a_47278_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20313 VDD a_23821_35279# a_29051_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20314 a_4123_16042# a_4215_15797# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20315 a_39015_47375# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X20316 VSS a_31793_41570# a_39387_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20317 a_29206_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20318 a_50290_59142# a_18546_59184# a_50198_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20319 a_11885_27497# a_5351_19913# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 a_9953_54223# a_9581_56079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X20320 a_2325_27765# a_2107_28169# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20321 a_40532_43781# a_39469_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20322 a_46578_18894# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20323 a_3415_9839# a_3142_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20324 a_16113_52271# a_15757_52535# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20325 VSS pmat.row_n[8] a_50594_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20326 vcm a_18162_9492# a_38242_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20327 a_17635_39605# a_12969_40175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20328 VSS a_18975_40871# a_20400_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20329 VDD a_10391_69653# a_10378_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2033 a_8452_77117# a_6292_69831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X20330 a_30514_23914# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20331 a_27106_22950# a_18162_22544# a_27198_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20332 VSS _1154_.A a_46804_51433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20333 VDD a_10651_44211# a_10677_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20334 VDD pmat.rowon_n[8] a_37146_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20335 a_31214_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20336 a_24186_19532# a_18546_19530# a_24094_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20337 a_42258_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20338 VDD a_4043_33535# a_4030_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20339 a_28907_43177# a_27785_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2034 VDD a_3207_65845# a_1823_68565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20340 VSS a_11067_64015# a_19488_52423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20341 a_19470_61190# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20342 a_4032_46983# a_2389_45859# a_4174_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X20343 vcm a_18162_55166# a_51294_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20344 a_21082_71190# a_18162_71230# a_21174_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20345 a_16285_29673# a_12437_28879# a_16213_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20346 a_51202_59142# pmat.row_n[3] a_51694_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20347 a_20474_15882# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20348 VSS pmat.row_n[10] a_23486_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20349 a_6829_27023# a_5320_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2035 VDD ANTENNA__1190__A1.DIODE a_40040_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.55e+11p ps=2.51e+06u w=1e+06u l=150000u
X20350 VDD a_31596_34191# a_31702_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20351 pmat.rowon_n[5] a_10515_13967# a_14738_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20352 a_33765_35877# a_33309_36039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20353 a_9207_47375# a_8583_47381# a_9099_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20354 VDD a_2672_43401# a_2847_43327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20355 a_38642_60508# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20356 a_46274_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20357 vcm a_18162_57174# a_24186_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20358 a_11881_16911# a_11711_16911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20359 VDD a_7999_31359# a_4259_31375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2036 a_20474_12870# pmat.rowoff_n[4] a_20078_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20360 VSS a_7693_22365# a_8859_22467# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20361 VDD a_45450_48695# a_45546_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20362 a_24490_14878# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20363 a_6639_23413# pmat.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20364 a_43170_24958# VDD a_43662_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20365 a_3879_42997# a_2021_26677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20366 VDD a_28189_37981# a_27795_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20367 a_28602_71552# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20368 a_36538_67214# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20369 a_49286_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2037 nmat.en_bit_n[2] pmat.en_bit_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X20370 a_10949_43124# a_10979_42390# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20371 VSS pmat.row_n[9] a_40554_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20372 a_9463_50877# a_9135_49257# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20373 VDD nmat.rowon_n[6] a_40158_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20374 a_7096_23145# a_7048_23277# a_7012_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20375 VDD a_3337_22325# a_3227_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20376 a_49590_66210# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20377 a_2319_74268# a_2163_74173# a_2464_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20378 a_23182_9492# a_18546_9490# a_23090_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20379 a_47186_23954# pmat.row_n[15] a_47678_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2038 vcm a_18162_7484# a_40250_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20380 VSS a_6283_31591# a_28455_47381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20381 a_47186_19938# a_18162_19532# a_47278_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20382 a_14578_51727# a_14452_51843# a_14174_51859# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20383 a_51694_21508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20384 VSS a_2375_16532# a_1895_15994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X20385 a_51294_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20386 VSS a_39781_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20387 VSS pmat.row_n[0] a_43566_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20388 a_37146_15922# pmat.row_n[7] a_37638_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20389 VSS pmat.row_n[13] a_37542_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2039 a_32035_43177# a_32072_42919# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X20390 a_38150_9898# a_18162_9492# a_38242_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20391 VDD nmat.rowon_n[7] a_44174_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20392 a_41654_13476# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20393 a_3119_22729# a_2603_22357# a_3024_22717# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X20394 a_29510_69222# pmat.rowon_n[13] a_29114_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20395 VSS pmat.row_n[10] a_26498_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20396 a_30514_64202# pmat.rowon_n[8] a_30118_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20397 VDD a_28507_52245# pmat.col[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X20398 a_24586_23516# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20399 a_24186_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X204 a_46182_71190# a_18162_71230# a_46274_71190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2040 a_38546_61190# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20400 a_31214_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20401 a_27198_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20402 a_20474_56170# pmat.rowon_n[0] a_20078_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20403 a_22879_41781# a_10949_42364# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20404 a_31518_72234# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20405 a_35230_65166# a_18546_65208# a_35138_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20406 a_11897_21813# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20407 a_35630_69544# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20408 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20409 a_27598_14480# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2041 VDD a_4976_16091# a_10305_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X20410 a_13163_10383# a_12539_10389# a_13055_10761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20411 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20412 a_14943_26703# a_14725_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X20413 a_25098_15922# a_18162_15516# a_25190_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20414 a_28202_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20415 VSS a_29217_41570# a_28281_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X20416 VDD pmat.rowoff_n[4] a_31122_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20417 a_48282_64162# a_18546_64204# a_48190_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20418 vcm a_18162_61190# a_45270_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20419 a_48682_68540# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2042 a_8851_63669# a_8656_63811# a_9161_64061# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X20420 VSS a_6343_18517# a_6277_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20421 a_9749_19061# a_7644_16341# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20422 a_7131_65149# a_6877_64822# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20423 a_24490_55166# VSS a_24094_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20424 a_12245_31061# a_12079_31061# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20425 a_8079_46519# a_8907_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20426 VDD a_11067_27239# a_35167_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20427 VSS a_10147_29415# a_36278_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20428 a_3960_19465# a_3045_19093# a_3613_19061# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X20429 a_36142_65166# pmat.row_n[9] a_36634_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2043 vcm a_18162_21540# a_22178_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20430 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=5.1e+06u w=1.89e+07u
X20431 a_28110_10902# pmat.row_n[2] a_28602_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20432 a_20629_30511# a_19439_30511# a_20520_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X20433 a_43566_58178# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20434 VSS a_26501_37462# a_26515_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20435 a_22178_61150# a_18546_61192# a_22086_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20436 a_9835_15279# a_9319_15279# a_9740_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X20437 a_12815_26409# a_11927_27399# a_12987_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X20438 VSS a_12851_28853# a_12407_28853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20439 vcm a_18162_60186# a_49286_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2044 a_25190_24552# a_18546_24550# a_25098_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20440 a_27618_27247# a_18243_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20441 a_41593_49871# a_30663_50087# a_34705_51959# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X20442 VDD pmat.rowon_n[12] a_25098_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20443 a_49194_64162# pmat.row_n[8] a_49686_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20444 a_7729_22467# a_7693_22365# a_7657_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20445 a_23182_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20446 a_37960_42693# a_36801_42405# a_37923_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20447 VDD a_2839_38101# a_3431_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20448 VDD clk_ena a_20787_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20449 a_9020_7497# a_8105_7125# a_8673_7093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2045 a_8275_71689# a_7829_71317# a_8179_71689# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X20450 a_36538_20902# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20451 a_3105_11837# a_3061_11445# a_2939_11849# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X20452 vcm a_18162_72234# a_26194_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20453 a_39154_56130# pmat.row_n[0] a_39646_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20454 a_30210_70186# a_18546_70228# a_30118_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20455 a_2369_28157# a_2325_27765# a_2203_28169# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20456 vcm a_18162_22544# a_44266_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20457 a_26194_60146# a_18546_60188# a_26102_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20458 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20459 VDD pmat.rowon_n[11] a_29114_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2046 a_45574_62194# pmat.rowon_n[6] a_45178_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20460 a_26594_64524# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20461 a_23090_61150# pmat.row_n[5] a_23582_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20462 VDD pmat.rowon_n[6] a_30118_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20463 a_44266_10496# a_18546_10494# a_44174_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20464 VDD a_22963_35041# a_22787_34709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20465 a_51598_69222# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20466 a_12247_20175# a_11995_20291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X20467 a_2985_74941# a_2950_74707# a_2747_74549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20468 a_15549_39867# a_15093_39638# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X20469 a_13723_3087# a_10883_3303# nmat.col[1] VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X2047 a_6557_35105# a_6339_34863# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X20470 a_29510_22910# nmat.rowon_n[1] a_29114_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20471 VSS pmat.row_n[14] a_38546_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20472 a_14035_39958# a_13853_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20473 a_21174_22544# a_18546_22542# a_21082_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20474 a_31122_70186# pmat.row_n[14] a_31614_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20475 VSS a_2411_33749# a_2369_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20476 a_22874_28585# a_20616_27791# a_22792_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20477 a_27106_60146# pmat.row_n[4] a_27598_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20478 a_36234_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20479 a_9675_10396# a_13795_10687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2048 VSS a_17996_40743# a_17959_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X20480 a_4591_28335# a_4241_28335# a_4496_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20481 a_35138_68178# a_18162_68218# a_35230_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20482 a_23883_40693# a_12116_40871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20483 VSS a_12500_68021# a_9545_66567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X20484 a_2250_70045# a_2163_69821# a_1846_69931# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20485 VDD VDD a_44174_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20486 VSS VDD a_40554_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20487 a_6787_55535# a_5211_57172# a_6424_55687# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X20488 a_49286_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20489 VDD a_3339_59879# a_10751_72917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2049 a_40158_71190# a_18162_71230# a_40250_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20490 VSS a_2199_13887# a_4025_6397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20491 VSS a_2944_59048# a_2882_59165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20492 a_3423_74549# a_3228_74691# a_3733_74941# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X20493 a_50594_7850# VDD a_50198_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20494 a_38546_17890# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20495 a_25190_21540# a_18546_21538# a_25098_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20496 a_43262_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20497 a_45574_18894# nmat.rowon_n[5] a_45178_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20498 a_5455_22057# a_3305_15823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20499 VSS pmat.row_n[7] a_42562_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 a_32126_58138# a_18162_58178# a_32218_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2050 a_31122_10902# pmat.row_n[2] a_31614_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20500 VSS a_19873_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20501 a_21478_9858# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20502 nmat.col_n[31] ANTENNA__1197__A.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20503 a_9664_47753# a_8583_47381# a_9317_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20504 VDD a_10575_15253# a_10562_15645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20505 a_12248_42583# a_12344_42325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20506 vcm a_18162_69222# a_46274_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20507 a_14460_60137# a_10239_14183# a_14369_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20508 a_11204_71855# a_10699_72943# a_11104_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X20509 a_50290_67174# a_18546_67216# a_50198_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2051 VSS pmat.row_n[10] a_42562_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20510 VSS pmat.row_n[1] a_31518_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20511 a_46274_57134# a_18546_57176# a_46182_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20512 a_5991_23983# a_5547_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X20513 a_7819_25731# a_7779_22583# a_7747_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20514 a_9556_69679# a_9139_68841# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20515 a_43170_58138# pmat.row_n[2] a_43662_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20516 VSS a_7040_8725# a_6998_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20517 VDD pmat.rowon_n[3] a_50198_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20518 a_40371_31393# a_39939_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20519 VSS pmat.row_n[6] a_46578_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2052 a_39013_42693# a_38737_41814# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X20520 a_43566_11866# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20521 a_14107_39631# a_13853_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20522 a_12020_40871# a_10927_41245# a_12162_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20523 a_7364_63303# a_7796_62723# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X20524 a_42166_7890# a_18162_7484# a_42258_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20525 a_32522_56170# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20526 a_4517_35407# a_4257_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20527 VDD VDD a_37146_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20528 a_29114_18934# pmat.row_n[10] a_29606_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20529 VSS VDD a_29510_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2053 a_28506_72234# VDD a_28110_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20530 VSS a_4399_51157# a_4075_68583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X20531 a_23182_69182# a_18546_69224# a_23090_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20532 vcm a_18162_66210# a_20170_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20533 a_33622_16488# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20534 a_30118_13914# pmat.row_n[5] a_30610_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20535 VSS a_2263_43719# a_39169_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20536 a_6369_39465# a_5687_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20537 a_12079_63695# a_11797_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20538 a_3784_62607# a_3305_62607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X20539 a_19166_59142# a_18546_59184# a_19074_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2054 a_2672_39049# a_1591_38677# a_2325_38645# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X20540 vcm a_18162_63198# a_51294_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20541 a_20570_19500# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20542 VSS a_10873_36341# a_24895_35253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20543 VSS a_6424_55687# a_5955_55223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20544 a_51202_67174# pmat.row_n[11] a_51694_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20545 VSS pmat.row_n[8] a_19470_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20546 VDD a_11007_58229# a_10965_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X20547 a_23486_14878# nmat.rowon_n[9] a_23090_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20548 a_28202_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20549 VSS a_13319_35507# a_13259_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X2055 a_9195_7423# a_9020_7497# a_9374_7485# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X20550 a_7099_74313# a_9655_74216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20551 VSS a_34942_51701# a_34883_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20552 vcm a_18162_65206# a_24186_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20553 a_51598_22910# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20554 a_24094_69182# pmat.row_n[13] a_24586_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20555 a_35534_67214# pmat.rowon_n[11] a_35138_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20556 a_8669_54281# a_7479_53909# a_8560_54281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20557 vcm a_18162_9492# a_46274_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20558 a_26460_40517# a_25301_40229# a_26423_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20559 VDD a_30699_29397# a_30645_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2056 vcm a_18162_20536# a_35230_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20560 a_45270_18528# a_18546_18526# a_45178_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20561 vcm a_18162_15516# a_42258_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20562 a_5349_77071# a_4429_76751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20563 a_3423_74549# a_3267_74817# a_3568_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X20564 a_8477_49257# a_7373_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20565 a_6861_77117# a_6795_76989# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20566 a_48586_66210# pmat.rowon_n[10] a_48190_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20567 VDD a_3951_77055# a_3938_76751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20568 VDD pmat.rowoff_n[15] a_46182_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20569 VDD a_19970_46287# a_20076_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2057 VDD pmat.rowon_n[2] a_24094_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20570 a_20438_35431# a_27566_43805# a_27757_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20571 a_25190_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20572 a_18795_47491# a_16083_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20573 pmat.rowoff_n[5] a_13814_59663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20574 vcm a_18162_14512# a_46274_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20575 VDD pmat.rowoff_n[7] a_36142_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20576 a_41709_31599# a_38913_31055# a_41637_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20577 VSS a_5731_17455# a_2564_21959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20578 a_8563_7119# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20579 a_8471_73487# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2058 a_4395_46831# a_2389_45859# a_4032_46983# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X20580 a_8268_56445# a_4843_54826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20581 a_7040_8725# a_6872_8725# a_7444_9117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20582 a_47278_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20583 a_2629_31599# a_2250_31965# a_2557_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20584 VSS a_1586_8439# a_1591_8213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20585 VDD a_33007_38771# a_33033_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20586 a_40554_61190# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20587 a_2107_43401# a_1591_43029# a_2012_43389# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X20588 a_5136_19783# a_4523_21276# a_5278_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20589 vcm a_18162_16520# a_19166_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2059 VSS _1183_.A2 nmat.col[13] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X20590 VSS a_1674_68047# a_5547_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20591 a_37146_66170# a_18162_66210# a_37238_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20592 a_4588_30511# a_4471_30724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20593 a_23182_14512# a_18546_14510# a_23090_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20594 a_6817_29199# a_4068_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20595 a_23486_71230# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20596 vcm a_18162_11500# a_20170_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20597 a_37638_11468# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20598 a_30514_72234# VDD a_30118_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20599 a_37238_8488# a_18546_8486# a_37146_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 VSS a_9839_47679# a_9773_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X2060 VSS a_1586_8439# a_3063_14741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20600 vcm a_18162_10496# a_33222_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20601 a_4225_71311# a_4265_71543# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X20602 a_27198_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20603 a_44570_60186# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20604 a_44570_19898# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20605 a_27502_70226# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20606 VDD a_10651_37683# a_10677_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20607 a_20492_35529# a_20438_35431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20608 vcm a_18162_8488# a_35230_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20609 a_25098_23954# a_18162_23548# a_25190_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2061 a_24490_11866# nmat.rowon_n[12] a_24094_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20610 a_30412_31751# a_31210_31751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20611 a_23847_40183# a_22725_40229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20612 a_48282_72194# a_18546_72236# a_48190_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20613 VDD a_6699_76983# a_5047_76983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20614 VDD pmat.rowon_n[9] a_35138_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20615 a_5711_33053# a_5087_32687# a_5603_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20616 a_25691_52521# _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20617 a_46182_9898# a_18162_9492# a_46274_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20618 a_4399_51157# a_4175_49667# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X20619 a_45670_22512# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2062 pmat.col_n[27] _1194_.B1 a_45475_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X20620 a_2464_52815# a_2250_52815# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20621 a_35230_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20622 VDD pmat.rowon_n[8] a_48190_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20623 a_47764_51433# ANTENNA__1196__A2.DIODE a_47591_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20624 a_24490_63198# pmat.rowon_n[7] a_24094_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20625 VSS pmat.row_n[4] a_21478_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20626 VSS pmat.row_n[11] a_21478_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20627 VSS a_2411_43301# a_6785_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20628 VSS a_1959_10615# a_1959_10383# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X20629 VSS a_2411_16101# a_2369_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2063 a_26194_7484# a_18546_7482# a_26102_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20630 VDD a_2672_36873# a_2847_36799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20631 a_47775_52815# a_24867_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20632 a_32126_71190# a_18162_71230# a_32218_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20633 a_35630_14480# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20634 a_35534_20902# pmat.rowoff_n[12] a_35138_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20635 VSS pmat.row_n[10] a_34530_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20636 VDD pmat.rowon_n[0] a_38150_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20637 a_6895_48981# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20638 a_2012_16189# a_1895_15994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20639 a_49194_72194# VDD a_49686_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2064 VSS a_18107_53034# pmat.rowoff_n[3] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X20640 VDD a_1923_53055# a_2464_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20641 VDD nmat.rowon_n[1] a_22086_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20642 vcm a_18162_58178# a_22178_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20643 VSS a_2199_13887# a_8717_7485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20644 a_46182_14918# a_18162_14512# a_46274_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20645 a_27405_52245# a_16311_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20646 a_49686_60508# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20647 a_50290_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20648 VDD a_13909_39605# a_13853_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20649 VSS a_19584_52423# a_22522_50247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2065 a_29041_40747# a_28975_40871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20650 a_3149_40303# a_3295_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20651 vcm a_18162_57174# a_35230_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20652 a_50594_69222# pmat.rowon_n[13] a_50198_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20653 a_5658_54991# a_2791_57703# a_5578_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X20654 a_2163_69821# a_1674_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20655 VDD a_35007_44527# a_35113_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20656 a_36142_10902# pmat.row_n[2] a_36634_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20657 a_12309_36483# a_22357_35877# a_23420_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20658 a_35534_14878# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20659 VDD a_44447_45431# a_42024_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.25e+11p ps=2.85e+06u w=1e+06u l=150000u
X2066 vcm a_18162_57174# a_43262_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20660 VSS a_12447_16143# a_14441_57533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20661 a_19074_20942# pmat.row_n[12] a_19566_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20662 a_26594_72556# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20663 a_43347_52047# a_24867_53135# pmat.col[24] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20664 a_19074_16926# a_18162_16520# a_19166_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20665 VDD pmat.rowon_n[14] a_30118_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20666 VSS a_22199_30287# a_28352_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20667 a_23182_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20668 a_20078_11906# a_18162_11500# a_20170_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20669 VDD pmat.rowon_n[4] a_26102_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2067 a_44174_70186# a_18162_70226# a_44266_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20670 a_26102_62154# a_18162_62194# a_26194_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20671 a_47582_67214# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20672 a_40402_52521# ANTENNA__1184__B1.DIODE a_40099_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20673 a_30210_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20674 a_5417_11445# a_5746_11703# a_5704_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20675 VSS pmat.row_n[9] a_51598_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20676 VSS a_4703_24527# a_7479_22467# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20677 a_29477_36395# a_24833_34191# a_29391_36395# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20678 a_24873_27791# a_17139_30503# nmat.col_n[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20679 a_6829_46607# a_2935_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2068 a_43566_14878# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20680 VDD nmat.rowon_n[6] a_51202_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20681 a_19459_35279# a_19282_35279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20682 a_12311_54135# a_9581_56079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20683 VSS a_39469_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20684 a_6904_34863# a_5823_34863# a_6557_35105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X20685 a_25393_38053# a_23700_38567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X20686 VDD a_22499_49783# a_22449_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20687 a_37542_59182# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20688 VDD pmat.rowoff_n[4] a_29114_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20689 VSS _1194_.B1 a_23935_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2069 a_4124_18231# a_3305_15823# a_4266_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20690 vcm a_18162_19532# a_21174_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20691 VSS pmat.row_n[1] a_41558_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20692 VDD a_1923_69823# a_3568_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20693 VSS pmat.row_n[11] a_24490_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20694 vcm a_18162_18528# a_34226_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20695 a_48190_15922# pmat.row_n[7] a_48682_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20696 a_42258_66170# a_18546_66212# a_42166_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20697 VDD nmat.rowon_n[4] a_42166_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20698 a_2215_38671# a_1591_38677# a_2107_39049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20699 a_13345_35303# a_13653_35516# a_13319_35507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X207 a_10697_75218# a_14071_74879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2070 a_2419_69455# a_4025_54965# a_3891_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X20700 VDD pmat.rowon_n[7] a_24094_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20701 VSS a_21621_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20702 a_30687_48071# a_30999_48071# a_30957_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20703 a_25090_46831# a_25189_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20704 a_8471_73487# a_7847_73493# a_8363_73865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20705 a_31518_56170# pmat.rowon_n[0] a_31122_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20706 VDD nmat.rowon_n[5] a_28110_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20707 a_20752_39429# a_19689_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20708 a_12341_57141# a_12613_57141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X20709 a_46274_65166# a_18546_65208# a_46182_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2071 VDD a_27789_36039# a_28112_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X20710 vcm a_18162_62194# a_43262_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20711 a_46674_69544# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20712 a_11978_67279# a_11883_62063# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20713 a_43170_66170# pmat.row_n[10] a_43662_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20714 a_35752_43781# a_34593_43493# a_35656_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20715 a_15439_48071# a_15711_47899# a_15669_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20716 a_2163_61761# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20717 VDD pmat.rowon_n[11] a_50198_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20718 VSS a_2411_43301# a_2369_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20719 VDD a_2046_30184# a_9595_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2072 a_32522_59182# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20720 a_19689_42405# a_18272_42693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X20721 a_44562_45743# a_29937_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20722 VDD a_2122_17455# a_2228_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20723 a_20170_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20724 a_46182_59142# a_18162_59182# a_46274_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20725 a_5043_57399# a_4025_54965# a_5277_57533# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20726 a_50290_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20727 a_5659_38127# a_5687_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20728 a_39646_8456# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20729 a_29114_69182# a_18162_69222# a_29206_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2073 a_5705_22057# a_3305_15823# a_5633_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X20730 a_33222_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20731 a_19166_67174# a_18546_67216# a_19074_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20732 a_2397_14013# a_1687_13621# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20733 a_28456_29673# a_15667_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20734 a_50594_22910# nmat.rowon_n[1] a_50198_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20735 VDD pmat.rowon_n[13] a_23090_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20736 a_83276_12015# _1194_.B1 a_82971_11989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X20737 a_37238_17524# a_18546_17522# a_37146_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20738 a_47186_65166# pmat.row_n[9] a_47678_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20739 a_10957_14191# a_10791_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2074 a_30111_47911# a_46968_45743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X20740 a_6175_60039# a_8569_60405# a_8599_60751# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u M=2
X20741 a_23182_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20742 a_20078_56130# a_18162_56170# a_20170_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20743 VSS a_2839_38101# a_4505_40125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20744 a_47120_27247# ANTENNA__1395__A1.DIODE a_46817_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20745 a_77528_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_2.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20746 VSS a_12217_66389# a_12199_62621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20747 a_4349_62063# a_4317_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20748 a_37146_57134# pmat.row_n[1] a_37638_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20749 VDD a_39079_40947# a_39105_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X2075 VDD nmat.rowon_n[2] a_34134_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20750 a_41654_55488# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20751 a_21891_47081# a_21837_46983# a_21797_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X20752 a_47582_20902# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20753 a_21082_23954# pmat.row_n[15] a_21574_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20754 a_40349_40726# a_39469_43493# a_40532_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20755 a_21082_19938# a_18162_19532# a_21174_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20756 vcm a_18162_23548# a_42258_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20757 a_51202_12910# pmat.row_n[4] a_51694_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20758 a_24586_65528# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20759 a_2676_29941# a_2500_30345# a_2820_30333# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2076 vcm a_18162_69222# a_20170_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20760 vcm a_18162_13508# a_38242_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20761 a_9337_15033# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20762 VSS a_3325_20175# a_5547_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20763 a_42258_11500# a_18546_11498# a_42166_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20764 a_34134_22950# pmat.row_n[14] a_34626_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20765 a_35290_44527# a_35113_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20766 a_3175_59585# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20767 a_6487_5629# a_1586_8439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20768 VSS a_11261_43421# a_10953_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20769 a_24094_55126# a_18162_55166# a_24186_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2077 a_30118_16926# pmat.row_n[8] a_30610_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20770 a_37542_12870# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20771 a_18546_20534# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X20772 VDD a_7263_42453# a_7250_42845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20773 a_5626_72105# a_3866_57399# a_5323_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20774 a_10489_20291# a_4976_16091# a_10417_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20775 VSS a_11521_64239# a_11713_64899# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20776 a_44570_13874# nmat.rowon_n[10] a_44174_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20777 VSS pmat.row_n[2] a_41558_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20778 VDD config_2_in[15] a_1591_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X20779 a_27502_23914# pmat.rowoff_n[15] a_27106_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2078 VDD a_37525_27221# nmat.col_n[17] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20780 a_5233_40553# a_4831_40303# a_5069_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X20781 a_24094_14918# pmat.row_n[6] a_24586_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20782 VSS pmat.row_n[12] a_24490_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20783 a_27598_56492# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20784 VDD a_12092_42895# a_12198_42895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20785 a_9581_73487# a_9103_73791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20786 VDD a_5383_48783# a_5785_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20787 a_18546_18526# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X20788 VSS pmat.row_n[14] a_49590_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20789 a_32218_22544# a_18546_22542# a_32126_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2079 a_44729_35773# a_35244_32411# a_44647_35520# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20790 VSS pmat.row_n[0] a_20474_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20791 VDD nmat.rowon_n[15] a_24094_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20792 a_50198_18934# pmat.row_n[10] a_50690_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20793 VSS a_43720_32143# a_44927_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20794 a_47278_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20795 a_14301_27023# a_13145_26935# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20796 a_13807_72399# a_13183_72405# a_13699_72777# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20797 VDD a_10864_68565# a_10822_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20798 a_6265_37039# a_6099_37039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20799 VDD a_3659_39733# a_4031_40455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X208 a_24673_52271# a_13459_28111# pmat.col[3] VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2080 VSS a_45432_46983# a_44774_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X20800 vcm a_18162_24552# a_19166_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20801 VSS pmat.row_n[6] a_39550_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20802 a_30514_8854# nmat.rowon_n[15] a_30118_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20803 a_47147_44655# a_46896_44905# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20804 a_41254_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20805 a_43566_60186# pmat.rowon_n[4] a_43170_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20806 a_43566_19898# nmat.rowon_n[4] a_43170_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20807 VSS a_6800_44629# a_6830_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20808 VDD a_10985_35516# a_10591_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20809 VSS a_1923_69823# a_8625_73853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2081 a_24118_27791# a_17139_30503# a_23815_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X20810 a_26498_70226# pmat.rowon_n[14] a_26102_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20811 a_6412_8725# a_6956_8965# a_6914_9117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20812 a_28116_37479# a_26957_37691# a_28079_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20813 a_44266_58138# a_18546_58180# a_44174_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20814 a_22725_38053# a_20848_38341# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20815 a_22733_47381# a_22567_47381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20816 VSS a_5579_12394# a_6845_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20817 a_22086_8894# a_18162_8488# a_22178_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20818 a_30514_57174# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20819 VDD a_10515_61839# a_12907_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2082 a_47678_71552# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20820 VDD config_1_in[9] a_1591_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X20821 vcm a_18162_10496# a_41254_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20822 a_56106_40254# comp.adc_nor_latch_0.NOR_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20823 a_33386_30485# a_7415_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20824 a_12595_31433# a_12079_31061# a_12500_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X20825 a_35230_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20826 VDD VDD a_48190_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20827 VDD a_45921_42167# a_44966_43255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X20828 a_32218_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20829 a_11041_38772# a_11347_36950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2083 VSS a_33436_34191# a_33542_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20830 a_34226_69182# a_18546_69224# a_34134_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20831 a_42258_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20832 a_45270_8488# a_18546_8486# a_45178_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20833 a_14637_27247# a_11091_26311# a_14553_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20834 a_48282_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20835 a_2953_33237# a_2787_33237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20836 a_31614_19500# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20837 VDD nmat.rowon_n[13] a_35138_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20838 a_12592_18365# a_11145_17999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20839 a_46182_22950# a_18162_22544# a_46274_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2084 VDD pmat.rowoff_n[12] a_47186_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20840 a_2672_39049# a_1757_38677# a_2325_38645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20841 VDD a_1586_18231# a_1591_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X20842 VSS a_18823_50247# a_24638_49159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20843 vcm a_18162_16520# a_40250_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20844 a_43262_19532# a_18546_19530# a_43170_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20845 a_50290_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20846 comp_latch comp.adc_nor_latch_0.QN VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20847 vcm a_18162_65206# a_35230_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20848 a_11889_27907# a_10814_29111# a_11793_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20849 VSS a_10814_29111# a_11711_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2085 VDD a_16083_50069# a_16219_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20850 a_13327_70741# a_14439_72703# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20851 a_35138_69182# pmat.row_n[13] a_35630_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20852 a_46578_67214# pmat.rowon_n[11] a_46182_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20853 a_33869_31599# a_33331_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20854 a_19074_24958# a_18162_24552# a_19166_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20855 a_7131_64822# a_6451_67655# a_7131_65149# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X20856 a_23182_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20857 a_36538_59182# pmat.rowon_n[3] a_36142_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20858 a_19166_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20859 a_7073_63695# a_5081_53135# a_6639_63927# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2086 VSS pmat.row_n[4] a_19470_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20860 a_12445_58229# a_12227_58633# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20861 a_44923_32687# a_38851_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20862 VDD a_14839_20871# a_14839_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X20863 a_7258_34863# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20864 a_31210_31751# a_31217_29429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X20865 a_26957_38779# a_26276_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X20866 a_2215_20175# a_1591_20181# a_2107_20553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20867 a_2107_36873# a_1591_36501# a_2012_36861# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X20868 a_26498_24918# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20869 VDD a_36419_28023# nmat.col_n[16] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X2087 VSS a_1717_13647# a_4338_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X20870 a_32522_17890# nmat.rowon_n[6] a_32126_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20871 a_7295_62063# a_2215_47375# a_7201_62063# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X20872 VDD pmat.rowon_n[4] a_34134_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20873 VSS VDD a_37542_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20874 a_30118_55126# VDD a_30610_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20875 vcm a_18162_7484# a_24186_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20876 a_83922_9615# ANTENNA__1196__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20877 a_20170_57134# a_18546_57176# a_20078_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20878 a_22085_36374# a_21621_35515# a_22743_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20879 VSS a_25209_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X2088 a_30857_39425# a_23821_35279# a_30771_39425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20880 a_48190_66170# a_18162_66210# a_48282_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20881 a_3219_69455# a_1591_69679# a_3029_69135# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X20882 a_34226_14512# a_18546_14510# a_34134_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20883 VSS a_2199_13887# a_2157_14013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X20884 VSS pmat.row_n[6] a_20474_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20885 a_33222_56130# a_18546_56172# a_33130_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20886 a_78802_40202# a_78898_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20887 VDD a_4259_31375# a_5331_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20888 a_34226_7484# a_18546_7482# a_34134_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20889 VDD a_44763_34293# a_46811_33927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2089 VSS pmat.row_n[11] a_19470_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20890 VSS a_43720_32143# a_46027_44905# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X20891 a_29510_15882# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20892 a_34611_36649# a_33309_36039# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20893 a_14289_66421# a_13919_65871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20894 VSS pmat.row_n[5] a_33526_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20895 a_30514_10862# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20896 a_6821_18543# a_6343_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20897 a_4169_10089# a_3609_9295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20898 VDD a_25647_38695# a_18975_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X20899 nmat.rowoff_n[14] a_14839_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X209 a_45574_15882# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2090 a_21174_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20900 VDD pmat.rowon_n[15] a_24094_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20901 a_42258_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20902 vcm a_18162_70226# a_43262_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20903 VSS pmat.row_n[10] a_45574_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20904 a_27881_38341# a_28189_37981# a_12585_39355# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X20905 VSS a_19505_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X20906 VSS a_5403_67655# a_5183_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20907 VDD a_31695_43439# a_31801_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20908 a_42462_48071# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20909 VDD a_5497_62839# a_6613_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2091 a_47186_61150# a_18162_61190# a_47278_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20910 a_40158_20942# pmat.row_n[12] a_40650_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20911 a_43662_23516# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20912 a_43262_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20913 a_40158_16926# a_18162_16520# a_40250_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20914 a_21082_9898# pmat.row_n[1] a_21574_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20915 VDD pmat.rowon_n[9] a_46182_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20916 a_11969_62063# a_5651_66975# a_11883_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20917 VSS a_1923_61759# a_1881_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X20918 a_50290_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20919 a_28506_62194# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2092 a_18235_41271# a_17625_42902# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X20920 VDD a_8031_13353# a_9414_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20921 a_15065_31599# a_15021_31841# a_14899_31599# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20922 a_46274_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20923 a_31614_9460# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20924 a_30118_72194# a_18162_72234# a_30210_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20925 VSS pmat.row_n[4] a_32522_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20926 VSS pmat.row_n[11] a_32522_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20927 a_22482_66210# pmat.rowon_n[10] a_22086_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20928 VDD pmat.rowon_n[1] a_36142_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20929 a_9557_17705# a_9155_17455# a_9393_17455# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X2093 a_26331_44535# a_25209_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X20930 a_46674_14480# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20931 VDD nmat.rowon_n[6] a_49194_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20932 a_46578_20902# pmat.rowoff_n[12] a_46182_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20933 VDD pmat.rowoff_n[15] a_20078_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20934 VSS a_44733_44431# a_45003_43343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20935 a_12488_36367# a_12237_36596# a_12267_36694# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X20936 a_2563_34837# a_2847_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20937 a_44174_15922# a_18162_15516# a_44266_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20938 VDD pmat.rowoff_n[4] a_50198_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20939 a_4901_30753# a_4683_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2094 a_20170_12504# a_18546_12502# a_20078_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20940 a_22963_42657# a_10781_42869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20941 a_29606_24520# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20942 a_20078_64162# a_18162_64202# a_20170_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20943 a_9643_66389# a_10921_64786# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20944 a_19166_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20945 VDD nmat.rowon_n[1] a_33130_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20946 vcm a_18162_58178# a_33222_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20947 a_36538_12870# pmat.rowoff_n[4] a_36142_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20948 a_12587_30838# a_6927_30503# a_12128_30663# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20949 a_19470_64202# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2095 a_23582_9460# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20950 VDD a_45119_32661# a_44923_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20951 a_44183_27497# a_18243_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20952 VDD nmat.rowon_n[9] a_23090_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20953 vcm a_18162_21540# a_38242_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20954 a_47186_10902# pmat.row_n[2] a_47678_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20955 a_21174_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20956 a_41254_61150# a_18546_61192# a_41162_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20957 VDD pmat.rowon_n[12] a_44174_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20958 a_24094_63158# a_18162_63198# a_24186_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20959 a_45574_68218# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2096 VDD pmat.rowoff_n[4] a_37146_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20960 a_3399_24787# a_3325_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X20961 a_34226_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20962 a_10591_35561# a_10985_35516# a_10651_35507# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X20963 VSS a_2529_44409# a_2463_44477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20964 a_29510_56170# pmat.rowon_n[0] a_29114_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20965 VSS a_4720_58487# a_4719_58255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20966 VDD nmat.rowon_n[10] a_27106_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20967 a_24586_10464# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20968 VDD a_31425_37218# a_30489_36893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X20969 a_46108_32687# a_43776_30287# a_45805_32661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2097 a_11116_18695# a_5351_19913# a_11258_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20970 a_2080_72221# a_1643_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20971 a_45270_60146# a_18546_60188# a_45178_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20972 VDD a_3613_19061# a_3503_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20973 VSS pmat.row_n[12] a_22482_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20974 a_45670_64524# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20975 a_48586_59182# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20976 a_42166_61150# pmat.row_n[5] a_42658_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20977 VDD a_5320_30199# a_4951_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20978 vcm a_18162_19532# a_32218_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20979 VDD a_3838_70455# a_3795_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2098 a_16966_29423# a_12437_28879# a_16966_29673# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X20980 a_50198_69182# a_18162_69222# a_50290_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20981 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20982 a_8086_52093# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20983 a_31518_18894# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20984 a_4070_47375# a_3799_47375# a_3987_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X20985 a_43659_28853# a_43451_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20986 a_35630_56492# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20987 a_36380_34191# a_36203_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20988 a_37238_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20989 a_7999_31359# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2099 vcm a_18162_68218# a_24186_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20990 a_11752_52931# a_10641_52815# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20991 a_40250_22544# a_18546_22542# a_40158_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20992 a_15259_31029# clk_ena a_15690_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X20993 a_29931_30517# a_23021_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20994 a_47321_37289# a_30571_50959# a_47035_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20995 a_4491_53511# a_4243_54991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20996 a_38972_39655# a_37813_39867# a_38935_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20997 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20998 VDD pmat.rowon_n[8] a_22086_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20999 a_36234_12504# a_18546_12502# a_36142_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u M=1806
X210 VSS pmat.row_n[10] a_48586_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2100 a_35230_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21000 a_46182_60146# pmat.row_n[4] a_46674_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21001 VDD VDD a_38150_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21002 a_50198_7890# VDD a_50690_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21003 VDD a_4220_62037# a_2944_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21004 a_19689_35877# a_18272_35077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21005 a_13158_71285# a_8491_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21006 a_4031_37191# a_3325_36495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21007 VSS a_10423_64786# a_10707_64783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21008 VDD a_3615_71631# a_14749_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21009 VSS a_13329_47893# a_12328_48168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2101 VDD a_20879_47893# a_12447_16143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X21010 a_4432_42313# a_4149_41941# a_4337_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21011 a_26102_7890# VDD a_26594_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21012 a_34530_70226# pmat.rowon_n[14] a_34134_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21013 a_20267_50345# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21014 a_19074_62154# pmat.row_n[6] a_19566_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21015 VSS pmat.row_n[2] a_29510_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21016 a_23582_60508# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21017 VDD a_2325_8181# a_2215_8207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21018 a_31214_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21019 a_32522_7850# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2102 a_82815_54965# ANTENNA_fanout52_A.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21020 a_38150_21946# a_18162_21540# a_38242_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21021 VSS a_4075_31591# a_14816_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21022 a_2319_74268# a_2124_74299# a_2629_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X21023 VDD a_19417_43990# a_20752_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X21024 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X21025 a_13553_50461# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21026 a_23663_36649# a_23700_36391# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21027 a_24719_37429# a_24895_37429# a_24847_37455# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21028 a_37542_61190# pmat.rowon_n[5] a_37146_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21029 VSS a_11019_71543# a_11204_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2103 clk_comp a_40399_36911# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X21030 a_14833_28585# a_14645_28381# a_14751_28341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21031 a_21478_67214# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21032 a_34226_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21033 a_51598_56170# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21034 VSS VDD a_48586_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21035 a_45574_21906# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21036 vcm a_18162_24552# a_40250_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21037 a_39015_47375# a_38391_47381# a_38907_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21038 a_34530_66210# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21039 a_48190_57134# pmat.row_n[1] a_48682_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2104 VDD a_6612_15797# a_1586_8439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21040 a_38242_59142# a_18546_59184# a_38150_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21041 a_23043_28335# a_22792_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21042 a_32126_23954# pmat.row_n[15] a_32618_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21043 a_32126_19938# a_18162_19532# a_32218_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21044 VSS a_10873_38517# a_22963_35041# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21045 a_20752_38341# a_19689_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21046 VSS pmat.row_n[8] a_38546_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21047 a_9602_10749# a_2021_11043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21048 VSS a_25647_37607# a_21219_36885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X21049 VDD a_1923_61759# a_2464_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2105 a_2244_20871# config_1_in[12] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21050 a_42562_14878# nmat.rowon_n[9] a_42166_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21051 VDD a_1586_18231# a_9411_15831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X21052 a_36234_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21053 a_35138_55126# a_18162_55166# a_35230_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21054 VDD a_12715_51420# a_12646_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21055 a_22086_15922# pmat.row_n[7] a_22578_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21056 a_48586_12870# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21057 a_1979_9661# a_1725_9334# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21058 a_25590_18496# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21059 a_25494_24918# VSS a_25098_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2106 VSS a_7999_31359# a_7933_31433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X21060 VSS pmat.row_n[13] a_22482_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21061 VDD a_5156_28335# a_5331_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21062 a_19166_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21063 a_4165_67503# a_2791_57703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21064 a_33412_52271# ANTENNA__1395__A1.DIODE a_33109_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21065 a_1644_59861# a_1591_58799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21066 vcm a_18162_55166# a_39246_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21067 VSS a_27913_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21068 a_35138_14918# pmat.row_n[6] a_35630_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21069 VSS a_14528_48114# a_14486_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2107 a_43561_47893# a_30111_47911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21070 a_39154_59142# pmat.row_n[3] a_39646_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21071 a_2250_52815# a_2163_53057# a_1846_52947# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21072 VSS a_19233_41479# a_20075_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21073 VDD _1179_.X a_83362_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X21074 a_10498_19631# a_10151_19637# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X21075 a_28506_15882# pmat.rowoff_n[7] a_28110_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21076 a_4031_32852# a_4123_32661# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X21077 VSS pmat.row_n[7] a_37542_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21078 a_11133_44581# a_10651_44211# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X21079 a_20170_65166# a_18546_65208# a_20078_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2108 a_4956_59317# a_2879_57487# a_5179_59663# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X21080 a_20570_69544# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21081 a_14462_61839# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21082 a_5197_16121# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X21083 a_10423_16055# a_10167_16950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21084 vcm a_18162_66210# a_29206_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21085 a_33222_64162# a_18546_64204# a_33130_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21086 vcm a_18162_61190# a_30210_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21087 a_47731_36103# a_47207_35951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21088 VDD a_2972_9991# a_4003_7663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21089 a_21174_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2109 VDD ANTENNA__1395__A1.DIODE a_83007_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X21090 VDD a_30278_30511# a_33299_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21091 a_33622_68540# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21092 a_29606_58500# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21093 a_6794_64015# a_4985_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21094 a_25688_32117# a_11067_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21095 VSS pmat.row_n[3] a_29510_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21096 a_35036_32375# a_35244_32411# a_35178_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21097 a_42258_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21098 a_21082_65166# pmat.row_n[9] a_21574_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21099 a_12053_27497# a_11235_26159# a_11969_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X211 VSS a_6283_31591# a_22567_47381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2110 a_25209_36965# a_22059_37683# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X21100 a_4801_69929# a_4991_69831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21101 a_42562_71230# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21102 vcm a_18162_60186# a_34226_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21103 a_34134_64162# pmat.row_n[8] a_34626_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21104 a_40158_24958# a_18162_24552# a_40250_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21105 a_39646_21508# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21106 VSS a_15259_31029# a_5535_29980# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21107 a_39246_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21108 a_25190_9492# a_18546_9490# a_25098_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21109 VSS a_33765_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X2111 VSS a_4032_46983# a_3793_47479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21110 a_8673_7093# a_8455_7497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21111 a_4583_18038# a_3305_15823# a_4124_18231# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21112 a_21478_20902# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21113 a_46274_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21114 VSS a_4048_74549# a_3986_74575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X21115 a_43170_60146# a_18162_60186# a_43262_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21116 VSS a_1923_31743# a_10373_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21117 a_24094_56130# pmat.row_n[0] a_24586_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21118 VDD a_23329_37462# a_22393_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X21119 a_2215_27791# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2112 VDD nmat.rowon_n[14] a_33130_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21120 VDD a_6608_60663# a_5053_59575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21121 VSS a_1586_18231# a_2603_22357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21122 a_13361_68841# a_13173_68597# a_13279_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21123 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X21124 a_3325_26159# a_2847_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21125 a_46578_70226# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21126 a_3116_77117# a_2999_76922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21127 a_28202_15516# a_18546_15514# a_28110_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21128 vcm a_18162_12504# a_25190_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21129 VSS a_9441_20189# a_12353_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2113 a_12999_3855# _1194_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X21130 a_44174_23954# a_18162_23548# a_44266_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21131 a_14399_12879# a_10239_14183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X21132 a_6339_40303# a_5989_40303# a_6244_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21133 VDD nmat.rowon_n[13] a_46182_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21134 a_24197_42405# a_23741_42567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X21135 a_15107_40183# a_13985_40229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21136 a_19166_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21137 a_36538_62194# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21138 VSS pmat.row_n[4] a_40554_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21139 VSS pmat.row_n[11] a_40554_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2114 vcm a_18162_18528# a_42258_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21140 a_10239_20291# a_4523_21276# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21141 a_19470_72234# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21142 VSS pmat.row_n[14] a_23486_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21143 a_49590_61190# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21144 VSS a_10878_58487# a_11149_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X21145 VSS a_19487_53034# pmat.rowoff_n[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21146 a_51202_71190# a_18162_71230# a_51294_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21147 a_13909_67279# a_13432_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21148 vcm a_18162_71230# a_37238_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21149 a_3399_62607# a_3345_62839# a_3305_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X2115 a_24895_39605# a_12116_39783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21150 a_50594_15882# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21151 VDD a_45432_46983# a_44774_48695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X21152 a_5633_46831# a_5221_45199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21153 VSS a_30999_48071# a_30947_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21154 vcm a_18162_11500# a_29206_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21155 a_21174_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21156 a_13801_34427# a_12568_35077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21157 VDD comp.adc_nor_latch_0.QN a_55418_40254# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21158 a_1644_58229# a_1823_58237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21159 vcm a_18162_58178# a_41254_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2116 a_8697_57167# a_4128_64391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X21160 VDD comp.adc_comp_circuit_0.adc_comp_buffer_0.in a_54790_39936# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X21161 a_22725_40229# a_22269_40391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21162 a_37638_63520# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21163 a_7129_57685# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21164 VDD config_1_in[8] a_1591_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X21165 a_34226_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21166 VDD pmat.rowon_n[5] a_41162_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21167 a_6917_27907# a_4516_21531# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21168 VDD a_6467_29415# a_7939_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21169 a_38935_39913# a_37813_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2117 a_48282_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21170 VSS pmat.row_n[5] a_26498_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21171 a_23486_17890# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21172 VSS a_6927_30503# a_11004_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21173 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X21174 a_30514_18894# nmat.rowon_n[5] a_30118_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21175 a_4061_63303# a_3784_62607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21176 a_20393_41046# a_20221_40835# a_20179_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X21177 VDD a_4032_46983# a_3793_47479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21178 a_11634_48285# a_11508_48187# a_11230_48171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X21179 nmat.rowoff_n[3] a_13551_8751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2118 a_41573_51701# a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X21180 nmat.col[14] a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21181 VSS a_19405_28853# a_30699_29397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21182 a_45670_72556# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21183 vcm a_18162_69222# a_31214_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21184 VDD a_13319_35507# a_13345_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X21185 VDD pmat.rowon_n[4] a_45178_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21186 vcm a_18162_59182# a_27198_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21187 a_8455_7497# a_7939_7125# a_8360_7485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21188 a_19487_53034# a_19579_52789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21189 a_31214_57134# a_18546_57176# a_31122_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2119 a_38095_32143# a_2007_25597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X21190 a_27502_16886# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21191 a_41795_30511# a_41321_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21192 a_25190_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21193 a_21279_48999# a_44870_48437# a_44806_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21194 VSS pmat.row_n[6] a_31518_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21195 a_25098_10902# a_18162_10496# a_25190_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21196 a_25287_32117# clk_ena VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21197 VDD VDD a_22086_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21198 a_36234_20536# a_18546_20534# a_36142_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21199 VDD a_1923_61759# a_3476_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X212 VSS a_31095_42367# a_31041_42689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2120 a_24186_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21200 VSS a_2046_30184# a_19439_32149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21201 a_48586_9858# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21202 a_39550_69222# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21203 a_12227_12937# a_11877_12565# a_12132_12925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21204 VSS pmat.row_n[11] a_43566_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21205 a_40554_64202# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21206 VDD a_1828_25589# a_1858_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21207 VDD a_4955_40277# a_4831_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21208 a_9601_51005# a_9427_50095# a_9529_51005# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21209 a_18973_29199# a_8583_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.1295e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2121 a_48586_69222# pmat.rowon_n[13] a_48190_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21210 VSS a_6559_33767# a_9963_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21211 a_22811_32521# a_22365_32149# a_22715_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21212 a_5123_52423# a_2389_45859# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21213 a_19074_70186# pmat.row_n[14] a_19566_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21214 VSS a_1591_14735# a_1769_14735# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X21215 a_46934_35951# a_30571_50959# a_46765_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21216 a_14803_31599# a_14287_31599# a_14708_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21217 a_17113_42405# a_16657_42567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21218 a_20474_67214# pmat.rowon_n[11] a_20078_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21219 a_29114_11906# a_18162_11500# a_29206_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2122 VDD a_5462_62215# a_5553_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X21220 a_30210_18528# a_18546_18526# a_30118_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21221 a_50594_56170# pmat.rowon_n[0] a_50198_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21222 VDD nmat.rowon_n[5] a_47186_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21223 a_14174_51859# a_14491_51969# a_14449_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21224 a_44666_15484# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21225 a_7352_65149# a_5307_67655# a_7131_64822# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21226 VSS a_9983_32385# a_9944_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21227 a_8025_24233# a_4703_24527# a_7929_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21228 a_6553_53047# a_6787_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21229 a_33526_66210# pmat.rowon_n[10] a_33130_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2123 a_41558_17890# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21230 VDD pmat.rowoff_n[15] a_31122_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21231 a_5225_34685# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21232 VDD a_9552_67191# a_8819_67197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X21233 VSS a_3576_17143# a_5463_17027# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21234 a_35534_9858# nmat.rowon_n[14] a_35138_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21235 VDD a_2672_64073# a_2847_63999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21236 a_9668_10651# a_9655_6335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21237 a_6557_40545# a_6339_40303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21238 VSS a_13909_39605# a_17811_39605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21239 a_2012_43389# a_1895_43194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2124 a_4043_59861# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X21240 a_46936_44111# a_43720_32143# a_46763_44431# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21241 vcm a_18162_14512# a_31214_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21242 VDD pmat.rowoff_n[7] a_21082_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21243 a_38242_67174# a_18546_67216# a_38150_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21244 a_45178_11906# pmat.row_n[3] a_45670_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21245 VDD a_33839_46805# a_40047_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21246 comp.adc_inverter_1.in clk_comp VDD VDD sky130_fd_pr__pfet_01v8 ad=2.394e+11p pd=2.82e+06u as=0p ps=0u w=420000u l=150000u M=2
X21247 VDD pmat.rowon_n[13] a_42166_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21248 a_28110_21946# pmat.row_n[13] a_28602_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21249 a_28110_17930# a_18162_17524# a_28202_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2125 VDD a_14653_53458# a_19595_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21250 VDD pmat.rowon_n[3] a_38150_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21251 a_32218_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21252 a_39209_29423# a_37827_30793# a_39127_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21253 VDD nmat.rowon_n[7] nmat.rowoff_n[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X21254 a_12705_10389# a_12539_10389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21255 VSS pmat.row_n[1] a_33526_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21256 a_35138_63158# a_18162_63198# a_35230_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21257 a_25190_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21258 a_22086_66170# a_18162_66210# a_22178_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21259 a_27502_57174# pmat.rowon_n[1] a_27106_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2126 a_25190_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21260 pmat.col_n[20] ANTENNA__1184__B1.DIODE a_39301_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21261 a_2080_65693# a_1643_65301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21262 a_22578_11468# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21263 vcm a_18162_63198# a_39246_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21264 a_7176_8751# a_7040_8725# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21265 a_44174_7890# a_18162_7484# a_44266_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21266 a_39154_67174# pmat.row_n[11] a_39646_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21267 a_43662_65528# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21268 a_40158_62154# pmat.row_n[6] a_40650_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21269 a_14289_59049# a_10515_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2127 a_12003_52815# a_11752_52931# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X21270 a_10969_71631# a_11115_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21271 a_19413_40229# a_17996_40743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21272 a_12196_44869# a_11133_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21273 a_12449_23145# a_5899_21807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21274 a_39550_22910# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21275 VDD a_22499_49783# a_37471_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21276 a_10898_77661# a_10811_77437# a_10494_77547# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21277 VSS pmat.row_n[12] a_43566_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21278 VDD a_4031_20884# a_3183_19258# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X21279 a_33222_72194# a_18546_72236# a_33130_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2128 a_22086_21946# a_18162_21540# a_22178_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21280 a_46674_56492# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21281 VDD pmat.rowon_n[9] a_20078_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21282 a_26102_24958# VDD a_26594_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21283 a_29206_62154# a_18546_62196# a_29114_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21284 a_41558_71230# pmat.rowon_n[15] a_41162_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21285 a_30610_22512# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21286 a_30118_8894# pmat.row_n[0] a_30610_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21287 a_29606_66532# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21288 a_51294_22544# a_18546_22542# a_51202_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21289 a_12757_39126# a_12585_39355# a_12543_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2129 VDD pmat.rowon_n[14] a_28110_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21290 a_20170_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21291 VSS a_17113_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21292 VDD pmat.rowon_n[8] a_33130_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21293 a_47278_12504# a_18546_12502# a_47186_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21294 VDD a_79085_40202# a_78898_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21295 a_4081_76457# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X21296 a_29676_40517# a_28613_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21297 a_29114_56130# a_18162_56170# a_29206_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21298 VDD a_19049_41959# a_17154_43671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21299 VDD a_5779_13255# a_5131_13255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X213 ANTENNA__1197__B.DIODE a_25695_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=0p ps=0u w=650000u l=150000u M=8
X2130 VDD nmat.sample_n a_18162_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X21300 a_20570_14480# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21301 a_20474_20902# pmat.rowoff_n[12] a_20078_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21302 VSS a_32305_51335# a_31631_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21303 VDD pmat.rowon_n[0] a_23090_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21304 a_14657_46403# nmat.sw a_14562_46403# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21305 VSS a_28915_50959# a_32871_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21306 a_34134_72194# VDD a_34626_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21307 a_45574_70226# pmat.rowon_n[14] a_45178_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21308 a_31122_14918# a_18162_14512# a_31214_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21309 a_34626_60508# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2131 VDD nmat.rowon_n[5] a_36142_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21310 a_14328_39631# a_12969_40175# a_14107_39958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X21311 VDD a_6087_67655# a_4396_66933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X21312 a_35534_62194# pmat.rowon_n[6] a_35138_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21313 a_21082_10902# pmat.row_n[2] a_21574_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21314 VDD a_2163_65469# a_2124_65595# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X21315 VDD VSS a_27106_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21316 nmat.col_n[10] a_14458_5487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21317 VDD a_2847_23743# a_2834_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21318 vcm a_18162_20536# a_25190_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21319 a_28202_23548# a_18546_23546# a_28110_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2132 a_8577_18115# a_8305_20871# a_8481_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21320 VSS a_2952_25045# a_6747_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21321 a_48586_61190# pmat.rowon_n[5] a_48190_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21322 VSS a_31210_31751# a_31479_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21323 a_32522_67214# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21324 VDD a_1923_31743# a_2464_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21325 a_6720_49007# a_5805_49007# a_6373_49249# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21326 a_39246_8488# a_18546_8486# a_39154_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21327 a_5423_67191# a_2419_53351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21328 a_4903_64015# a_4351_55527# a_4809_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21329 VSS a_4128_46983# a_5747_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2133 a_12266_48285# a_11508_48187# a_11703_48156# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X21330 vcm a_18162_66210# a_50290_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21331 a_27502_10862# nmat.rowon_n[13] a_27106_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21332 VSS a_18823_50247# a_21970_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21333 a_2417_45173# a_2199_45577# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21334 a_49286_59142# a_18546_59184# a_49194_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21335 a_1953_5059# a_1761_6031# a_1857_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21336 VDD a_2419_53351# a_4162_64561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21337 a_50690_19500# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21338 a_5455_22057# a_3351_27249# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21339 VSS a_17336_43439# a_17442_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2134 VSS a_3956_72373# a_3894_72399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X21340 a_22482_59182# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21341 a_4071_47919# a_4075_50087# a_4071_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21342 VSS pmat.row_n[8] a_49590_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21343 a_20078_16926# pmat.row_n[8] a_20570_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21344 a_47278_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21345 a_37638_71552# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21346 VDD a_9305_58229# a_5535_57993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X21347 a_2944_56872# a_3514_57167# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X21348 VDD pmat.rowoff_n[12] a_37146_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21349 a_28112_35303# a_27049_35515# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2135 VSS a_23823_47679# a_15899_47939# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X21350 a_3871_6031# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21351 a_33130_15922# pmat.row_n[7] a_33622_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21352 a_4450_24310# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X21353 a_37146_61150# a_18162_61190# a_37238_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21354 a_2834_43023# a_1757_43029# a_2672_43401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21355 a_12981_74581# a_12815_74581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21356 VSS a_16890_36911# a_18999_35279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21357 VSS a_4075_31591# a_14816_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21358 VSS a_27421_41814# a_27895_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21359 a_26498_58178# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2136 a_50594_72234# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21360 VSS a_20787_30199# a_20591_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X21361 a_26498_16886# nmat.rowon_n[7] a_26102_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21362 VDD a_9655_6335# a_9642_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21363 a_5462_30333# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21364 a_8695_12801# a_3571_13627# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21365 vcm a_18162_67214# a_27198_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21366 a_38242_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21367 a_38546_69222# pmat.rowon_n[13] a_38150_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21368 a_31214_65166# a_18546_65208# a_31122_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21369 a_31614_69544# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2137 VDD a_7436_60039# a_6816_60699# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21370 a_27198_55126# a_18546_55168# a_27106_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21371 vcm a_18162_17524# a_45270_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21372 a_2425_36201# a_1899_35051# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X21373 a_27598_59504# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21374 VSS a_5565_19605# a_5499_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21375 a_28626_29423# a_28812_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21376 a_31122_59142# a_18162_59182# a_31214_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21377 VSS a_15667_27239# a_45923_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21378 VDD a_35382_34191# a_36203_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21379 a_40554_72234# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2138 a_28202_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21380 VSS pmat.row_n[9] a_39550_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21381 VSS a_37820_30485# a_41593_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21382 a_22178_17524# a_18546_17522# a_22086_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21383 vcm a_18162_16520# a_49286_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21384 a_32126_65166# pmat.row_n[9] a_32618_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21385 a_7645_53909# a_7479_53909# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21386 a_6981_28879# a_4068_25615# a_6909_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21387 vcm a_18162_11500# a_50290_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21388 a_37238_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21389 a_10057_67753# a_5363_70543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2139 a_12489_58621# a_12445_58229# a_12323_58633# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X21390 a_45645_45895# a_31675_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21391 a_4036_70741# a_4421_70741# a_4165_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X21392 VSS a_14379_46287# a_14486_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21393 a_46427_39009# a_40837_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21394 VSS a_2199_13887# a_3105_11837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21395 nmat.col_n[13] a_14734_4175# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21396 VSS a_2411_33749# a_4549_34685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21397 a_22086_57134# pmat.row_n[1] a_22578_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21398 a_32522_20902# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21399 VSS a_2659_35015# a_2509_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X214 a_10791_26409# a_9579_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X2140 VSS pmat.row_n[9] a_49590_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21400 VSS a_13985_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21401 VDD pmat.rowon_n[5] a_39154_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21402 a_35138_56130# pmat.row_n[0] a_35630_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21403 a_26194_16520# a_18546_16518# a_26102_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21404 a_44266_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21405 vcm a_18162_13508# a_23182_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21406 VSS _1196_.B1 a_32305_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21407 a_6060_49007# a_5785_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21408 a_41784_52271# a_11067_27239# a_41481_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21409 VSS pmat.row_n[7] a_25494_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2141 a_32218_17524# a_18546_17522# a_32126_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21410 a_22482_12870# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21411 VSS a_24719_43957# a_14773_43746# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21412 a_6757_75663# a_6051_74183# a_5497_73719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21413 a_2104_45565# a_1987_45370# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X21414 a_47582_62194# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21415 a_13519_55369# a_13073_54997# a_13423_55369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21416 VSS pmat.row_n[4] a_51598_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21417 VSS pmat.row_n[11] a_51598_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21418 VDD a_12053_27497# a_22874_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21419 a_5081_13103# a_5227_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2142 a_39469_43493# a_39013_43655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21420 VSS pmat.row_n[14] a_34530_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21421 a_26102_58138# pmat.row_n[2] a_26594_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21422 a_4313_44111# a_3911_44431# a_4149_44431# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X21423 a_33033_37479# a_33341_37692# a_33007_37683# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21424 vcm a_18162_71230# a_48282_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21425 VDD pmat.rowon_n[11] a_38150_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21426 VDD a_18975_40871# a_20393_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21427 a_26498_11866# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21428 a_32218_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21429 VSS a_2319_72092# a_2250_72221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2143 a_22199_30287# a_41731_49525# a_46395_29199# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X21430 VDD a_2847_50069# a_2834_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21431 a_48682_24520# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21432 a_38242_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21433 VSS a_11067_30287# a_40966_46653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21434 VDD a_3496_51701# a_3434_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21435 a_7578_48553# a_8091_49192# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=0p ps=0u w=650000u l=150000u
X21436 VSS pmat.row_n[6] a_24490_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21437 a_47035_43817# a_7109_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21438 VSS a_29036_41831# a_28999_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21439 a_16552_46805# a_16403_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2144 pmat.rowoff_n[7] a_14340_19783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X21440 VDD a_4025_54965# a_6583_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21441 a_38546_22910# nmat.rowon_n[1] a_38150_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21442 a_37542_8854# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21443 a_36142_21946# pmat.row_n[13] a_36634_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21444 VSS a_1591_74031# a_1985_76001# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21445 VDD nmat.rowon_n[9] a_42166_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21446 a_36142_17930# a_18162_17524# a_36234_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21447 a_40158_70186# pmat.row_n[14] a_40650_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21448 VDD a_39413_40956# a_39019_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21449 a_40250_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2145 VDD nmat.rowon_n[15] a_49194_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21450 a_17503_32143# a_10055_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21451 a_8941_22467# a_5899_21807# a_8859_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21452 VDD VSS a_25098_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21453 VDD a_3663_9269# a_3609_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21454 VDD a_10781_42364# a_10725_42390# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X21455 a_49194_20942# pmat.row_n[12] a_49686_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21456 a_49194_16926# a_18162_16520# a_49286_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21457 VSS pmat.row_n[0] a_47582_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21458 a_50198_11906# a_18162_11500# a_50290_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21459 VDD a_4383_7093# a_10741_17782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2146 VSS pmat.row_n[0] a_45574_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21460 VSS a_34277_38550# a_33341_38780# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X21461 VDD a_15049_36374# a_14113_36604# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X21462 a_39154_12910# pmat.row_n[4] a_39646_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21463 a_43662_10464# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21464 a_29206_70186# a_18546_70228# a_29114_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21465 VDD pmat.rowoff_n[15] a_29114_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21466 a_47947_27247# ANTENNA__1195__A1.DIODE nmat.col_n[27] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21467 a_20170_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21468 a_26594_20504# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21469 VDD VDD a_33130_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2147 VDD a_15049_42902# a_14113_43132# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X21470 VSS pmat.row_n[12] a_41558_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21471 a_26194_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21472 a_47278_20536# a_18546_20534# a_47186_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21473 vcm a_18162_19532# a_51294_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21474 a_33227_52047# ANTENNA__1195__A1.DIODE pmat.col_n[13] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21475 a_29114_64162# a_18162_64202# a_29206_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21476 a_33222_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21477 a_9651_62985# a_9301_62613# a_9556_62973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21478 a_40650_8456# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21479 a_40129_29423# a_38905_28853# a_39496_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2148 VDD a_3061_11445# a_2951_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X21480 VDD pmat.rowoff_n[7] a_19074_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21481 VSS a_23933_32143# a_25423_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21482 a_17113_35877# a_13503_36893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21483 VDD a_1586_18231# a_1591_23445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X21484 a_12585_37179# a_17113_35877# a_18176_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X21485 VDD nmat.rowon_n[13] a_20078_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21486 VDD a_7779_22583# a_9385_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21487 VSS a_2046_30184# a_5087_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21488 a_31122_22950# a_18162_22544# a_31214_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21489 VSS a_11271_73085# a_11232_73211# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2149 a_82736_4943# ANTENNA__1190__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X21490 VSS pmat.row_n[3] a_44570_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21491 VDD nmat.rowon_n[15] a_50198_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21492 a_38150_18934# pmat.row_n[10] a_38642_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21493 a_27106_12910# a_18162_12504# a_27198_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21494 a_11910_47197# a_11823_46973# a_11506_47083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21495 a_42658_16488# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21496 VSS pmat.row_n[13] a_27502_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21497 a_44783_45743# a_44635_46025# a_44420_45895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21498 a_6933_77117# a_6799_75637# a_6861_77117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21499 a_31518_67214# pmat.rowon_n[11] a_31122_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X215 a_6283_31591# a_7387_33231# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X2150 a_47278_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21500 a_10613_8573# a_10047_8751# a_10541_8573# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21501 a_31412_43439# a_31235_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21502 VDD a_12263_50959# a_16403_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21503 a_3061_11445# a_2843_11849# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21504 a_32522_8854# nmat.rowon_n[15] a_32126_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21505 a_10693_25321# a_9528_20407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21506 a_21478_59182# pmat.rowon_n[3] a_21082_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21507 VSS pmat.row_n[2] a_48586_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21508 a_45574_55166# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21509 a_1644_77813# a_1823_77821# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2151 VSS a_10139_32117# a_10070_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X21510 a_50290_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21511 a_6009_74281# a_5931_74183# a_4601_74005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21512 a_36234_68178# a_18546_68220# a_36142_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21513 a_28506_65206# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21514 VDD a_1591_16367# a_1739_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21515 a_7213_19407# a_4976_16091# a_7131_19407# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21516 a_9869_62581# a_9651_62985# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21517 VDD a_4328_6409# a_4503_6335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21518 a_49286_67174# a_18546_67216# a_49194_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21519 a_18546_66212# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X2152 VDD a_4613_19087# a_5179_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21520 VSS a_2199_13887# a_9177_6397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21521 a_2559_44150# a_1739_47893# a_2100_44343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21522 a_5357_62779# a_6583_61519# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21523 a_4588_30511# a_4471_30724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21524 a_39550_71230# pmat.rowon_n[15] a_39154_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21525 a_20078_67174# a_18162_67214# a_20170_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21526 a_25494_58178# pmat.rowon_n[2] a_25098_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21527 VSS VDD a_22482_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21528 a_21621_35515# a_20848_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X21529 a_50198_56130# a_18162_56170# a_50290_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2153 a_22325_36950# a_22153_37179# a_22111_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X21530 a_22787_34165# a_11317_36924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21531 a_28602_61512# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21532 a_24094_8894# a_18162_8488# a_24186_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21533 a_33130_66170# a_18162_66210# a_33222_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21534 VSS a_33845_27765# nmat.col_n[14] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21535 VDD comp_latch a_10443_12879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21536 VSS a_44420_45895# a_41926_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21537 a_19566_19500# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21538 VSS a_4383_7093# a_10741_17782# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21539 a_22377_51727# ANTENNA__1196__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2154 a_26102_20942# a_18162_20536# a_26194_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21540 a_51202_23954# pmat.row_n[15] a_51694_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21541 a_28971_47753# a_28621_47381# a_28876_47741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21542 a_51202_19938# a_18162_19532# a_51294_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21543 a_34226_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21544 a_6612_66933# a_2407_49289# a_6832_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21545 a_26671_46831# a_26321_46831# a_26576_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21546 a_37542_23914# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21547 a_36324_46983# a_36532_46805# a_36466_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21548 a_44570_24918# VSS a_44174_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21549 a_41162_15922# pmat.row_n[7] a_41654_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2155 a_2672_20553# a_1757_20181# a_2325_20149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X21550 VSS pmat.row_n[13] a_41558_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21551 a_20329_35431# a_20534_35431# a_20492_35529# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21552 a_38242_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21553 VSS pmat.row_n[10] a_30514_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21554 a_44666_57496# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21555 VSS a_17113_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21556 a_11149_59887# a_11007_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21557 a_27198_63158# a_18546_63200# a_27106_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21558 a_22085_37479# a_22393_37692# a_22059_37683# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21559 a_27598_67536# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2156 VSS a_37823_34191# nmat.sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X21560 a_9731_9839# a_9583_10121# a_9368_9991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X21561 VSS a_21239_47349# a_18547_51565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X21562 VDD pmat.rowon_n[9] a_31122_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21563 a_34530_16886# nmat.rowon_n[7] a_34134_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21564 a_45563_31055# a_45019_38645# a_45345_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21565 a_27106_57134# a_18162_57174# a_27198_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21566 VDD a_2411_33749# a_9231_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21567 a_14833_29967# a_12851_28853# a_14465_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21568 a_31214_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21569 VDD a_5211_57172# a_5043_57399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2157 a_12542_47197# a_11823_46973# a_11979_47068# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X21570 a_47582_15882# pmat.rowoff_n[7] a_47186_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21571 VSS pmat.row_n[4] a_44570_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21572 a_10325_69679# a_9135_69679# a_10216_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X21573 a_25226_28335# a_8583_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21574 VDD pmat.rowon_n[1] a_21082_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21575 VSS pmat.row_n[14] a_27502_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21576 a_35230_55126# a_18546_55168# a_35138_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21577 a_31614_14480# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21578 a_31518_20902# pmat.rowoff_n[12] a_31122_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21579 vcm a_18162_24552# a_49286_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2158 vcm a_18162_19532# a_19166_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21580 a_10378_70045# a_9301_69679# a_10216_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21581 a_35630_59504# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21582 VDD a_5331_53511# a_4081_61127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X21583 a_9361_47741# a_9317_47349# a_9195_47753# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21584 VSS a_1586_33927# a_1591_36501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21585 VSS a_3891_25623# a_4068_25615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21586 VDD a_2840_55509# a_2787_55535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21587 VDD a_11921_35286# a_10985_35516# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X21588 a_45829_35407# a_45475_35520# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21589 a_48682_58500# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2159 a_37146_69182# a_18162_69222# a_37238_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21590 a_48190_9898# pmat.row_n[1] a_48682_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21591 a_24719_35253# a_11041_36596# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21592 VSS a_22199_30287# a_31203_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21593 a_21478_12870# pmat.rowoff_n[4] a_21082_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21594 VSS pmat.row_n[3] a_48586_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21595 VSS a_12437_28585# a_15585_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21596 vcm a_18162_7484# a_50290_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21597 VDD a_3305_27791# a_4443_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21598 a_6159_77295# a_5713_77295# a_6063_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21599 a_26194_24552# a_18546_24550# a_26102_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X216 vcm a_18162_58178# a_36234_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2160 VSS pmat.row_n[1] a_39550_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21600 vcm a_18162_21540# a_23182_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21601 a_25190_66170# a_18546_66212# a_25098_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21602 a_46578_62194# pmat.rowon_n[6] a_46182_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21603 a_32126_10902# pmat.row_n[2] a_32618_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21604 VDD a_24719_36341# a_15049_36374# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21605 vcm a_18162_7484# a_26194_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21606 a_30514_68218# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21607 a_12135_16367# a_11619_16367# a_12040_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X21608 a_38601_49035# ANTENNA_fanout52_A.DIODE a_38515_49035# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X21609 a_3657_19453# a_3613_19061# a_3491_19465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2161 VDD a_16083_50069# a_17203_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21610 VDD pmat.rowon_n[2] a_25098_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21611 VSS a_2931_40277# a_1895_41018# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21612 a_19166_9492# a_18546_9490# a_19074_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21613 VDD a_13091_28327# a_24873_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21614 a_15144_35077# a_13985_34789# a_15048_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X21615 a_25494_11866# nmat.rowon_n[12] a_25098_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21616 a_9602_10422# a_2021_11043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X21617 a_12067_67279# a_3923_68021# a_11895_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X21618 a_4308_24135# a_4516_21531# a_4450_24310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21619 VDD a_14163_55295# a_14150_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2162 VDD a_4865_12533# a_5445_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.315e+12p ps=1.063e+07u w=1e+06u l=150000u M=2
X21620 VDD a_9075_28023# a_11961_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21621 VSS a_9075_28023# a_11711_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21622 a_17996_41831# a_16837_42043# a_17959_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X21623 a_45178_70186# a_18162_70226# a_45270_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21624 vcm a_18162_62194# a_26194_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21625 a_26102_66170# pmat.row_n[10] a_26594_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21626 a_37542_64202# pmat.rowon_n[8] a_37146_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21627 a_30210_60146# a_18546_60188# a_30118_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21628 VDD nmat.rowon_n[14] a_35138_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21629 a_30610_64524# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2163 a_10641_52815# a_10363_53153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21630 a_33526_59182# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21631 vcm a_18162_12504# a_44266_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21632 a_2834_36495# a_1757_36501# a_2672_36873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21633 VDD nmat.rowon_n[2] a_35138_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21634 VSS a_12715_51420# a_12646_51549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21635 a_38242_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21636 VDD pmat.rowoff_n[12] a_48190_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21637 a_20570_56492# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21638 a_22178_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21639 a_48190_61150# a_18162_61190# a_48282_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2164 a_32126_57134# pmat.row_n[1] a_32618_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21640 a_4124_28023# a_4068_25615# a_4266_28157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21641 VDD a_1899_35051# a_6641_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21642 a_11409_28585# a_5991_23983# a_11337_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21643 a_21174_12504# a_18546_12502# a_21082_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21644 a_33622_9460# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21645 a_31122_60146# pmat.row_n[4] a_31614_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21646 VDD pmat.rowoff_n[4] a_38150_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21647 a_40250_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21648 VSS a_36341_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21649 vcm a_18162_68218# a_25190_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2165 vcm a_18162_14512# a_20170_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21650 a_36234_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21651 a_49194_24958# a_18162_24552# a_49286_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21652 a_8695_63937# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21653 a_12335_58255# a_1957_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21654 vcm a_18162_18528# a_43262_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21655 a_41321_30511# a_40967_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21656 a_6978_58799# a_3339_70759# a_7168_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21657 a_49286_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21658 VSS a_17536_38567# a_17499_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21659 a_6128_59887# a_5731_58951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2166 a_19267_28879# a_18795_28882# a_19165_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X21660 a_26272_41831# a_25209_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21661 VSS pmat.row_n[5] a_45574_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21662 VSS a_6607_10615# a_5768_9527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X21663 a_42562_17890# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21664 a_41237_28585# a_24747_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21665 VSS pmat.row_n[15] a_28506_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21666 a_25190_11500# a_18546_11498# a_25098_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21667 a_3295_40277# a_3659_39733# a_3431_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X21668 a_7829_71317# a_7663_71317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21669 a_23090_21946# a_18162_21540# a_23182_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2167 a_41254_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21670 a_26194_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21671 a_2099_8725# a_1979_9334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21672 a_29915_51183# a_13091_28327# pmat.col[10] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21673 a_35161_49007# a_26891_28327# nmat.col[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21674 cgen.dlycontrol1_in[1] a_1591_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21675 vcm a_18162_59182# a_46274_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21676 VSS a_9335_51727# a_10491_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X21677 a_2629_67503# a_2250_67869# a_2557_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21678 a_6891_15279# a_6541_15279# a_6796_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21679 a_28876_47741# a_28639_47081# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2168 a_43566_55166# VSS a_43170_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21680 a_29206_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21681 a_50290_57134# a_18546_57176# a_50198_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21682 a_22482_61190# pmat.rowon_n[5] a_22086_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21683 a_19166_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21684 a_46578_16886# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21685 VDD a_11611_50332# a_11542_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21686 a_1899_76001# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X21687 VSS a_11697_56775# a_8749_57141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21688 VSS pmat.row_n[6] a_50594_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21689 a_44174_10902# a_18162_10496# a_44266_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2169 a_43261_48783# a_33423_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X21690 VSS VDD a_33526_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21691 a_30514_21906# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21692 a_27106_20942# a_18162_20536# a_27198_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21693 a_38150_69182# a_18162_69222# a_38242_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21694 VDD pmat.rowon_n[6] a_37146_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21695 VSS config_1_in[8] a_1591_6031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21696 a_33130_57134# pmat.row_n[1] a_33622_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21697 a_42258_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21698 a_23182_59142# a_18546_59184# a_23090_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21699 vcm a_18162_56170# a_20170_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X217 VDD pmat.rowon_n[15] a_40158_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2170 a_46845_44111# a_40105_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=0p ps=0u w=1e+06u l=150000u
X21700 a_83094_10089# _1184_.A2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21701 a_36270_50095# _1154_.A pmat.col_n[16] VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u w=650000u l=150000u
X21702 a_8291_23983# a_7847_24233# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X21703 a_5197_16121# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21704 a_19470_18894# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21705 VSS a_1586_18231# a_1591_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21706 VSS pmat.row_n[8] a_23486_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21707 a_28572_44007# a_27509_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21708 VSS a_2595_13621# a_2526_13647# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21709 a_20474_13874# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2171 VSS ANTENNA__1395__A2.DIODE a_31847_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X21710 VDD a_18823_50247# a_19439_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21711 VDD a_39981_37462# a_39045_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X21712 a_21174_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21713 VDD a_16045_37692# a_15651_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21714 VDD a_38905_28853# a_38933_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21715 a_33526_12870# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21716 a_45574_63198# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21717 VSS pmat.row_n[13] a_35534_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21718 vcm a_18162_55166# a_24186_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21719 a_24921_27221# _1192_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2172 a_26498_65206# pmat.rowon_n[9] a_26102_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21720 a_24094_59142# pmat.row_n[3] a_24586_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21721 VSS a_34002_34191# a_34639_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21722 VDD config_2_in[4] a_1591_35951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X21723 VSS VDD a_36538_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21724 a_1846_59051# a_2124_59067# a_2080_59165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21725 a_9367_50871# a_9463_50877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21726 VSS a_6821_18543# a_9227_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21727 a_43170_22950# pmat.row_n[14] a_43662_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21728 a_36234_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21729 VDD pmat.rowoff_n[15] a_50198_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2173 VDD pmat.rowon_n[5] a_49194_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21730 VSS pmat.row_n[7] a_22482_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21731 VSS a_10641_52815# a_11829_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21732 a_46578_7850# VDD a_46182_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21733 a_19166_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21734 a_50198_64162# a_18162_64202# a_50290_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21735 a_35559_30209# a_6283_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21736 a_36538_65206# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21737 a_26456_41605# a_25393_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21738 a_49286_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21739 a_36634_17492# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2174 vcm a_18162_13508# a_33222_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21740 a_36538_23914# pmat.rowoff_n[15] a_36142_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21741 a_25190_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21742 a_10233_7913# a_10378_7637# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21743 VDD a_12905_17973# a_12795_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21744 vcm.sky130_fd_sc_hd__buf_4_2.A vcm.sky130_fd_sc_hd__dlymetal6s6s_1_5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21745 VDD pmat.rowoff_n[7] a_40158_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21746 a_23301_47349# a_23083_47753# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21747 VSS config_2_in[14] a_1591_50639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21748 a_49590_64202# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21749 a_34530_7850# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2175 a_4433_40125# a_2935_38279# a_4351_39872# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21750 VSS a_2283_39189# a_1895_38842# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X21751 a_47186_21946# pmat.row_n[13] a_47678_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21752 VSS a_2791_57703# a_2757_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21753 a_47186_17930# a_18162_17524# a_47278_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21754 VSS a_22269_40391# a_22743_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21755 VSS pmat.row_n[1] a_27502_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21756 a_51294_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21757 a_39550_56170# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21758 a_13253_42693# a_13561_42333# a_13227_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21759 a_41162_66170# a_18162_66210# a_41254_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2176 VDD a_9317_47349# a_9207_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X21760 a_37146_13914# pmat.row_n[5] a_37638_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21761 a_38150_7890# a_18162_7484# a_38242_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21762 a_7186_25615# a_6747_25731# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X21763 a_29510_67214# pmat.rowon_n[11] a_29114_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21764 a_41654_11468# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21765 VSS pmat.row_n[8] a_26498_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21766 a_13768_22325# a_13467_21263# a_13717_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=0p ps=0u w=1e+06u l=150000u
X21767 VSS a_10055_31591# a_15916_52277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21768 a_24586_21508# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21769 a_24186_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2177 VDD a_79368_39738# a_79181_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21770 a_32589_47375# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21771 a_27106_65166# a_18162_65206# a_27198_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21772 VSS a_44444_32233# a_46897_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21773 VSS a_26957_37691# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21774 a_31214_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21775 a_19470_59182# pmat.rowon_n[3] a_19074_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21776 a_31518_70226# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21777 VSS a_10569_64489# a_10707_64783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21778 a_35230_63158# a_18546_63200# a_35138_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21779 VDD a_20310_28029# a_22265_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2178 a_20170_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21780 a_47453_36815# a_38851_28327# a_46636_36469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21781 a_11981_14191# a_10791_14191# a_11872_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X21782 a_35630_67536# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21783 a_27598_12472# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21784 a_4254_7351# a_4003_7663# a_4241_7663# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X21785 a_40678_31599# a_38913_31055# a_40592_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21786 a_25098_13914# a_18162_13508# a_25190_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21787 VDD nmat.rowon_n[13] a_31122_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21788 a_48282_62154# a_18546_62196# a_48190_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21789 a_48682_66532# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2179 VDD ANTENNA__1190__A2.DIODE a_14289_4649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X21790 a_45178_63158# pmat.row_n[7] a_45670_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21791 a_17959_42089# a_16837_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21792 a_21478_62194# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21793 a_15324_41831# a_14261_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21794 a_34530_61190# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21795 VSS pmat.row_n[14] a_35534_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21796 a_4918_34319# a_4831_34561# a_4514_34451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21797 vcm a_18162_71230# a_22178_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21798 a_16911_51959# a_17183_51817# a_17141_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21799 VSS a_11902_56775# a_11697_56775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_32126_17930# pmat.row_n[9] a_32618_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2180 a_10319_7663# a_9668_10651# a_9827_8181# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X21800 VDD pmat.rowon_n[0] a_42166_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21801 VDD a_5307_67655# a_7073_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21802 a_2867_43541# a_1957_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21803 a_4719_69929# a_2419_69455# a_4801_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21804 a_46217_52815# a_11067_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X21805 a_4583_27830# a_4068_25615# a_4124_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21806 VDD pmat.rowon_n[10] a_25098_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21807 a_22578_63520# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21808 VSS a_33109_52245# pmat.col[13] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21809 a_33925_29199# a_13641_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2181 VSS a_1644_34293# a_1586_33927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21810 a_49194_62154# pmat.row_n[6] a_49686_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21811 a_3983_47919# a_4128_46983# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21812 VDD a_1858_25615# a_2511_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21813 a_23182_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21814 a_25190_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21815 a_47278_68178# a_18546_68220# a_47186_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21816 a_18180_38341# a_17021_38053# a_18084_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X21817 a_36617_43131# a_35752_43781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21818 a_6649_41935# a_6619_41909# a_6554_43255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X21819 vcm a_18162_70226# a_26194_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2182 a_2107_28169# a_1591_27797# a_2012_28157# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X21820 VSS a_20695_32447# a_20629_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21821 vcm a_18162_9492# a_41254_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21822 a_37542_72234# VDD a_37146_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21823 a_44801_35773# a_43776_30287# a_44729_35773# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21824 a_30610_72556# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21825 vcm a_18162_20536# a_44266_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21826 VDD pmat.rowon_n[9] a_29114_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21827 a_26594_62516# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21828 VSS a_9963_13967# a_13814_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X21829 a_44562_46070# a_29937_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2183 VDD a_2791_57703# a_2971_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X21830 VDD pmat.rowon_n[4] a_30118_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21831 a_9823_10749# a_9675_10396# a_9460_10615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21832 VSS a_40105_47375# a_47026_45519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21833 a_51294_9492# a_18546_9490# a_51202_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21834 a_51598_67214# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21835 VSS a_9463_8439# a_8243_7290# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21836 VDD a_9919_57863# a_9577_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X21837 VSS a_19582_46983# a_19531_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21838 VDD pmat.rowon_n[1] a_19074_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21839 a_13335_31359# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 a_32522_12870# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21840 nmat.rowoff_n[3] a_13551_8751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21841 a_29510_20902# pmat.rowoff_n[12] a_29114_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21842 VDD a_14071_74879# a_14058_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21843 a_47207_35951# a_46934_35951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21844 a_41558_59182# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21845 a_21174_20536# a_18546_20534# a_21082_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21846 VSS a_9581_73487# a_9873_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21847 a_41558_17890# nmat.rowon_n[6] a_41162_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21848 a_5603_18543# a_5253_18543# a_5508_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21849 a_24490_69222# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2185 a_44570_63198# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21850 a_25743_49783# a_25802_48169# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21851 a_48586_23914# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21852 a_29183_36919# a_28061_36965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21853 a_19470_12870# pmat.rowoff_n[4] a_19074_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21854 a_49286_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21855 VDD a_7405_32441# a_7435_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21856 VDD a_15439_48071# a_14528_48114# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X21857 a_42258_56130# a_18546_56172# a_42166_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21858 VDD a_2764_45577# a_2939_45503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21859 a_25098_58138# a_18162_58178# a_25190_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2186 a_4679_28853# a_5038_28853# a_4815_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X21860 VSS a_33341_37692# a_33033_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21861 a_39154_71190# a_18162_71230# a_39246_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21862 a_38546_15882# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21863 VSS a_1858_25615# a_15065_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21864 a_11559_68619# a_10864_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21865 a_45574_16886# nmat.rowon_n[7] a_45178_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21866 VSS pmat.row_n[5] a_42562_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21867 a_32507_47695# a_30999_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21868 VSS a_1957_43567# a_12489_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21869 a_25098_17930# pmat.row_n[9] a_25590_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2187 VSS a_25575_31055# a_41121_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21870 VDD cgen.dlycontrol4_in[0] a_1945_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21871 VDD nmat.rowon_n[5] a_32126_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21872 vcm a_18162_67214# a_46274_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21873 VDD a_27313_51701# pmat.col_n[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21874 a_13446_14191# a_9963_13967# a_13277_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21875 a_2325_38645# a_2107_39049# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21876 a_31303_27497# a_25879_31591# a_31085_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21877 VSS a_35465_32441# a_35399_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21878 a_50290_65166# a_18546_65208# a_50198_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21879 a_50690_69544# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2188 VSS a_18563_27791# a_41192_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21880 a_46274_55126# a_18546_55168# a_46182_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21881 a_46674_59504# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21882 VSS a_3339_59879# a_10989_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21883 a_2464_74397# a_2250_74397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21884 VDD a_12557_30485# a_12587_30838# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21885 a_29536_47753# a_28455_47381# a_29189_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21886 vcm a_18162_8488# a_30210_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21887 VDD pmat.rowon_n[14] a_37146_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21888 vcm a_18162_69222# a_19166_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21889 a_29114_16926# pmat.row_n[8] a_29606_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2189 a_3158_13647# a_2439_13889# a_2595_13621# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X21890 a_9460_10615# a_9675_10396# a_9602_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21891 a_6612_65845# a_2407_49289# a_6832_66191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21892 a_27236_46831# a_26155_46831# a_26889_47073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21893 a_41162_9898# a_18162_9492# a_41254_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21894 a_44976_47349# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21895 a_23182_67174# a_18546_67216# a_23090_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21896 a_30118_11906# pmat.row_n[3] a_30610_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21897 vcm a_18162_64202# a_20170_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21898 a_14655_53359# a_11067_64015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21899 VSS a_4337_22351# a_4259_24643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X219 VSS pmat.row_n[15] a_32522_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2190 a_11793_71311# a_9279_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21900 a_20078_68178# pmat.row_n[12] a_20570_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21901 a_19166_57134# a_18546_57176# a_19074_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21902 VSS a_17154_43671# a_17159_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21903 a_41254_17524# a_18546_17522# a_41162_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21904 a_51202_65166# pmat.row_n[9] a_51694_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21905 VDD pmat.rowon_n[3] a_23090_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21906 VDD a_6979_51157# a_6883_51335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21907 VSS a_18769_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21908 a_51294_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21909 VSS pmat.row_n[6] a_19470_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2191 a_7167_52105# a_6651_51733# a_7072_52093# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X21910 a_3026_41213# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21911 VSS a_25695_28111# a_37737_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21912 a_22522_50247# a_22499_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21913 a_35007_44527# a_34830_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21914 a_12034_14557# a_10957_14191# a_11872_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21915 VDD a_39089_27765# nmat.col[20] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21916 a_41162_57134# pmat.row_n[1] a_41654_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21917 VSS a_12079_9615# a_14839_9295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21918 a_37754_30511# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21919 VSS pmat.rowon_n[7] a_14734_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2192 a_47186_8894# a_18162_8488# a_47278_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21920 a_4993_77071# a_4951_76983# a_4123_76181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X21921 vcm a_18162_63198# a_24186_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21922 a_20310_28029# a_20695_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21923 VSS a_6179_65479# a_5495_65479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X21924 a_51598_20902# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21925 a_24094_67174# pmat.row_n[11] a_24586_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21926 a_10287_24759# a_10651_24617# a_10586_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21927 a_35534_65206# pmat.rowon_n[9] a_35138_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21928 a_45270_16520# a_18546_16518# a_45178_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21929 vcm a_18162_13508# a_42258_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2193 vcm a_18162_72234# a_45270_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21930 a_11149_40188# a_33255_43777# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21931 a_2847_8511# a_2672_8585# a_3026_8573# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21932 a_48586_64202# pmat.rowon_n[8] a_48190_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21933 VDD a_11910_43047# a_11915_42895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21934 a_41558_12870# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21935 VDD nmat.rowon_n[2] a_46182_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21936 a_30457_37479# a_30765_37692# a_30431_37683# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21937 a_24490_22910# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21938 VSS a_18272_39429# a_18235_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21939 a_49286_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2194 a_42166_7890# VDD a_42658_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21940 a_3123_69135# a_3069_69367# a_3029_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X21941 a_38546_56170# pmat.rowon_n[0] a_38150_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21942 a_46815_37013# a_35244_32411# a_47321_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21943 a_31614_56492# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21944 a_49590_72234# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21945 a_14370_15279# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21946 VDD nmat.rowon_n[10] a_36142_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21947 a_33489_42043# a_30523_41245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X21948 a_11703_48156# a_11547_48061# a_11848_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21949 a_47861_51727# a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2195 a_11207_31764# a_11299_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21950 a_9919_51959# a_9213_53903# a_10388_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21951 a_32218_12504# a_18546_12502# a_32126_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21952 a_7201_62063# a_5784_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21953 a_51294_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21954 a_6723_37405# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21955 a_47278_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21956 VDD a_2563_34837# a_5043_37191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21957 a_43965_27221# a_27763_27221# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21958 VDD a_11113_39747# a_34552_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X21959 VSS a_4383_7093# a_3551_6202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2196 a_42166_22950# pmat.row_n[14] a_42658_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21960 VSS pmat.row_n[6] a_43566_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21961 a_40554_18894# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21962 vcm a_18162_14512# a_19166_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21963 a_37542_9858# nmat.rowon_n[14] a_37146_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21964 a_10422_24643# a_9528_20407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21965 VSS VDD a_26498_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21966 a_29635_31029# a_30219_29967# a_30205_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.1e+11p pd=3.22e+06u as=0p ps=0u w=1e+06u l=150000u
X21967 a_30514_70226# pmat.rowon_n[14] a_30118_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21968 a_44266_71190# a_18546_71232# a_44174_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21969 VDD a_10864_68565# a_11541_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2197 a_35230_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21970 a_10233_50639# a_8385_51727# a_9457_51163# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21971 a_10209_22351# a_10071_17999# a_10055_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21972 VDD VSS a_44174_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21973 a_2241_39465# a_1899_35051# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21974 a_20474_62194# pmat.rowon_n[6] a_20078_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21975 a_36373_50095# a_30663_50087# a_36270_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X21976 VSS a_13091_50095# a_13278_51549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21977 a_31323_29967# a_31072_30083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21978 a_33526_61190# pmat.rowon_n[5] a_33130_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21979 a_6628_77295# a_5547_77295# a_6281_77537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2198 pmat.row_n[8] a_19675_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X21980 a_41883_47081# a_13275_48783# a_41665_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21981 VDD a_2007_49770# a_1895_50308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X21982 a_3583_11775# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21983 a_48282_70186# a_18546_70228# a_48190_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21984 a_44082_31599# a_41949_30761# a_43996_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21985 VDD a_3331_59317# a_3262_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21986 a_11358_73309# a_11271_73085# a_10954_73195# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21987 a_45178_71190# pmat.row_n[15] a_45670_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21988 a_46182_7890# a_18162_7484# a_46274_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21989 a_45670_20504# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2199 VSS a_33839_46805# a_40047_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21990 a_8703_6202# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21991 a_45270_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21992 a_3569_72765# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21993 a_10999_36694# a_10817_36694# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21994 VSS a_36341_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X21995 VDD pmat.rowon_n[6] a_48190_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21996 a_17867_44535# a_16745_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21997 a_34226_59142# a_18546_59184# a_34134_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21998 a_11230_48171# a_11547_48061# a_11505_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21999 a_35630_12472# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u M=1806
X220 VSS a_10985_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X2200 VDD pmat.rowon_n[11] a_48190_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22000 VDD a_2683_22089# a_8097_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22001 a_10391_62911# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22002 VSS pmat.row_n[8] a_34530_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22003 VDD a_6283_31591# a_26155_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22004 a_32218_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22005 VSS a_25997_42902# a_25061_43132# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X22006 a_22578_71552# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22007 a_39246_22544# a_18546_22542# a_39154_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22008 a_49194_70186# pmat.row_n[14] a_49686_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22009 VDD pmat.rowoff_n[12] a_22086_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2201 VSS pmat.row_n[7] a_21478_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22010 a_28812_29575# a_37795_29111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22011 a_46182_12910# a_18162_12504# a_46274_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22012 VSS a_14497_42658# a_13561_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X22013 a_12133_9001# a_11051_8903# a_12061_9001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22014 a_25190_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22015 a_22086_61150# a_18162_61190# a_22178_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22016 VSS pmat.row_n[13] a_46578_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22017 a_43566_66210# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22018 a_8378_63827# a_8656_63811# a_8612_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22019 a_32126_8894# pmat.row_n[0] a_32618_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2202 a_36538_7850# VDD a_36142_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22020 a_50594_67214# pmat.rowon_n[11] a_50198_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22021 vcm a_18162_55166# a_35230_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22022 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22023 a_5547_24233# a_4337_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22024 a_14691_29575# a_14751_28341# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X22025 a_35138_59142# pmat.row_n[3] a_35630_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22026 a_2369_39037# a_2325_38645# a_2203_39049# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22027 VDD a_24867_53135# a_35269_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22028 VDD a_4503_70455# a_4421_70741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X22029 a_26498_8854# nmat.rowon_n[15] a_26102_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2203 a_18162_68218# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X22030 a_14734_4175# _1183_.A2 a_14565_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22031 a_11713_64899# a_10921_64786# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22032 a_13961_72765# a_13917_72373# a_13795_72777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22033 a_26594_70548# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22034 a_47278_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22035 a_19074_14918# a_18162_14512# a_19166_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22036 a_40554_59182# pmat.rowon_n[3] a_40158_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22037 a_23182_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22038 a_5069_40303# a_4705_39759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22039 VDD a_3429_76725# a_3319_76751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2204 a_21087_43177# a_21124_42919# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X22040 a_23486_69222# pmat.rowon_n[13] a_23090_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22041 a_26102_60146# a_18162_60186# a_26194_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22042 VSS a_2319_52789# a_2250_52815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22043 VSS a_19405_28853# a_19083_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22044 VSS a_4955_40277# a_5921_44629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22045 a_5257_69679# a_4719_69929# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22046 a_47582_65206# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22047 vcm a_18162_17524# a_30210_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22048 a_47678_17492# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22049 a_9651_62985# a_9135_62613# a_9556_62973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2205 a_48282_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22050 VDD pmat.rowoff_n[7] a_51202_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22051 a_45178_18934# a_18162_18528# a_45270_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22052 a_9225_71855# a_9183_72007# a_8283_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X22053 a_37542_57174# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22054 VDD a_22059_37683# a_22085_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22055 VDD nmat.rowon_n[13] a_29114_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22056 a_44570_58178# pmat.rowon_n[2] a_44174_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22057 VSS a_21219_36885# a_21031_37217# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22058 VSS VDD a_41558_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22059 VSS a_34948_50069# pmat.col[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X2206 a_40041_27791# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X22060 VDD a_24937_36039# a_25628_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22061 VSS a_2944_69928# a_2882_70045# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22062 a_27502_68218# pmat.rowon_n[12] a_27106_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22063 a_2325_20149# a_2107_20553# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22064 VSS pmat.row_n[9] a_24490_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22065 vcm a_18162_16520# a_34226_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22066 VDD a_2319_72092# a_2250_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22067 vcm a_18162_66210# a_38242_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22068 a_48190_13914# pmat.row_n[5] a_48682_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22069 VSS a_20616_27791# a_23021_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2207 VDD a_5363_33551# a_6651_33239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22070 a_22178_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22071 a_42258_64162# a_18546_64204# a_42166_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22072 nmat.rowoff_n[13] a_11067_16359# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22073 a_38642_19500# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22074 a_42658_68540# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22075 VDD a_4553_18297# a_4583_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22076 a_3568_74575# a_3354_74575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22077 VDD a_45019_38645# a_44515_38645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22078 VSS a_2847_41151# a_2781_41225# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X22079 VDD a_6283_31591# a_22567_47381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2208 a_6242_67503# a_5403_67655# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X22080 VSS pmat.row_n[0] a_27502_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22081 VDD pmat.rowon_n[5] a_24094_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22082 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22083 VDD nmat.rowon_n[7] a_28110_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22084 a_19487_49159# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22085 a_4241_13653# a_4075_13653# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22086 a_14000_47695# a_11067_64015# a_13697_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22087 VSS a_21977_52245# pmat.col[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22088 a_2655_72373# a_2858_72531# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22089 a_46274_63158# a_18546_63200# a_46182_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2209 a_7935_20719# a_7048_23277# a_7935_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=4.1e+11p ps=2.82e+06u w=1e+06u l=150000u
X22090 vcm a_18162_60186# a_43262_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22091 a_5760_54991# a_5730_54965# a_5658_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22092 a_46674_67536# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22093 a_43170_64162# pmat.row_n[8] a_43662_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22094 a_6641_44111# a_2659_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22095 VDD a_45325_38127# a_47357_38127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22096 VDD pmat.rowon_n[9] a_50198_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22097 a_55770_39250# comp.adc_nor_latch_0.R VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22098 a_79085_39738# a_79181_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22099 a_46182_57134# a_18162_57174# a_46274_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X221 a_29206_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2210 VSS pmat.row_n[6] a_34530_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22100 VSS nmat.sw a_10383_13077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X22101 a_32522_62194# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22102 VSS a_3688_17179# a_8399_18115# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22103 VDD a_4383_7093# a_12069_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22104 a_7258_8751# a_7040_8725# a_7176_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22105 a_10702_32143# a_9944_32259# a_10139_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22106 VDD a_2046_30184# a_2787_33237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22107 a_29114_67174# a_18162_67214# a_29206_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22108 vcm a_18162_72234# a_20170_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22109 a_16926_46261# a_12447_16143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2211 a_35630_17492# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22110 a_10140_67503# a_9545_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22111 a_19166_65166# a_18546_65208# a_19074_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22112 VDD pmat.rowon_n[1] a_40158_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22113 VSS pmat.row_n[14] a_46578_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22114 VDD a_7899_67477# a_7803_67655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22115 a_19566_69544# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22116 a_50690_14480# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22117 a_40250_8488# a_18546_8486# a_40158_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22118 a_50594_20902# pmat.rowoff_n[12] a_50198_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22119 vcm a_18162_71230# a_33222_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2212 a_35534_23914# pmat.rowoff_n[15] a_35138_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22120 VDD pmat.rowon_n[11] a_23090_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22121 a_37238_15516# a_18546_15514# a_37146_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22122 VSS a_10515_15055# pmat.rowon_n[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22123 a_19074_59142# a_18162_59182# a_19166_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22124 a_33622_24520# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22125 a_2199_45577# a_1683_45205# a_2104_45565# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X22126 VSS a_12345_39100# a_12764_39453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22127 a_23182_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22128 a_44420_45895# a_44635_46025# a_44562_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22129 a_39550_17890# nmat.rowon_n[6] a_39154_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2213 a_22178_72194# a_18546_72236# a_22086_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22130 VSS a_13503_43421# a_13443_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22131 a_40554_12870# pmat.rowoff_n[4] a_40158_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22132 a_7809_17705# a_7407_17455# a_7645_17455# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X22133 a_6799_75637# a_6803_77269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22134 a_37146_55126# VDD a_37638_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22135 a_12568_35077# a_11409_34789# a_12472_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22136 VSS a_2944_61493# a_2882_61519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22137 a_23486_22910# nmat.rowon_n[1] a_23090_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22138 a_21082_21946# pmat.row_n[13] a_21574_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22139 a_21082_17930# a_18162_17524# a_21174_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2214 VSS pmat.sample a_18546_70228# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X22140 vcm a_18162_21540# a_42258_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22141 a_45270_24552# a_18546_24550# a_45178_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22142 a_51202_10902# pmat.row_n[2] a_51694_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22143 vcm a_18162_11500# a_38242_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22144 a_15420_41831# a_14261_42043# a_15383_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22145 VSS a_4313_44111# a_4837_45519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22146 VDD a_29536_47753# a_29711_47679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22147 a_48586_72234# VDD a_48190_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22148 a_34134_20942# pmat.row_n[12] a_34626_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22149 a_34134_16926# a_18162_16520# a_34226_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2215 a_28602_7452# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22150 a_45475_52271# _1192_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22151 a_5451_14557# a_5271_14557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22152 VDD pmat.rowon_n[2] a_44174_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22153 a_37542_10862# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22154 a_5779_13255# a_4895_12559# a_6013_13103# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X22155 VDD a_27236_46831# a_27411_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22156 a_44570_11866# nmat.rowon_n[12] a_44174_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22157 a_3939_16950# a_3688_17179# a_3480_17143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22158 VSS a_37519_46983# a_36539_47113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X22159 a_24094_12910# pmat.row_n[4] a_24586_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2216 a_24490_7850# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X22160 a_27502_21906# nmat.rowon_n[2] a_27106_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22161 VSS a_2419_53351# a_5157_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22162 vcm a_18162_22544# a_28202_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22163 a_18546_16518# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X22164 a_83362_12265# _1194_.A2 a_82971_11989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22165 a_32218_20536# a_18546_20534# a_32126_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22166 VSS a_24937_43655# a_26331_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22167 vcm a_18162_69222# a_40250_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22168 a_9367_50871# a_8385_51727# a_9601_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22169 a_50198_16926# pmat.row_n[8] a_50690_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2217 VSS a_26479_32117# a_42307_31756# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=5.88e+06u w=650000u l=150000u M=2
X22170 a_35534_69222# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22171 VSS a_44444_32233# a_44320_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22172 a_45554_52815# ANTENNA__1190__B1.DIODE a_45251_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22173 a_5683_30333# a_5535_29980# a_5320_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22174 VDD a_2007_8916# a_1895_8378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22175 a_37146_72194# a_18162_72234# a_37238_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22176 a_24015_36911# cgen.dlycontrol3_in[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X22177 VSS pmat.row_n[4] a_39550_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22178 a_46027_44905# a_44966_43255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22179 VSS pmat.row_n[11] a_39550_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2218 a_48586_22910# nmat.rowon_n[1] a_48190_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22180 a_41254_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22181 a_14647_51701# a_14491_51969# a_14792_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22182 a_27598_9460# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22183 VDD a_5266_17143# a_5451_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22184 VSS a_2122_19087# a_2228_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22185 a_10873_36341# a_29391_36395# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X22186 a_40250_12504# a_18546_12502# a_40158_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22187 a_23090_18934# pmat.row_n[10] a_23582_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22188 vcm a_18162_68218# a_44266_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22189 a_2672_41225# a_1591_40853# a_2325_40821# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2219 a_46182_21946# pmat.row_n[13] a_46674_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22190 VDD _1154_.A a_47449_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22191 a_5297_34685# a_4918_34319# a_5225_34685# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X22192 a_4713_38377# a_3325_40847# a_4617_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22193 a_44266_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22194 a_45469_53135# _1192_.B1 a_45251_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22195 a_8197_76757# a_8031_76757# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22196 a_27198_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22197 VSS pmat.row_n[2] a_33526_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22198 a_30514_55166# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22199 VDD a_9411_2215# a_25139_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X222 a_39154_7890# a_18162_7484# a_39246_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2220 VSS a_5323_71829# a_5271_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22200 a_26501_37462# a_25393_38053# a_26456_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22201 a_45077_32687# a_38851_28327# a_45005_32687# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X22202 VSS a_2163_65469# a_2124_65595# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22203 a_21174_68178# a_18546_68220# a_21082_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22204 a_15857_27791# a_14947_26159# a_15667_28111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22205 a_29635_31029# a_30412_31751# a_30121_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22206 a_39550_8854# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22207 a_42166_21946# a_18162_21540# a_42258_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22208 a_45270_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22209 VSS a_2007_21482# a_1895_20346# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2221 a_50198_70186# pmat.row_n[14] a_50690_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22210 VDD pmat.rowon_n[14] a_48190_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22211 a_7210_11837# a_2021_9563# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22212 a_38150_11906# a_18162_11500# a_38242_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22213 a_34226_67174# a_18546_67216# a_34134_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22214 a_3797_14709# a_3579_15113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22215 a_24861_52047# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22216 a_27106_19938# pmat.row_n[11] a_27598_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22217 a_7824_31433# a_6743_31061# a_7477_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22218 a_29067_47753# a_28621_47381# a_28971_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22219 a_48282_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2222 VDD a_12985_62581# a_5462_62215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X22220 VSS pmat.row_n[0] a_49590_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22221 a_40868_29423# a_24747_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22222 a_24490_71230# pmat.rowon_n[15] a_24094_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22223 cgen.dlycontrol2_in[1] a_1591_38127# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22224 a_4843_54826# a_8477_57141# a_8507_57487# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u M=2
X22225 VSS a_3325_40847# a_3659_39733# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X22226 a_46182_20942# a_18162_20536# a_46274_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22227 a_4220_62037# a_4509_62037# a_4443_62063# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X22228 vcm a_18162_19532# a_39246_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22229 vcm a_18162_14512# a_40250_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2223 a_46182_17930# a_18162_17524# a_46274_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22230 vcm a_18162_63198# a_35230_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22231 a_35138_67174# pmat.row_n[11] a_35630_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22232 a_46578_65206# pmat.rowon_n[9] a_46182_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22233 a_4149_41941# a_3983_41941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22234 a_19086_34343# a_19565_35279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22235 a_23823_47679# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X22236 a_40250_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22237 a_22482_23914# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22238 a_19074_22950# a_18162_22544# a_19166_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22239 a_41192_28995# a_24747_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2224 a_4075_31591# a_7939_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X22240 a_23182_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22241 a_36538_57174# pmat.rowon_n[1] a_36142_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22242 a_35534_22910# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22243 a_2834_63695# a_1757_63701# a_2672_64073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22244 a_6281_77537# a_6063_77295# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22245 a_29206_18528# a_18546_18526# a_29114_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22246 VSS a_22199_30287# a_42151_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22247 VDD a_13227_42333# a_13253_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22248 a_2999_76922# a_4123_76181# a_4081_76457# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22249 a_6424_55687# a_5682_56311# a_6566_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2225 VSS a_12557_32441# a_12491_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22250 a_44665_45519# a_40105_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22251 a_43781_52245# a_16311_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22252 a_31299_29673# a_21365_27247# a_31217_29429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22253 VSS pmat.row_n[9] a_28506_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22254 a_32522_15882# pmat.rowoff_n[7] a_32126_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22255 a_3325_43023# a_2847_43327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22256 VSS pmat.row_n[7] a_41558_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22257 a_38242_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22258 VDD a_6612_66933# a_4298_67191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22259 VDD a_82789_26677# nmat.col[29] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2226 a_17927_48437# a_17397_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X22260 a_12581_69455# a_12719_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22261 a_20170_55126# a_18546_55168# a_20078_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22262 vcm a_18162_24552# a_34226_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22263 a_20570_59504# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22264 a_28506_7850# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22265 VDD a_7456_15279# a_7631_15253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22266 vcm a_18162_56170# a_29206_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22267 a_42258_72194# a_18546_72236# a_42166_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22268 a_14369_50345# a_13432_62581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22269 a_34828_36165# a_33765_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2227 a_50290_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22270 a_33622_58500# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22271 a_29510_13874# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22272 a_10111_30511# a_9761_30511# a_10016_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22273 VSS pmat.row_n[3] a_33526_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22274 a_38150_56130# a_18162_56170# a_38242_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22275 a_14749_47197# a_14486_46831# a_14336_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22276 a_50198_8894# a_18162_8488# a_50290_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22277 a_31518_62194# pmat.rowon_n[6] a_31122_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22278 VDD a_3571_13627# a_11619_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22279 VSS pmat.row_n[8] a_45574_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2228 VSS VDD a_34530_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22280 a_39154_23954# pmat.row_n[15] a_39646_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22281 VSS a_3423_74549# a_3354_74575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22282 a_43170_72194# VDD a_43662_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22283 a_39154_19938# a_18162_19532# a_39246_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22284 a_26102_8894# a_18162_8488# a_26194_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22285 a_43662_21508# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22286 a_40158_14918# a_18162_14512# a_40250_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22287 a_21082_7890# VDD a_21574_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22288 a_43262_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22289 a_14816_47919# a_5363_70543# a_14336_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2229 VDD pmat.sample_n a_18162_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X22290 VSS a_3615_71631# a_14197_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22291 a_46182_65166# a_18162_65206# a_46274_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22292 a_50290_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22293 VSS pmat.row_n[0] a_35534_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22294 a_32035_42089# a_30913_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22295 a_28506_60186# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22296 a_28506_19898# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22297 VDD a_6244_71829# a_5521_72373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22298 a_31614_7452# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22299 a_30118_70186# a_18162_70226# a_30210_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X223 VDD pmat.rowon_n[5] a_36142_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2230 a_13719_36649# a_13779_36595# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X22300 a_8267_49159# a_3746_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22301 a_18546_61192# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X22302 a_14094_60751# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22303 a_10965_58255# a_10878_58487# a_10090_58093# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22304 a_22482_64202# pmat.rowon_n[8] a_22086_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22305 VDD pmat.en_bit_n[0] a_36142_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22306 a_37238_23548# a_18546_23546# a_37146_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22307 VDD pmat.rowoff_n[7] a_49194_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22308 a_46674_12472# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22309 VSS a_9675_10396# a_11167_11177# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2231 a_36142_13914# pmat.row_n[5] a_36634_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22310 VDD nmat.rowon_n[2] a_20078_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22311 a_22015_48579# a_21215_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22312 a_44174_13914# a_18162_13508# a_44266_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22313 VDD nmat.rowon_n[13] a_50198_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22314 a_23182_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22315 a_20078_62154# a_18162_62194# a_20170_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22316 a_29606_22512# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22317 a_10754_15279# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22318 VSS a_11067_16359# pmat.rowon_n[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22319 a_19166_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2232 VSS a_4523_21276# a_11091_26311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X22320 VSS ANTENNA__1196__A2.DIODE a_13723_3087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22321 VDD pmat.rowoff_n[12] a_33130_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22322 VDD a_2149_45717# a_6093_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22323 a_7377_65577# a_4583_68021# a_5399_65479# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22324 a_33130_61150# a_18162_61190# a_33222_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22325 a_36538_10862# nmat.rowon_n[13] a_36142_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22326 a_19566_14480# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22327 vcm a_18162_71230# a_41254_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22328 a_14458_14191# a_10239_14183# a_14372_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22329 VDD pmat.rowoff_n[4] a_23090_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2233 a_40650_11468# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22330 vcm a_18162_61190# a_37238_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22331 VSS a_16837_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22332 a_21174_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22333 a_34134_24958# a_18162_24552# a_34226_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22334 a_28613_40229# a_28116_39655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22335 VDD pmat.rowon_n[10] a_44174_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22336 a_41654_63520# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22337 a_51598_59182# pmat.rowon_n[3] a_51202_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22338 a_34226_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22339 a_1895_36666# a_2467_35925# a_2425_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2234 VSS pmat.row_n[8] a_25494_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22340 VSS a_33007_38771# a_32947_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22341 a_14486_47919# a_11067_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22342 a_9207_47375# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22343 VSS pmat.row_n[5] a_30514_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22344 a_2250_74397# a_2163_74173# a_1846_74283# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22345 a_8479_11484# a_8511_10422# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22346 VDD nmat.rowon_n[12] a_27106_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22347 VSS a_5363_33551# a_19439_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22348 a_48586_57174# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22349 a_45670_62516# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2235 a_39646_55488# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22350 VSS a_8851_12533# a_8782_12559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X22351 a_50198_67174# a_18162_67214# a_50290_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22352 vcm a_18162_59182# a_31214_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22353 VSS a_2791_57703# a_3315_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X22354 VSS a_36753_46805# a_36687_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22355 a_31518_16886# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22356 a_10957_28879# a_10609_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X22357 a_40158_59142# a_18162_59182# a_40250_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22358 a_49686_19500# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22359 vcm a_18162_22544# a_36234_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2236 a_19074_23954# pmat.row_n[15] a_19566_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22360 a_23301_47349# a_23083_47753# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22361 a_40250_20536# a_18546_20534# a_40158_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22362 a_23090_69182# a_18162_69222# a_23182_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22363 VDD pmat.rowon_n[6] a_22086_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22364 a_36234_10496# a_18546_10494# a_36142_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22365 a_1644_76181# a_1823_76181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22366 VDD ANTENNA__1197__A.DIODE a_43999_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22367 a_6641_37583# a_6061_38377# a_6403_37252# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22368 VDD nmat.rowon_n[14] a_37146_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22369 a_27421_41814# a_26773_40955# a_27836_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2237 a_23090_72194# VDD a_23582_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22370 a_4608_41909# a_4432_42313# a_4752_42301# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22371 VDD a_5351_60663# a_4317_62215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X22372 VDD a_5455_22057# a_5899_21807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22373 a_6732_44111# a_4257_34319# a_6559_44431# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22374 VDD nmat.rowon_n[4] a_26102_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22375 a_44174_58138# a_18162_58178# a_44266_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22376 a_2939_11849# a_2493_11477# a_2843_11849# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22377 a_23663_39913# a_22541_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22378 a_30514_63198# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22379 a_19074_60146# pmat.row_n[4] a_19566_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2238 a_11785_16367# a_11619_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22380 a_27106_68178# a_18162_68218# a_27198_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22381 VSS a_6467_29415# a_7939_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X22382 VSS pmat.row_n[13] a_20474_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22383 VSS a_4705_39759# a_5757_40097# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22384 a_44174_17930# pmat.row_n[9] a_44666_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22385 VSS pmat.row_n[15] a_44570_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22386 a_13457_64757# a_13239_65161# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22387 a_20170_9492# a_18546_9490# a_20078_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22388 a_32802_47695# a_31152_48071# a_32507_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22389 a_19509_39638# a_19505_38779# a_20568_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2239 a_19074_19938# a_18162_19532# a_19166_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22390 a_39666_30287# a_39127_29423# a_39580_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22391 VDD pmat.rowon_n[1] a_51202_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22392 a_12149_56399# a_6927_30503# a_11711_56079# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X22393 a_20776_51959# a_18823_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22394 a_21174_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22395 a_35230_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22396 a_37542_18894# nmat.rowon_n[5] a_37146_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22397 a_9919_57863# a_10191_57691# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22398 a_13985_35877# a_13319_35507# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22399 a_21478_65206# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X224 a_1923_61759# a_4043_59861# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X2240 VDD a_1923_69823# a_2747_74549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22400 a_34226_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22401 VSS a_15420_44007# a_15383_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22402 a_21574_17492# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22403 a_21478_23914# pmat.rowoff_n[15] a_21082_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22404 a_11149_59887# a_9135_60967# a_10286_60405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22405 a_51598_12870# pmat.rowoff_n[4] a_51202_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22406 VDD a_2847_33749# a_2834_34141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22407 VSS config_2_in[4] a_1591_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22408 VDD a_13837_37981# a_13443_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22409 a_34530_64202# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2241 a_49194_12910# pmat.row_n[4] a_49686_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22410 a_48190_55126# VDD a_48682_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22411 VDD a_30431_37683# a_30457_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22412 a_38242_57134# a_18546_57176# a_38150_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22413 a_11837_68591# a_11559_68619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X22414 a_32126_21946# pmat.row_n[13] a_32618_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22415 a_32126_17930# a_18162_17524# a_32218_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22416 a_10405_64239# a_9405_66627# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22417 VDD pmat.rowon_n[3] a_42166_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22418 VDD a_24895_36341# a_24719_36341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22419 VSS a_10873_40693# a_10817_41046# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2242 a_23582_21508# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22420 VSS pmat.row_n[6] a_38546_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22421 VSS ANTENNA__1395__B1.DIODE a_22745_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22422 VSS a_45529_51157# pmat.col_n[26] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22423 a_10216_69679# a_9301_69679# a_9869_69921# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22424 a_24490_56170# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22425 a_27605_42693# a_27913_42333# a_27329_42902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X22426 VDD a_6168_18543# a_6343_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22427 a_3024_22717# a_2907_22522# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22428 VDD a_44966_43255# a_44917_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22429 a_25590_16488# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2243 _1196_.B1 a_44533_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u M=16
X22430 a_22086_13914# pmat.row_n[5] a_22578_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22431 a_48586_10862# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22432 VDD a_3576_17143# a_5545_17027# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22433 VDD a_2007_42644# a_1895_43194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22434 VDD a_9411_2215# a_34063_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22435 a_2500_30345# a_2217_29973# a_2405_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22436 VDD a_6281_77537# a_6171_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X22437 a_11004_55535# a_11202_55687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22438 a_35138_12910# pmat.row_n[4] a_35630_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22439 VDD a_2944_59048# a_2882_59165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2244 a_20078_14918# a_18162_14512# a_20170_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22440 a_4429_76751# a_3951_77055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22441 VSS a_4553_28089# a_4487_28157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22442 a_13319_26703# a_12449_22895# a_13211_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22443 VSS a_47731_36103# a_47592_35643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22444 a_10867_43447# a_10927_43421# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22445 a_1907_12342# a_1725_12342# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22446 a_2781_41225# a_1591_40853# a_2672_41225# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X22447 a_30913_42043# a_29036_41831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22448 a_7373_48695# a_7578_48553# a_7536_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22449 a_28506_13874# nmat.rowon_n[10] a_28110_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2245 a_23182_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22450 VSS a_18243_28327# a_28628_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22451 a_22307_27791# a_22056_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22452 a_20170_63158# a_18546_63200# a_20078_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22453 a_20570_67536# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22454 VDD a_4901_30753# a_4791_30877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22455 a_48190_72194# a_18162_72234# a_48282_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22456 VDD a_1781_9308# a_36919_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X22457 a_18603_47081# a_12263_50959# a_18521_46837# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22458 vcm a_18162_64202# a_29206_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22459 a_50690_56492# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2246 a_44266_21540# a_18546_21538# a_44174_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22460 a_13643_22671# a_13768_22325# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22461 a_29114_68178# pmat.row_n[12] a_29606_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22462 VDD a_5363_73807# a_5361_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22463 a_33222_62154# a_18546_62196# a_33130_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22464 a_33622_66532# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22465 a_15107_34743# a_13985_34789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22466 a_30118_63158# pmat.row_n[7] a_30610_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22467 VDD pmat.rowoff_n[15] a_38150_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22468 a_20170_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22469 a_51294_12504# a_18546_12502# a_51202_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2247 pmat.col[23] a_28131_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X22470 a_8283_71829# a_9183_72007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22471 VSS a_1923_53055# a_1881_53181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22472 VSS VDD a_38546_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22473 VDD a_13973_66933# a_13909_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22474 a_38150_64162# a_18162_64202# a_38242_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22475 a_26425_52521# ANTENNA__1190__B1.DIODE pmat.col_n[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22476 VSS pmat.row_n[14] a_20474_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22477 a_42258_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22478 VSS a_2163_58941# a_2124_59067# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22479 a_43566_9858# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 VDD a_5325_9269# a_4989_11079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22480 a_10478_25045# a_9441_20189# a_10693_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22481 a_48586_7850# VDD a_48190_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22482 VSS VDD a_45574_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22483 a_34134_62154# pmat.row_n[6] a_34626_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22484 a_19470_9858# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22485 a_40158_22950# a_18162_22544# a_40250_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22486 a_22195_52521# _1194_.A2 a_21977_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22487 a_39246_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22488 VSS a_3688_17179# a_7213_19407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22489 a_11987_24847# a_7026_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2249 a_26102_65166# a_18162_65206# a_26194_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22490 a_32218_68178# a_18546_68220# a_32126_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22491 a_19948_51959# a_12263_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22492 VSS pmat.row_n[1] a_29510_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22493 a_22482_72234# VDD a_22086_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22494 VSS a_2192_49159# a_2099_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22495 a_28202_13508# a_18546_13506# a_28110_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22496 vcm a_18162_10496# a_25190_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22497 VSS a_2215_47375# a_2879_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22498 a_24747_29967# a_24214_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X22499 a_13529_68841# a_12719_69367# a_13456_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 a_40250_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2250 VDD a_4383_7093# a_4341_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X22500 a_7355_31433# a_6909_31061# a_7259_31433# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X22501 a_6447_35229# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22502 a_19166_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22503 a_36538_60186# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22504 a_14372_5487# ANTENNA__1187__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22505 a_40532_39429# a_39469_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22506 a_36538_19898# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22507 a_3354_74575# a_3267_74817# a_2950_74707# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22508 a_19470_70226# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22509 vcm a_18162_56170# a_50290_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2251 a_31978_43439# a_31801_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22510 a_3583_11775# a_3408_11849# a_3762_11837# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22511 a_49590_18894# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22512 a_22541_44581# a_21032_44007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X22513 a_12605_28879# a_8583_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22514 a_24847_36367# a_12237_36596# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22515 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22516 a_2651_29098# a_2743_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X22517 a_50594_13874# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22518 a_51294_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22519 a_41654_71552# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2252 VDD vcm.sky130_fd_sc_hd__buf_4_3.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+11p ps=4.74e+06u w=500000u l=500000u M=2
X22520 a_33526_23914# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22521 VDD a_1586_8439# a_3063_14741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22522 a_4036_67477# a_1591_67503# a_4259_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22523 a_37638_61512# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22524 VDD a_1923_53055# a_1643_56597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22525 a_38906_32509# a_2007_25597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22526 a_27198_19532# a_18546_19530# a_27106_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22527 a_34226_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22528 a_6636_72105# a_6602_72007# a_6381_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22529 a_41162_61150# a_18162_61190# a_41254_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2253 a_15107_40183# a_15093_39638# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X22530 a_9195_58951# a_6927_30503# a_9369_58827# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22531 a_2847_16127# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22532 a_13501_65149# a_13457_64757# a_13335_65161# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22533 a_3325_36495# a_2847_36799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22534 a_24094_71190# a_18162_71230# a_24186_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22535 a_29510_62194# pmat.rowon_n[6] a_29114_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22536 a_2203_16201# a_1757_15829# a_2107_16201# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22537 VSS pmat.row_n[10] a_26498_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22538 a_23486_15882# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22539 a_30514_16886# nmat.rowon_n[7] a_30118_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2254 a_30210_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22540 VDD a_5043_37191# a_4127_37013# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22541 VSS a_2007_49770# a_1895_50308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22542 a_9797_9813# a_1717_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X22543 VSS a_38041_30485# a_37975_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22544 a_45670_70548# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22545 vcm a_18162_67214# a_31214_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22546 a_49286_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22547 cgen.dlycontrol2_in[0] a_1591_37039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22548 vcm a_18162_57174# a_27198_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22549 VSS a_2411_43301# a_9361_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2255 VSS a_30765_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22550 a_42562_69222# pmat.rowon_n[13] a_42166_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22551 a_39111_38825# a_39505_38780# a_22153_37179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X22552 VDD a_1781_9308# a_1725_9334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X22553 a_14335_16519# a_12447_16143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22554 a_31214_55126# a_18546_55168# a_31122_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22555 a_31614_59504# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22556 a_27502_14878# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22557 VDD a_32957_30287# a_33299_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22558 a_25190_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22559 a_4837_45519# a_2983_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2256 VSS pmat.row_n[12] a_51598_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22560 a_15477_31055# a_13479_26935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22561 a_2219_4943# a_1775_5059# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22562 a_7442_42479# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22563 a_36637_27497# a_24591_28327# nmat.col[17] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22564 VDD pmat.rowon_n[14] a_22086_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22565 a_39550_67214# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22566 a_4032_64391# a_4162_64561# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22567 VSS pmat.row_n[9] a_43566_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22568 VDD nmat.rowon_n[6] a_43170_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22569 a_41254_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2257 VDD a_3859_22655# a_3846_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22570 VSS a_25287_51157# pmat.col_n[5] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22571 a_3116_77117# a_2999_76922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22572 a_31469_40726# a_30913_39867# a_32035_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22573 VSS a_39045_37692# a_38737_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22574 a_4985_74895# a_4259_73807# a_4505_74005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22575 a_9655_74216# a_9581_73487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22576 VSS a_7313_74005# a_7247_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22577 VDD a_2007_76970# a_1823_77821# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22578 vcm a_18162_18528# a_26194_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22579 a_49590_59182# pmat.rowon_n[3] a_49194_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2258 a_20848_38341# a_19689_38053# a_20811_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X22580 a_20474_65206# pmat.rowon_n[9] a_20078_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22581 VSS pmat.row_n[0] a_46578_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22582 a_30210_16520# a_18546_16518# a_30118_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22583 VDD nmat.rowon_n[7] a_47186_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22584 a_44666_13476# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22585 a_33949_39867# a_33007_38771# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22586 VSS pmat.row_n[10] a_29510_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22587 VDD a_6612_65845# a_5267_65479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22588 a_33526_64202# pmat.rowon_n[8] a_33130_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22589 VDD nmat.rowon_n[4] a_34134_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2259 a_18176_36165# a_12585_37179# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X22590 a_38996_50959# _1154_.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22591 a_27598_23516# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22592 a_83094_10383# ANTENNA__1190__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22593 VDD a_8767_16055# a_8767_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22594 a_27198_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22595 a_10081_52299# a_4259_31375# a_9995_52299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X22596 VDD nmat.rowon_n[2] a_31122_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22597 VSS a_12375_42895# a_12481_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22598 VDD a_4259_73807# a_4509_62037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22599 a_34226_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X226 vcm a_18162_57174# a_49286_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2260 VSS pmat.row_n[2] a_39550_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22600 a_51598_62194# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22601 a_23486_56170# pmat.rowon_n[0] a_23090_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22602 VSS a_4124_18231# a_2467_18517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22603 a_34530_72234# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22604 VDD nmat.rowon_n[10] a_21082_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22605 a_38242_65166# a_18546_65208# a_38150_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22606 a_38642_69544# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22607 VDD a_21124_36391# a_21028_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22608 VDD a_2325_40821# a_2215_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22609 VDD pmat.rowon_n[11] a_42166_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2261 VDD a_10873_38517# a_10817_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X22610 a_28110_15922# a_18162_15516# a_28202_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22611 vcm a_18162_61190# a_48282_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22612 a_6133_60137# a_5497_62839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22613 a_32218_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22614 VSS a_16311_28327# a_26149_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22615 VDD a_7658_71543# a_12815_74581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22616 a_11872_14191# a_10957_14191# a_11525_14433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22617 a_25190_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22618 a_27502_55166# VSS a_27106_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22619 a_14816_46831# a_3615_71631# a_14336_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2262 a_9919_57863# a_7521_47081# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X22620 VDD pmat.rowon_n[7] a_13547_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22621 vcm a_18162_8488# a_32218_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22622 a_42562_22910# nmat.rowon_n[1] a_42166_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22623 a_39154_65166# pmat.row_n[9] a_39646_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22624 a_27001_30511# a_23933_32143# a_26899_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X22625 a_40158_60146# pmat.row_n[4] a_40650_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22626 a_11041_36596# a_12267_36694# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22627 VDD pmat.rowon_n[12] a_28110_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22628 VDD a_1586_8439# a_7939_7125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22629 a_6981_28879# a_6579_29199# a_6817_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X2263 a_7809_17705# a_4976_16091# a_7737_17705# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X22630 VSS config_2_in[15] a_1591_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22631 a_39550_20902# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22632 a_43451_29423# a_41949_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22633 a_47861_27497# a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22634 vcm a_18162_72234# a_29206_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22635 VDD pmat.rowon_n[1] a_49194_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22636 VSS pmat.row_n[15] a_37542_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22637 a_33222_70186# a_18546_70228# a_33130_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22638 a_3894_72399# a_3136_72515# a_3331_72373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22639 a_26102_22950# pmat.row_n[14] a_26594_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2264 a_36485_49007# a_33957_48437# a_22499_49783# VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X22640 vcm a_18162_22544# a_47278_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22641 a_1644_34293# a_1591_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22642 a_30118_71190# pmat.row_n[15] a_30610_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22643 a_29206_60146# a_18546_60188# a_29114_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22644 a_30610_20504# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22645 a_37987_32521# a_37637_32149# a_37892_32509# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X22646 a_7847_20719# a_8197_20871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22647 a_29606_64524# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22648 a_30210_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22649 a_51294_20536# a_18546_20534# a_51202_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2265 VSS a_11927_27399# a_17323_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X22650 a_15395_31375# a_11067_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22651 VDD a_2046_30184# a_2051_29973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22652 VDD pmat.rowon_n[6] a_33130_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22653 a_47278_10496# a_18546_10494# a_47186_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22654 a_14565_63695# a_11067_64015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22655 a_19470_23914# pmat.rowoff_n[15] a_19074_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22656 a_14289_4649# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22657 a_9395_27791# a_8951_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22658 a_20570_12472# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22659 a_49590_12870# pmat.rowoff_n[4] a_49194_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2266 VSS a_37731_44527# pmat.sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X22660 a_7180_37039# a_6265_37039# a_6833_37281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22661 a_2107_64073# a_1591_63701# a_2012_64061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X22662 a_19566_56492# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22663 a_14486_46831# a_11067_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22664 a_42791_32375# a_44082_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22665 a_24186_22544# a_18546_22542# a_24094_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22666 VDD a_78802_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_1.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22667 VDD a_9020_7497# a_9195_7423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22668 a_33084_40743# a_31925_40955# a_33047_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22669 a_34134_70186# pmat.row_n[14] a_34626_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2267 a_23179_47753# a_22733_47381# a_23083_47753# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X22670 VDD a_3325_20175# a_9109_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22671 a_42166_18934# pmat.row_n[10] a_42658_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22672 VSS VDD a_42562_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22673 a_31122_12910# a_18162_12504# a_31214_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22674 a_39246_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22675 VSS a_4383_7093# a_8031_13353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22676 VSS pmat.row_n[13] a_31518_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22677 a_12267_36694# a_12309_36483# a_12267_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22678 a_2215_38671# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22679 a_32305_51335# a_28915_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2268 VDD pmat.rowoff_n[7] a_29114_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22680 VSS a_28245_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22681 a_1644_62581# a_1591_61519# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22682 VDD a_24867_53135# a_42065_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22683 VSS a_38727_32447# a_38661_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22684 a_35534_60186# pmat.rowon_n[4] a_35138_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22685 VSS a_36946_34191# a_37823_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22686 a_35534_19898# nmat.rowon_n[4] a_35138_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22687 a_23700_44869# a_22541_44581# a_23663_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22688 a_32218_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22689 a_28202_21540# a_18546_21538# a_28110_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2269 VDD a_8907_48437# a_8267_49159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X22690 a_25393_35877# a_24937_36039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X22691 a_46274_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22692 a_10593_15823# a_10423_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22693 a_19491_47893# a_19647_48052# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X22694 a_48586_18894# nmat.rowon_n[5] a_48190_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22695 a_39550_9858# nmat.rowon_n[14] a_39154_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22696 a_11104_71855# a_9375_72007# a_11014_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X22697 a_51598_9858# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22698 a_40250_68178# a_18546_68220# a_40158_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22699 a_32522_65206# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X227 VDD a_11115_71285# a_11322_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X2270 a_26594_12472# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22700 a_36234_58138# a_18546_58180# a_36142_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22701 a_32618_17492# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22702 vcm a_18162_69222# a_49286_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22703 a_30118_18934# a_18162_18528# a_30210_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22704 vcm a_18162_64202# a_50290_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22705 a_46182_19938# pmat.row_n[11] a_46674_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22706 a_29187_27791# a_21739_29415# a_28969_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22707 a_37975_30511# a_37827_30793# a_37612_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X22708 a_50198_68178# pmat.row_n[12] a_50690_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22709 a_49286_57134# a_18546_57176# a_49194_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2271 VSS a_19049_41959# a_17154_43671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22710 a_21124_39655# a_19965_39867# a_21087_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22711 a_2861_76757# a_2695_76757# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22712 VSS a_7405_32441# a_7339_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22713 a_22482_57174# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22714 a_78448_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_1.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22715 VSS pmat.row_n[6] a_49590_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22716 a_14923_34473# a_13801_34427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22717 VSS a_22449_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22718 a_2769_22357# a_2603_22357# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22719 a_39826_48829# a_2263_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2272 a_2672_20553# a_1591_20181# a_2325_20149# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X22720 a_35534_56170# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22721 VDD a_4516_21531# a_9595_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22722 a_22459_28879# a_22015_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22723 VSS a_16800_47213# a_16552_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22724 VSS a_10932_21959# a_10814_29111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X22725 a_26194_69182# a_18546_69224# a_26102_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22726 vcm a_18162_66210# a_23182_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22727 a_33130_13914# pmat.row_n[5] a_33622_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22728 VDD a_14465_29575# a_14471_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22729 a_9282_73853# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2273 a_24094_13914# a_18162_13508# a_24186_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22730 a_23582_19500# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22731 VDD a_15435_29111# a_15393_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22732 a_2507_29673# a_2648_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22733 VDD a_42240_29423# a_43451_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22734 a_21395_50857# a_22199_49667# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22735 a_33327_52521# _1184_.A2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22736 a_26498_14878# nmat.rowon_n[9] a_26102_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22737 a_36634_8456# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22738 VDD a_2244_20871# cgen.dlycontrol4_in[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22739 a_41558_23914# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2274 VDD nmat.rowon_n[13] a_30118_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22740 a_3207_65845# a_3410_66003# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22741 a_35230_19532# a_18546_19530# a_35138_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22742 vcm a_18162_65206# a_27198_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22743 VSS pmat.row_n[0] a_42562_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22744 VDD nmat.rowon_n[15] a_46182_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22745 a_27106_69182# pmat.row_n[13] a_27598_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22746 a_38546_67214# pmat.rowon_n[11] a_38150_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22747 a_31214_63158# a_18546_63200# a_31122_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22748 a_48282_18528# a_18546_18526# a_48190_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22749 a_31614_67536# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2275 VDD pmat.en_bit_n[2] nmat.en_bit_n[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X22750 vcm a_18162_15516# a_45270_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22751 VDD a_2879_60975# a_2727_58470# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22752 a_31122_57134# a_18162_57174# a_31214_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22753 VSS a_37612_30663# a_37143_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22754 pmat.col[21] a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22755 a_34134_8894# pmat.row_n[0] a_34626_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22756 VSS a_7373_49007# a_8309_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X22757 VSS a_3909_17209# a_3843_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22758 a_20811_44535# a_19689_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22759 a_4985_51433# a_4351_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X2276 a_8305_20871# a_12047_14165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X22760 a_10491_51183# a_9463_50877# a_10395_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22761 a_28506_8854# nmat.rowon_n[15] a_28110_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22762 VSS pmat.row_n[14] a_31518_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22763 a_28202_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22764 a_40554_70226# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22765 VSS ANTENNA__1395__B1.DIODE a_46934_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22766 pmat.col_n[31] _1196_.B1 a_46217_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22767 VDD a_4553_28089# a_4583_27830# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22768 a_22178_15516# a_18546_15514# a_22086_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22769 vcm a_18162_14512# a_49286_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2277 VSS a_14887_46377# a_14699_46377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22770 a_7210_11510# a_2021_9563# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X22771 a_9421_28335# a_4339_27804# a_9339_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22772 a_24937_43655# a_25209_44581# a_26272_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22773 a_24490_17890# nmat.rowon_n[6] a_24094_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22774 a_25393_41317# a_24937_41479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22775 a_12463_22351# a_12212_22467# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X22776 a_3970_55311# a_1823_58237# a_3884_55311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22777 a_22086_55126# VDD a_22578_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22778 a_43566_61190# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22779 VSS a_43533_30761# a_44801_35773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2278 a_44174_63158# pmat.row_n[7] a_44666_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22780 a_30210_24552# a_18546_24550# a_30118_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22781 a_50594_62194# pmat.rowon_n[6] a_50198_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22782 a_14466_28879# a_14287_28995# a_14466_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X22783 a_26194_14512# a_18546_14510# a_26102_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22784 vcm a_18162_11500# a_23182_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22785 a_19605_32149# a_19439_32149# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22786 a_25190_56130# a_18546_56172# a_25098_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22787 a_33526_72234# VDD a_33130_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22788 VSS pmat.row_n[5] a_25494_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22789 a_22482_10862# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2279 vcm a_18162_7484# a_49286_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22790 VDD _1154_.X a_36637_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22791 a_15757_52535# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22792 a_14618_72765# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22793 a_47582_60186# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22794 a_11019_71543# a_10975_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22795 a_13181_54447# a_13139_54599# a_13091_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X22796 a_47582_19898# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22797 VSS a_5687_71829# a_6772_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22798 a_5508_32687# a_5391_32900# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22799 a_35630_23516# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X228 a_7803_67655# a_7899_67477# a_8201_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X2280 a_48190_18934# pmat.row_n[10] a_48682_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22800 a_35230_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22801 a_28110_23954# a_18162_23548# a_28202_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22802 VDD pmat.rowon_n[9] a_38150_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22803 a_19233_41479# a_18953_43493# a_20016_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22804 VDD a_2727_58470# a_2969_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22805 a_48682_22512# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22806 a_9983_32385# a_2046_30184# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22807 a_12227_58633# a_11877_58261# a_12132_58621# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22808 VDD a_4135_19391# a_4122_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22809 a_11225_35836# a_11071_36694# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2281 VDD a_13091_52047# a_17459_49641# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22810 a_38242_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22811 a_27502_63198# pmat.rowon_n[7] a_27106_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22812 VDD a_18241_31698# a_18243_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22813 a_22086_72194# a_18162_72234# a_22178_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22814 a_10521_60975# a_10190_60663# a_10449_60975# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22815 VSS pmat.row_n[4] a_24490_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22816 a_20855_36885# a_20605_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22817 VSS pmat.row_n[11] a_24490_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22818 a_46481_52271# _1194_.B1 a_46263_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22819 a_35138_71190# a_18162_71230# a_35230_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2282 a_42258_69182# a_18546_69224# a_42166_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22820 a_38642_14480# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22821 a_38546_20902# pmat.rowoff_n[12] a_38150_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22822 VSS a_14641_57711# a_14839_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22823 a_36142_15922# a_18162_15516# a_36234_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22824 VDD pmat.rowoff_n[4] a_42166_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22825 a_10921_64786# a_14289_66421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X22826 a_40250_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22827 VSS a_1586_50247# a_1683_45205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22828 VSS a_12197_41570# a_11261_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X22829 VSS _1184_.A2 a_83166_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2283 a_13605_71017# a_13203_70767# a_13441_70767# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X22830 VDD nmat.rowon_n[1] a_25098_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22831 vcm a_18162_58178# a_25190_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22832 a_49194_14918# a_18162_14512# a_49286_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22833 VDD a_10676_30511# a_10851_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22834 VSS a_2007_8916# a_1895_8378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22835 a_35621_27247# a_26891_28327# nmat.col[16] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22836 VSS a_35244_32411# a_46723_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22837 a_8013_56085# a_7847_56085# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22838 VDD a_31152_48071# a_30687_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22839 VDD a_9528_20407# _0467_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2284 VDD a_4031_32852# a_3091_33402# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22840 a_40532_38341# a_39469_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22841 VDD a_25473_52245# pmat.col[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22842 a_39154_10902# pmat.row_n[2] a_39646_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22843 a_9231_32117# a_9666_32275# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22844 a_2163_56765# a_1586_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22845 a_38907_48841# a_38557_48469# a_38812_48829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22846 a_29606_72556# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22847 a_37542_68218# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22848 a_30210_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22849 a_12219_63303# a_11883_62063# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2285 a_20983_37277# a_20605_40719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X22850 VDD nmat.rowon_n[2] a_29114_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22851 VDD pmat.rowon_n[14] a_33130_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22852 a_26194_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22853 a_23090_11906# a_18162_11500# a_23182_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22854 a_2215_20175# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22855 VDD nmat.rowon_n[5] a_41162_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22856 a_29114_62154# a_18162_62194# a_29206_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22857 VDD a_31675_47695# a_43349_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22858 a_33222_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22859 a_11071_36694# a_11113_36483# a_11071_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 a_22111_36950# a_22153_37179# a_22111_37277# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22860 VSS a_39469_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22861 VSS a_28705_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22862 pmat.rowoff_n[13] a_14839_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X22863 VDD ANTENNA__1196__A2.DIODE a_13185_2473# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22864 VDD nmat.rowon_n[10] a_19074_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22865 VDD a_11007_58229# a_11257_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22866 vcm a_18162_19532# a_24186_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22867 a_31122_20942# a_18162_20536# a_31214_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22868 VSS a_19399_48437# a_16800_47213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X22869 a_42166_69182# a_18162_69222# a_42258_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2287 a_2405_29967# a_2237_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=0p ps=0u w=840000u l=150000u
X22870 VSS pmat.row_n[1] a_44570_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22871 a_33765_36965# a_33007_37683# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22872 a_38150_16926# pmat.row_n[8] a_38642_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22873 a_28525_43655# a_27785_43131# a_28907_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22874 VSS a_12076_62839# a_12081_62723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22875 a_45545_33551# a_40951_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22876 a_43170_9898# pmat.row_n[1] a_43662_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22877 VSS pmat.row_n[11] a_27502_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22878 VSS a_5123_52423# a_4866_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22879 VSS a_39647_48767# a_39581_48841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2288 vcm a_18162_71230# a_21174_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22880 a_31518_65206# pmat.rowon_n[9] a_31122_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22881 a_1586_18231# a_3944_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X22882 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22883 VSS a_9103_73791# a_9037_73865# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22884 a_19074_9898# pmat.row_n[1] a_19566_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22885 VSS a_28049_50613# pmat.col_n[8] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22886 VDD nmat.rowon_n[4] a_45178_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22887 a_4031_37191# a_4127_37013# a_4429_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22888 a_1881_56623# a_1846_56875# a_1643_56597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22889 VDD clk_ena a_25090_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2289 a_4523_21276# a_5179_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X22890 vcm a_18162_7484# a_21174_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22891 a_21478_57174# pmat.rowon_n[1] a_21082_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22892 a_46182_68178# a_18162_68218# a_46274_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22893 a_5989_40303# a_5823_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22894 a_29606_9460# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22895 VDD pmat.rowon_n[7] a_27106_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22896 a_2012_36861# a_1895_36666# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22897 a_31214_7484# a_18546_7482# a_31122_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22898 vcm a_18162_72234# a_50290_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22899 a_16197_40517# a_16505_40157# a_16171_40157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X229 a_23182_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2290 a_39246_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22900 a_49286_65166# a_18546_65208# a_49194_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22901 a_49686_69544# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22902 VDD config_2_in[13] a_2235_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22903 a_13549_74549# a_13331_74953# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22904 a_40250_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22905 a_41878_29673# a_41443_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22906 a_49194_59142# a_18162_59182# a_49286_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22907 a_23182_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22908 a_40650_17492# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22909 a_40554_23914# pmat.rowoff_n[15] a_40158_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2291 a_13683_24847# a_13367_24527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.73e+11p pd=2.98e+06u as=0p ps=0u w=420000u l=150000u
X22910 a_46921_30761# a_30571_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22911 a_44449_31029# a_43533_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22912 a_4069_19465# a_2879_19093# a_3960_19465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22913 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22914 a_20078_24958# nmat.en_C0_n a_20570_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22915 a_15543_31573# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22916 a_8378_12691# a_8656_12675# a_8612_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22917 VSS a_11202_55687# a_12175_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22918 VDD pmat.rowon_n[13] a_26102_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22919 a_51202_21946# pmat.row_n[13] a_51694_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2292 a_3399_33609# a_2953_33237# a_3303_33609# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X22920 a_51202_17930# a_18162_17524# a_51294_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22921 VSS a_44791_43541# a_44739_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22922 VSS a_30571_50959# a_36373_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22923 a_26194_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22924 a_23090_56130# a_18162_56170# a_23182_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22925 a_26437_27791# a_16311_28327# nmat.col_n[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22926 a_37542_21906# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22927 VSS a_23329_37462# a_22393_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X22928 a_40628_39429# a_39469_39141# a_40532_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22929 VDD a_40349_40726# a_39413_40956# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X2293 VDD a_43720_32143# a_46936_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X22930 VDD a_11797_60431# a_12219_63303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22931 a_41162_13914# pmat.row_n[5] a_41654_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22932 a_3215_22729# a_2769_22357# a_3119_22729# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22933 a_26498_66210# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22934 a_3859_56311# a_3967_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22935 a_34425_50959# a_30571_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X22936 VSS pmat.row_n[8] a_30514_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22937 VDD a_3859_56311# a_3225_55509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X22938 a_44666_55488# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22939 a_24094_23954# pmat.row_n[15] a_24586_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2294 VDD pmat.rowon_n[10] a_24094_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22940 a_24094_19938# a_18162_19532# a_24186_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22941 vcm a_18162_23548# a_45270_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22942 a_11057_67503# a_5363_70543# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22943 VSS a_31596_34191# a_31702_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22944 VSS a_16837_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22945 VSS a_12967_12863# a_12901_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X22946 a_27598_65528# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22947 a_2215_26525# a_1591_26159# a_2107_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22948 a_20337_41831# a_20645_42044# a_14149_39747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X22949 a_31122_65166# a_18162_65206# a_31214_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2295 a_21574_63520# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22950 a_6883_55862# a_5682_56311# a_6424_55687# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22951 a_34530_14878# nmat.rowon_n[9] a_34134_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22952 a_2500_30345# a_2051_29973# a_2405_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X22953 a_8397_71285# a_8179_71689# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22954 a_27106_55126# a_18162_55166# a_27198_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22955 VSS a_47592_35643# a_47591_35407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22956 VSS pmat.row_n[0] a_20474_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22957 a_47582_13874# nmat.rowon_n[10] a_47186_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22958 a_4031_32852# a_4123_32661# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X22959 VSS pmat.row_n[2] a_44570_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2296 a_4491_26486# a_2952_25045# a_4032_26311# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X22960 a_17996_36391# a_16837_36603# a_17959_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22961 a_5352_65577# a_5267_65479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22962 VSS a_6787_47607# a_7111_74575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22963 VDD VSS a_21082_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22964 a_27106_14918# pmat.row_n[6] a_27598_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22965 VSS pmat.row_n[12] a_27502_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22966 VSS a_14439_72703# a_14373_72777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X22967 a_16679_51183# a_13091_52047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22968 VDD a_7840_27247# a_19439_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22969 a_22178_23548# a_18546_23546# a_22086_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2297 a_31518_59182# pmat.rowon_n[3] a_31122_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22970 a_3727_66113# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22971 a_31614_12472# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22972 VSS a_8305_20871# a_9749_19061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22973 a_6400_60137# a_5731_58951# a_5939_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X22974 VSS pmat.row_n[0] a_50594_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22975 a_48190_7890# VDD a_48682_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22976 a_12543_40214# a_12585_40443# a_12543_40541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22977 VSS a_11409_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X22978 a_21478_10862# nmat.rowon_n[13] a_21082_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22979 a_21341_28585# a_10223_26703# a_21269_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2298 VDD a_11921_41814# a_10985_42044# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X22980 a_27167_31375# a_15101_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22981 VSS a_20695_30485# a_20629_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22982 a_44266_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22983 a_46578_60186# pmat.rowon_n[4] a_46182_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22984 a_22871_29967# a_22459_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X22985 a_25190_64162# a_18546_64204# a_25098_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22986 vcm a_18162_61190# a_22178_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22987 a_46578_19898# nmat.rowon_n[4] a_46182_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22988 a_9931_15279# a_9485_15279# a_9835_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22989 a_25590_68540# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2299 a_46274_68178# a_18546_68220# a_46182_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22990 a_15325_32509# a_10055_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22991 VDD a_7779_22583# a_7729_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22992 a_38552_32521# a_37471_32149# a_38205_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22993 VSS clk_ena a_31235_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22994 a_51294_68178# a_18546_68220# a_51202_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22995 a_13801_38779# a_10927_37981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X22996 a_8443_20719# a_7935_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.35e+11p pd=2.67e+06u as=0p ps=0u w=1e+06u l=150000u
X22997 a_47278_58138# a_18546_58180# a_47186_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22998 VDD a_1957_43567# a_12124_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22999 a_20474_58178# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_26498_18894# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X230 a_49286_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2300 vcm a_18162_65206# a_43262_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23000 a_28020_37479# a_26957_37691# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23001 vcm a_18162_60186# a_26194_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23002 a_4450_21629# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23003 a_26102_64162# pmat.row_n[8] a_26594_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23004 a_2250_61519# a_2124_61635# a_1846_61651# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23005 a_33526_57174# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23006 VDD VDD a_35138_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23007 a_30610_62516# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23008 vcm a_18162_10496# a_44266_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23009 a_3026_33775# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2301 a_43170_69182# pmat.row_n[13] a_43662_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23010 a_3151_48285# a_2971_48285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23011 VDD a_77528_39738# a_77341_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23012 a_38242_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23013 a_2012_26159# a_1895_26372# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23014 a_41558_7850# VDD a_41162_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23015 a_1895_38842# a_1899_35051# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23016 a_3325_40847# a_2847_41151# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23017 a_20682_30877# a_19605_30511# a_20520_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23018 VSS a_2199_13887# a_8413_12925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23019 a_34626_19500# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2302 a_5245_56053# a_2407_49289# a_5498_56399# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X23020 vcm a_18162_22544# a_21174_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23021 a_17021_38053# a_13503_37981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X23022 a_36142_23954# a_18162_23548# a_36234_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23023 a_33622_7452# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23024 a_21174_10496# a_18546_10494# a_21082_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23025 VDD nmat.rowon_n[13] a_38150_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23026 VSS a_6853_55509# a_6787_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23027 VSS pmat.row_n[1] a_22482_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23028 a_49194_22950# a_18162_22544# a_49286_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23029 a_36538_68218# pmat.rowon_n[12] a_36142_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2303 a_3668_6397# a_3551_6202# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X23030 a_11795_64899# a_10569_64489# a_11713_64899# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23031 a_46274_19532# a_18546_19530# a_46182_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23032 vcm a_18162_16520# a_43262_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23033 a_3986_74575# a_3267_74817# a_3423_74549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23034 a_7068_11703# a_7283_11484# a_7210_11510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23035 VDD a_2315_44124# a_3151_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23036 VSS a_20475_49783# a_20175_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23037 a_42562_15882# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23038 VSS pmat.row_n[10] a_45574_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23039 a_44733_44431# a_7109_29423# a_44745_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2304 a_46182_9898# pmat.row_n[1] a_46674_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23040 VDD a_1643_54965# a_1591_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23041 a_11030_30511# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23042 VDD a_8908_14967# a_8767_16055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23043 a_26194_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23044 a_46636_36469# a_38851_28327# a_47293_36815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23045 a_27443_32143# a_24374_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X23046 a_47685_30517# a_35244_32411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23047 vcm a_18162_57174# a_46274_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23048 VDD a_2683_22089# a_7819_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23049 a_39826_47741# a_2263_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2305 a_2468_21959# a_1781_9308# a_2610_21807# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23050 a_47915_46506# a_47975_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23051 a_20170_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23052 a_19166_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23053 a_50690_59504# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23054 a_22482_18894# nmat.rowon_n[5] a_22086_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23055 a_46578_14878# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23056 a_14107_39958# a_14149_39747# a_14107_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23057 a_29510_24918# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23058 VSS a_21970_48071# a_21923_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X23059 VSS a_12213_53359# a_12895_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2306 VDD a_22537_36911# a_40399_36911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23060 VDD a_3751_64757# a_2944_65576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X23061 vcm a_18162_9492# a_37238_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23062 VSS a_2411_16101# a_2369_20541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23063 a_38150_67174# a_18162_67214# a_38242_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23064 VDD pmat.rowon_n[4] a_37146_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23065 vcm a_18162_59182# a_19166_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23066 a_33130_55126# VDD a_33622_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23067 a_23182_57134# a_18546_57176# a_23090_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23068 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23069 a_20078_58138# pmat.row_n[2] a_20570_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2307 VSS a_77980_38962# vcm.sky130_fd_sc_hd__buf_4_3.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X23070 a_47278_9492# a_18546_9490# a_47186_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23071 a_19470_16886# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23072 VSS pmat.row_n[6] a_23486_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23073 a_20474_11866# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23074 a_42658_24520# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23075 VSS a_22787_34709# a_12197_38306# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23076 a_33526_10862# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23077 a_2163_71997# a_1674_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23078 VSS pmat.row_n[11] a_35534_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23079 VDD pmat.rowon_n[15] a_27106_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2308 a_35269_49257# a_25695_28111# nmat.col[15] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X23080 a_5183_67503# a_5307_67655# a_5046_67655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23081 a_83741_26409# ANTENNA__1395__B1.DIODE nmat.col_n[29] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23082 VSS pmat.row_n[10] a_48586_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23083 a_10897_6825# a_10378_7637# a_9459_5461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23084 VDD a_25287_51157# pmat.col_n[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X23085 a_5603_18543# a_5087_18543# a_5508_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23086 VDD nmat.rowon_n[14] a_39154_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23087 a_43170_20942# pmat.row_n[12] a_43662_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23088 a_46674_23516# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23089 a_46274_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2309 a_28506_57174# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23090 a_43170_16926# a_18162_16520# a_43262_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23091 a_51202_9898# pmat.row_n[1] a_51694_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23092 VDD nmat.rowon_n[2] a_50198_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23093 a_50198_62154# a_18162_62194# a_50290_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23094 a_18891_47491# a_18547_51565# a_18795_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23095 a_38793_49007# a_38515_49035# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X23096 a_49286_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23097 a_12481_36694# a_12309_36483# a_12267_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23098 a_42562_56170# pmat.rowon_n[0] a_42166_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23099 VDD nmat.rowon_n[5] a_39154_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X231 a_25494_18894# nmat.rowon_n[5] a_25098_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2310 a_25590_62516# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23100 a_33130_72194# a_18162_72234# a_33222_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23101 a_36634_15484# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23102 a_36538_21906# nmat.rowon_n[2] a_36142_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23103 a_14058_74575# a_12981_74581# a_13896_74953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23104 VDD nmat.rowon_n[10] a_40158_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23105 VDD a_6412_8725# a_6548_8751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.184e+11p ps=2.2e+06u w=840000u l=150000u
X23106 a_25494_66210# pmat.rowon_n[10] a_25098_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23107 a_49686_14480# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23108 VDD pmat.rowoff_n[15] a_23090_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23109 a_17959_36649# a_16837_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2311 vcm a_18162_10496# a_39246_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23110 a_19834_34191# a_19657_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23111 a_47186_15922# a_18162_15516# a_47278_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23112 a_23090_64162# a_18162_64202# a_23182_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23113 a_51294_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23114 a_11216_17455# a_9441_20189# a_10995_17782# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X23115 a_1823_64213# a_2847_63999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23116 a_4785_38377# a_3325_36495# a_4713_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23117 a_14287_60975# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23118 a_2203_43401# a_1757_43029# a_2107_43401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23119 VSS a_14839_66103# a_14839_65871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2312 a_49590_71230# pmat.rowon_n[15] a_49194_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23120 pmat.rowoff_n[10] a_11067_64015# a_14830_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23121 a_2939_45503# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23122 a_37146_11906# pmat.row_n[3] a_37638_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23123 VSS VDD a_30514_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23124 VSS a_45119_32661# a_45077_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23125 a_29510_65206# pmat.rowon_n[9] a_29114_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23126 a_2107_33775# a_1591_33775# a_2012_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23127 VDD pmat.rowon_n[13] a_34134_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23128 a_37146_9898# a_18162_9492# a_37238_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23129 VDD a_11202_55687# a_13289_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2313 a_30118_67174# a_18162_67214# a_30210_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23130 VDD nmat.rowon_n[9] a_26102_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23131 VSS a_3571_13627# a_11619_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23132 a_4415_71631# a_1823_76181# a_4225_71311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23133 a_24186_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23134 a_20752_41605# a_19689_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23135 a_44266_61150# a_18546_61192# a_44174_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23136 a_11159_23145# a_6173_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23137 a_5821_32929# a_5603_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23138 VSS a_35186_47375# a_37519_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23139 VDD pmat.rowon_n[12] a_47186_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2314 VSS VDD a_32522_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23140 a_27106_63158# a_18162_63198# a_27198_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23141 a_48586_68218# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23142 a_16163_43413# a_16339_43745# a_16291_43805# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23143 a_47278_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23144 a_9485_15279# a_9319_15279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23145 a_19470_57174# pmat.rowon_n[1] a_19074_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23146 a_4687_28335# a_4241_28335# a_4591_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23147 VDD config_1_in[11] a_1626_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23148 a_11265_47919# a_11230_48171# a_10795_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23149 a_23884_40517# a_22725_40229# a_23847_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X2315 VDD a_19928_37253# a_19832_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X23150 a_3026_18365# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23151 a_35630_65528# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23152 a_27598_10464# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23153 a_28946_30287# a_28715_28879# a_27995_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23154 VSS pmat.row_n[2] a_42562_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23155 VDD a_2163_69821# a_2124_69947# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23156 pmat.rowon_n[12] a_14839_65871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23157 a_48282_60146# a_18546_60188# a_48190_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23158 a_7093_13353# a_5579_12394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X23159 a_48682_64524# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2316 a_41254_9492# a_18546_9490# a_41162_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23160 a_45178_61150# pmat.row_n[5] a_45670_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23161 a_21478_60186# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23162 VSS a_4956_59317# a_3956_59317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X23163 vcm a_18162_19532# a_35230_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23164 a_21478_19898# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23165 VSS a_2847_33749# a_2781_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23166 VSS a_9963_13967# nmat.rowoff_n[11] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23167 a_35717_28111# ANTENNA__1197__A.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23168 a_5989_34863# a_5823_34863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23169 a_15690_31375# a_15660_31029# a_15395_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2317 a_19605_30511# a_19439_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23170 a_34611_43177# a_33489_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23171 VSS pmat.row_n[12] a_35534_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23172 a_34530_18894# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23173 VDD a_13091_28327# a_35729_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23174 a_25190_72194# a_18546_72236# a_25098_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23175 a_38642_56492# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23176 VDD a_7907_52031# a_7894_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23177 a_23420_43781# a_22357_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23178 a_11205_77295# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23179 a_43262_22544# a_18546_22542# a_43170_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2318 a_18546_58180# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X23180 VDD pmat.rowon_n[8] a_25098_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23181 a_39246_12504# a_18546_12502# a_39154_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23182 a_22578_61512# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23183 a_49194_60146# pmat.row_n[4] a_49686_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23184 VSS pmat.row_n[13] a_50594_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23185 a_12092_42895# a_11915_42895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23186 a_26102_72194# VDD a_26594_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23187 a_6170_5739# a_6448_5755# a_6404_5853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23188 VSS a_39469_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23189 a_37542_70226# pmat.rowon_n[14] a_37146_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2319 a_6837_10499# a_2021_11043# a_6742_10499# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X23190 a_11071_40719# a_10817_41046# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23191 a_30610_70548# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23192 a_51294_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23193 a_45574_9858# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23194 a_26594_60508# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23195 VSS a_10873_40693# a_26459_42657# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23196 a_34226_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23197 VDD a_17559_51157# pmat.rowoff_n[15] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X23198 a_51598_65206# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23199 VSS a_33765_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X232 a_23604_36391# a_23700_36391# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X2320 a_3983_47919# a_4075_50087# a_4071_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23200 a_51694_17492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23201 a_51598_23914# pmat.rowoff_n[15] a_51202_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23202 VDD VSS a_19074_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23203 VSS a_39647_47679# a_39581_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X23204 VSS pmat.row_n[9] a_37542_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23205 VSS a_15101_29423# a_25352_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23206 a_41558_57174# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23207 a_11731_8751# a_11051_8903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23208 a_41558_15882# pmat.rowoff_n[7] a_41162_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23209 a_24490_67214# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2321 a_23763_27497# a_10883_3303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X23210 VDD a_33386_30485# a_31675_47695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X23211 VDD a_14439_72703# a_14426_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23212 a_48586_21906# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23213 VSS a_21621_35515# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23214 vcm a_18162_24552# a_43262_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23215 a_23846_27247# _1192_.B1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23216 a_45270_69182# a_18546_69224# a_45178_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23217 a_19470_10862# nmat.rowon_n[13] a_19074_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23218 vcm a_18162_66210# a_42258_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23219 a_41949_30761# a_38905_28853# a_41795_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2322 VSS ANTENNA__1395__A2.DIODE a_27616_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X23220 a_2629_53181# a_2250_52815# a_2557_53181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23221 vcm a_18162_56170# a_38242_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23222 a_35138_23954# pmat.row_n[15] a_35630_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23223 a_35138_19938# a_18162_19532# a_35230_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23224 a_18176_42693# a_17113_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23225 VSS a_3866_57399# a_6829_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23226 VSS a_46817_43541# a_46582_46519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23227 a_14261_44219# a_13805_43990# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X23228 a_42658_58500# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23229 a_38546_13874# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2323 a_44266_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23230 a_3026_50095# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23231 a_45574_14878# nmat.rowon_n[9] a_45178_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23232 VSS pmat.row_n[3] a_42562_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23233 a_17459_37143# a_17675_37001# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23234 a_39246_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23235 VSS pmat.row_n[0] a_31518_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23236 a_28602_18496# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23237 a_28506_24918# VSS a_28110_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23238 VDD a_2411_33749# a_10284_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23239 a_78802_39738# a_78898_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2324 a_7263_42453# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X23240 a_25098_15922# pmat.row_n[7] a_25590_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23241 a_38293_51727# a_24591_28327# pmat.col_n[18] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23242 VDD nmat.rowon_n[7] a_32126_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23243 vcm a_18162_65206# a_46274_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23244 a_39193_42043# a_38737_41814# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X23245 a_46182_69182# pmat.row_n[13] a_46674_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23246 a_50290_63158# a_18546_63200# a_50198_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23247 a_50690_67536# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23248 VSS a_13985_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23249 VSS pmat.row_n[1] a_30514_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2325 pmat.col_n[30] a_46934_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23250 a_28110_8894# pmat.row_n[0] a_28602_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23251 a_36175_50345# a_26891_28327# pmat.col_n[16] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X23252 a_22879_41781# a_23055_41781# a_23007_41807# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23253 VDD a_2407_49289# a_7377_65577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23254 a_1959_12791# a_1979_12342# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23255 vcm a_18162_67214# a_19166_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23256 a_41162_7890# a_18162_7484# a_41254_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23257 VSS config_2_in[5] a_1591_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X23258 a_23182_65166# a_18546_65208# a_23090_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23259 vcm a_18162_62194# a_20170_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 a_14803_31599# a_14453_31599# a_14708_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X23260 VSS pmat.row_n[14] a_50594_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23261 a_23582_69544# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23262 vcm a_18162_17524# a_37238_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23263 a_20078_66170# pmat.row_n[10] a_20570_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23264 a_19166_55126# a_18546_55168# a_19074_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23265 VSS a_28116_37479# a_28189_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X23266 a_33489_36603# a_30155_36893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X23267 a_39981_37462# a_39469_38053# a_40532_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23268 a_19566_59504# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23269 a_41254_15516# a_18546_15514# a_41162_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2327 VSS a_45282_32143# ANTENNA__1196__A2.DIODE VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u M=16
X23270 a_2672_41225# a_1757_40853# a_2325_40821# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23271 VSS a_13653_40956# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23272 vcm a_18162_61190# a_33222_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23273 a_51294_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23274 a_5715_16911# a_5463_17027# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X23275 a_24033_28111# a_13459_28111# a_23815_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23276 a_5260_67753# a_3866_57399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23277 VSS a_11261_37981# a_10953_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23278 a_12559_51325# a_5363_33551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23279 a_7521_31421# a_7477_31029# a_7355_31433# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2328 a_20078_59142# a_18162_59182# a_20170_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23280 a_41162_55126# VDD a_41654_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23281 cgen.dlycontrol2_in[4] a_2603_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23282 VDD config_2_in[11] a_1591_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23283 a_24094_65166# pmat.row_n[9] a_24586_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23284 a_17996_35303# a_16837_35515# a_17959_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X23285 a_11285_36694# a_11113_36483# a_11071_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23286 a_45270_14512# a_18546_14510# a_45178_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23287 vcm a_18162_11500# a_42258_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23288 a_45574_71230# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23289 VSS a_5081_53135# a_6334_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2329 a_29606_19500# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23290 a_43170_24958# a_18162_24552# a_43262_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23291 a_42709_27791# a_21739_29415# nmat.col_n[22] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23292 VDD a_3688_17179# a_10489_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23293 a_14647_51701# a_14452_51843# a_14957_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23294 a_11542_50461# a_11416_50363# a_11138_50347# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23295 a_41558_10862# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23296 a_2595_13621# a_2439_13889# a_2740_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23297 a_21478_8854# nmat.rowon_n[15] a_21082_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23298 a_11233_76207# a_11023_76359# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23299 a_24490_20902# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X233 VSS pmat.row_n[7] a_22482_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2330 a_30121_31599# a_28704_29568# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.46e+11p pd=5.58e+06u as=0p ps=0u w=650000u l=150000u
X23300 a_49286_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23301 a_1979_12342# a_1717_13647# a_1979_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23302 a_4446_65871# a_3688_65987# a_3883_65845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23303 a_7370_27791# a_7023_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X23304 a_27106_56130# pmat.row_n[0] a_27598_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23305 a_36234_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23306 a_12901_12937# a_11711_12565# a_12792_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23307 VSS pmat.row_n[15] a_22482_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23308 a_6242_70767# a_3339_70759# a_6432_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23309 a_11455_50237# a_5363_33551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2331 a_20170_20536# a_18546_20534# a_20078_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23310 a_49590_70226# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23311 VSS a_1923_61759# a_8413_64061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23312 VDD nmat.rowon_n[12] a_36142_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23313 vcm a_18162_22544# a_32218_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23314 a_2971_48285# a_2983_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23315 a_4591_14025# a_4241_13653# a_4496_14013# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23316 vcm a_18162_12504# a_28202_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23317 a_17054_28995# a_16863_29239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23318 VSS a_2847_18303# a_2781_18377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X23319 a_47186_23954# a_18162_23548# a_47278_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2332 a_40554_17890# nmat.rowon_n[6] a_40158_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23320 a_32218_10496# a_18546_10494# a_32126_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23321 VSS cgen.dlycontrol4_in[1] a_1945_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23322 vcm a_18162_59182# a_40250_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23323 VSS a_3325_43023# a_3983_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X23324 VSS a_5558_9527# a_5510_9615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23325 a_39550_62194# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23326 a_12875_16341# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23327 a_41162_72194# a_18162_72234# a_41254_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23328 VSS pmat.row_n[4] a_43566_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23329 a_14373_72777# a_13183_72405# a_14264_72777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2333 a_47582_23914# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23330 a_9502_53609# a_9463_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23331 VSS pmat.row_n[11] a_43566_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23332 a_40554_16886# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23333 VSS pmat.row_n[14] a_26498_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23334 VDD a_9103_56383# a_9090_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23335 VSS a_33957_48437# a_35306_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23336 a_33489_44219# a_32256_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X23337 a_45747_51433# a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23338 a_24186_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23339 a_44145_28363# a_38851_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2334 a_2467_35015# a_2563_34837# a_2865_34863# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23340 a_7302_34102# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23341 a_77528_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_2.X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23342 VDD a_1586_18231# a_1591_27797# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23343 a_36234_8488# a_18546_8486# a_36142_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23344 VDD nmat.rowon_n[1] a_44174_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23345 vcm a_18162_58178# a_44266_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23346 VSS a_3571_13627# a_4075_13653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23347 a_1881_31599# a_1846_31851# a_1643_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23348 a_20474_60186# pmat.rowon_n[4] a_20078_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23349 a_20474_19898# nmat.rowon_n[4] a_20078_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2335 a_44737_45199# a_29937_31055# a_44447_45431# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.4e+11p pd=2.88e+06u as=5.2e+11p ps=3.04e+06u w=1e+06u l=150000u
X23350 VSS pmat.row_n[5] a_29510_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23351 VDD a_1586_50247# a_6651_51733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23352 a_2325_26401# a_2107_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23353 a_31214_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23354 VDD nmat.rowon_n[9] a_34134_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23355 comp.adc_nor_latch_0.QN comp_latch a_56106_40254# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23356 a_33526_18894# nmat.rowon_n[5] a_33130_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23357 a_4579_47919# a_4071_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.35e+11p pd=2.67e+06u as=0p ps=0u w=1e+06u l=150000u
X23358 a_12691_31433# a_12245_31061# a_12595_31433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23359 vcm a_18162_8488# a_34226_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2336 a_51202_15922# pmat.row_n[7] a_51694_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23360 a_48682_72556# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23361 a_21174_58138# a_18546_58180# a_21082_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23362 vcm a_18162_69222# a_34226_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23363 a_45270_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23364 a_42166_11906# a_18162_11500# a_42258_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23365 VDD pmat.rowon_n[4] a_48190_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23366 a_31122_19938# pmat.row_n[11] a_31614_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23367 VDD a_4135_37815# a_2839_38101# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X23368 a_34226_57134# a_18546_57176# a_34134_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23369 pmat.rowon_n[2] a_11067_16359# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2337 VSS pmat.row_n[13] a_51598_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23370 VDD a_25688_32117# a_25287_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23371 VDD a_11067_27239# a_24118_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23372 a_2107_50095# a_1591_50095# a_2012_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23373 a_12629_68367# a_12597_68279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23374 a_35630_10464# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23375 VSS pmat.row_n[6] a_34530_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23376 a_28110_10902# a_18162_10496# a_28202_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23377 a_46896_44905# a_7109_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23378 VDD VDD a_25098_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23379 a_39246_20536# a_18546_20534# a_39154_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2338 a_39015_48463# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X23380 nmat.col_n[1] a_13354_2223# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23381 a_4682_6397# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23382 a_25190_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23383 VSS pmat.row_n[11] a_46578_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23384 a_43566_64202# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23385 VDD a_2215_47375# a_2879_60975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23386 VDD a_12069_36341# a_12481_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23387 a_50594_65206# pmat.rowon_n[9] a_50198_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23388 a_4491_47158# a_2315_44124# a_4032_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23389 VSS a_1586_63927# a_1591_63701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2339 vcm a_18162_16520# a_38242_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23390 a_1979_12342# a_1761_11471# a_1907_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X23391 VDD a_43533_30761# a_46765_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23392 VSS pmat.row_n[3] a_36538_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23393 a_19074_12910# a_18162_12504# a_19166_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23394 a_20170_19532# a_18546_19530# a_20078_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23395 a_40554_57174# pmat.rowon_n[1] a_40158_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23396 VDD a_31923_42367# a_31783_42689# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23397 a_18675_47081# a_18547_51565# a_18603_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23398 VSS pmat.row_n[13] a_19470_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23399 VSS a_2847_50069# a_2781_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X234 a_49590_14878# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2340 a_48282_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23400 a_23486_67214# pmat.rowon_n[11] a_23090_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23401 a_22541_36603# a_22085_36374# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X23402 vcm a_18162_15516# a_30210_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23403 a_33222_18528# a_18546_18526# a_33130_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23404 a_47678_15484# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23405 a_9274_76751# a_8197_76757# a_9112_77129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23406 a_2203_36873# a_1757_36501# a_2107_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23407 VDD nmat.rowon_n[10] a_51202_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23408 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23409 a_7072_62037# a_1823_68565# a_7295_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2341 VSS a_16607_36911# a_16713_36911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23410 a_2672_18377# a_1591_18005# a_2325_17973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23411 a_37542_55166# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23412 a_12162_39958# a_12116_39783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23413 a_2163_71997# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23414 a_25639_43957# a_25815_43957# a_25767_43983# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X23415 a_3315_69455# a_2727_58470# a_3219_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23416 vcm a_18162_14512# a_34226_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23417 a_48190_11906# pmat.row_n[3] a_48682_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23418 VSS a_9287_65087# a_9221_65161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23419 vcm a_18162_64202# a_38242_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2342 a_42258_14512# a_18546_14510# a_42166_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23420 VDD a_1643_71829# a_1591_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23421 a_47861_51727# ANTENNA__1395__B1.DIODE pmat.col[28] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23422 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=5.1e+06u w=1.89e+07u
X23423 a_38150_68178# pmat.row_n[12] a_38642_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23424 a_42258_62154# a_18546_62196# a_42166_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23425 VDD pmat.rowon_n[13] a_45178_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23426 a_42658_66532# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23427 a_46936_44111# a_7109_29423# a_46845_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23428 a_9037_56457# a_7847_56085# a_8928_56457# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23429 a_22578_9460# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2343 VSS a_10873_38517# a_10817_38870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23430 a_12249_71311# a_11893_71427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23431 a_45270_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23432 a_42166_56130# a_18162_56170# a_42258_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23433 VSS a_30699_29397# a_31072_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23434 a_7180_37039# a_6099_37039# a_6833_37281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23435 a_28202_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23436 a_25098_66170# a_18162_66210# a_25190_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23437 a_24719_39605# a_12228_39605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23438 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23439 VSS a_35244_32411# a_47499_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2344 a_41254_56130# a_18546_56172# a_41162_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23440 a_4403_51701# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X23441 VSS a_28189_37981# a_27881_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23442 a_19523_47491# a_12263_50959# a_19441_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23443 VSS a_1923_61759# a_8809_65149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23444 a_6179_69831# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23445 a_2398_51859# a_2676_51843# a_2632_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23446 a_46674_65528# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23447 a_43170_62154# pmat.row_n[6] a_43662_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23448 a_46182_55126# a_18162_55166# a_46274_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23449 a_17959_35561# a_16837_35515# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2345 VSS a_12449_22895# a_14301_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.24e+11p ps=5.82e+06u w=650000u l=150000u
X23450 a_32522_60186# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23451 a_32522_19898# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23452 vcm a_18162_70226# a_20170_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23453 a_36634_57496# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23454 a_38642_8456# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23455 a_19166_63158# a_18546_63200# a_19074_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23456 VDD VSS a_40158_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23457 a_46182_14918# pmat.row_n[6] a_46674_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23458 VSS pmat.row_n[12] a_46578_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23459 a_49590_23914# pmat.rowoff_n[15] a_49194_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2346 VSS a_33567_30199# a_32865_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23460 a_20570_23516# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23461 VDD a_1899_35051# a_1857_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23462 VSS a_12069_36341# a_12488_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23463 VSS comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.84e+07u l=3.9e+06u
X23464 a_19566_67536# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23465 a_20170_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23466 a_41254_23548# a_18546_23546# a_41162_23954# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23467 a_50690_12472# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23468 VDD pmat.rowon_n[9] a_23090_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23469 a_49686_56492# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2347 a_24094_58138# a_18162_58178# a_24186_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23470 a_37238_13508# a_18546_13506# a_37146_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23471 a_29114_24958# VDD a_29606_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23472 a_1979_12015# a_1725_12342# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23473 VSS pmat.row_n[0] a_44570_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23474 VDD nmat.rowon_n[15] a_48190_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23475 VSS a_40951_31599# a_45629_35773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23476 a_19074_57134# a_18162_57174# a_19166_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23477 a_33622_22512# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23478 a_23182_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23479 VSS a_3339_59879# a_13501_65149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2348 VSS a_5991_23983# a_10515_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X23480 a_39550_15882# pmat.rowoff_n[7] a_39154_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23481 VSS pmat.row_n[4] a_36538_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23482 a_13236_8573# a_12257_8527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23483 a_40554_10862# nmat.rowon_n[13] a_40158_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23484 VSS pmat.row_n[14] a_19470_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23485 a_9137_27253# a_4516_21531# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23486 a_23582_14480# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23487 a_23486_20902# pmat.rowoff_n[12] a_23090_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23488 a_46667_46287# a_29937_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23489 a_21082_15922# a_18162_15516# a_21174_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2349 a_37542_15882# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23490 VDD pmat.rowon_n[0] a_26102_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23491 vcm a_18162_61190# a_41254_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23492 VSS a_4679_28853# a_4379_28548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23493 a_48586_70226# pmat.rowon_n[14] a_48190_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23494 a_19233_40719# a_18963_41085# a_19143_41085# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23495 a_27249_28995# a_22459_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23496 a_34134_14918# a_18162_14512# a_34226_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23497 VDD a_5411_12167# a_5363_12015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23498 VSS a_34204_27765# a_37828_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23499 a_3229_14741# a_3063_14741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X235 VDD a_20329_35431# a_17675_37001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X2350 a_18546_23546# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X23500 a_38546_62194# pmat.rowon_n[6] a_38150_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23501 a_28867_40871# a_21981_34191# a_29041_40747# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23502 a_24094_10902# pmat.row_n[2] a_24586_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23503 a_22482_68218# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23504 vcm a_18162_20536# a_28202_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23505 VSS a_16800_47213# a_17187_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23506 a_6292_65479# a_12225_74575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23507 VSS a_11759_10615# a_11051_8903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23508 vcm a_18162_67214# a_40250_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23509 a_35534_67214# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2351 a_44570_16886# nmat.rowon_n[7] a_44174_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23510 VSS a_11067_16359# pmat.rowon_n[4] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23511 a_6346_65577# a_6292_65479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23512 a_19955_30511# a_19439_30511# a_19860_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23513 VDD a_19551_34191# a_19657_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23514 a_37146_70186# a_18162_70226# a_37238_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23515 a_2121_74031# a_1643_74005# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23516 VDD a_1586_8439# a_8399_6037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23517 a_5361_72399# a_5271_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23518 VSS a_2791_57703# a_4327_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23519 a_24131_29967# a_22628_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2352 VSS pmat.row_n[5] a_41558_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23520 a_27598_7452# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23521 a_23486_7850# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23522 a_2882_70045# a_2124_69947# a_2319_69916# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23523 a_25494_59182# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23524 vcm a_18162_12504# a_36234_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23525 a_9839_47679# a_9664_47753# a_10018_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23526 VDD config_1_in[6] a_1591_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23527 VDD a_10873_40693# a_10817_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X23528 a_40250_10496# a_18546_10494# a_40158_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23529 a_23090_16926# pmat.row_n[8] a_23582_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2353 a_24094_17930# pmat.row_n[9] a_24586_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23530 a_2099_24746# a_2191_24501# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23531 VDD nmat.rowon_n[4] a_30118_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23532 VSS a_10515_13967# a_20267_50345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23533 a_29510_58178# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23534 VSS a_34942_51701# a_35252_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23535 a_19405_28853# a_6664_26159# a_19526_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23536 a_31122_68178# a_18162_68218# a_31214_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23537 a_12245_21807# a_11897_21813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X23538 a_21082_8894# a_18162_8488# a_21174_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23539 VSS a_36854_44527# a_37731_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2354 VSS pmat.row_n[15] a_24490_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23540 a_7373_48695# a_6787_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23541 a_2882_74397# a_2163_74173# a_2319_74268# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23542 a_45270_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23543 a_39089_27765# a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23544 a_8397_71285# a_8179_71689# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23545 a_13729_10761# a_12539_10389# a_13620_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23546 a_34226_65166# a_18546_65208# a_34134_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23547 a_11167_11177# a_11207_11079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23548 a_31214_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23549 VDD a_13479_26935# a_14905_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2355 a_4634_32509# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X23550 a_34626_69544# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23551 vcm a_18162_17524# a_48282_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23552 VDD a_10873_36341# a_11285_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23553 a_12164_4175# _1194_.B1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23554 a_5749_57685# a_4351_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23555 a_34134_59142# a_18162_59182# a_34226_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23556 a_4450_21302# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23557 vcm a_18162_7484# a_48282_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23558 a_36209_49257# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X23559 a_25767_43983# a_11041_39860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2356 VSS a_33341_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23560 a_43566_72234# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23561 a_35138_65166# pmat.row_n[9] a_35630_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23562 a_39581_47753# a_38391_47381# a_39472_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23563 VDD a_13427_18303# a_13414_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23564 a_12949_18365# a_12905_17973# a_12783_18377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23565 VDD a_2655_59317# a_1823_60949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23566 a_36142_10902# a_18162_10496# a_36234_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23567 a_12245_31061# a_12079_31061# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23568 a_37739_42089# a_36617_42043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23569 VSS VDD a_25494_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2357 VDD a_6557_35105# a_6447_35229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X23570 a_22482_21906# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23571 a_19074_20942# a_18162_20536# a_19166_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23572 a_14460_12265# a_11435_58791# a_14369_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23573 a_25098_57134# pmat.row_n[1] a_25590_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23574 VDD a_22527_27221# nmat.col[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X23575 a_36538_55166# pmat.en_bit_n[0] a_36142_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23576 VSS vcm.sky130_fd_sc_hd__buf_4_3.A a_77980_38962# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23577 a_13203_70767# a_12809_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23578 a_30699_29397# a_21365_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23579 a_35534_20902# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2358 a_35715_29941# a_35559_30209# a_35860_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X23580 vcm a_18162_23548# a_30210_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23581 a_29206_16520# a_18546_16518# a_29114_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23582 a_47278_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23583 a_45178_9898# pmat.row_n[1] a_45670_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23584 a_30833_46805# a_31105_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X23585 a_76962_39738# a_77058_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23586 a_7160_33927# a_6007_33767# a_7302_34102# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23587 VSS pmat.row_n[7] a_28506_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23588 a_25494_12870# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23589 a_40785_29673# a_17842_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2359 VDD pmat.rowon_n[1] a_31122_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X23590 a_37542_63198# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23591 a_32035_36649# a_30913_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23592 a_32522_13874# nmat.rowon_n[10] a_32126_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23593 a_9583_10121# a_14071_8511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23594 VDD a_11872_14191# a_12047_14165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23595 a_40969_29967# a_17842_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23596 vcm a_18162_72234# a_38242_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23597 VSS a_5081_53135# a_6242_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23598 a_33299_32143# a_29163_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23599 VSS a_6975_76823# a_7092_74005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X236 VDD a_8723_67191# a_7899_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2360 VDD a_14839_66103# a_14839_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23600 a_44570_66210# pmat.rowon_n[10] a_44174_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23601 a_42258_70186# a_18546_70228# a_42166_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23602 a_29114_58138# pmat.row_n[2] a_29606_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23603 VDD a_11067_27239# a_30015_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23604 VDD pmat.rowoff_n[15] a_42166_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23605 a_23604_38567# a_22541_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23606 a_29510_11866# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23607 a_22792_28585# a_20616_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23608 a_33222_7484# a_18546_7482# a_33130_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23609 a_42166_64162# a_18162_64202# a_42258_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2361 a_45270_55126# a_18546_55168# a_45178_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23610 a_44453_53135# _1192_.B1 pmat.col_n[25] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23611 a_14521_69707# a_3615_71631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23612 a_47035_43817# a_46950_43719# a_46817_43541# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23613 VSS pmat.row_n[6] a_27502_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23614 a_13955_24847# a_11337_25071# a_13855_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23615 a_31518_60186# pmat.rowon_n[4] a_31122_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23616 a_31518_19898# nmat.rowon_n[4] a_31122_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23617 a_33141_51727# a_24591_28327# pmat.col_n[13] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23618 VDD a_5351_19913# a_13683_24847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23619 a_39154_21946# pmat.row_n[13] a_39646_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2362 a_22343_50613# a_22475_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X23620 a_39154_17930# a_18162_17524# a_39246_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23621 a_43170_70186# pmat.row_n[14] a_43662_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23622 VDD nmat.rowon_n[9] a_45178_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23623 VSS a_10873_36341# a_11292_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23624 a_9335_51727# a_9084_51843# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23625 a_43262_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23626 a_40158_12910# a_18162_12504# a_40250_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23627 a_5757_40097# a_4955_40277# a_5671_40097# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X23628 a_8084_71677# a_5779_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X23629 VDD a_19865_46983# a_19678_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2363 VDD ANTENNA__1190__A1.DIODE a_27531_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X23630 VDD VSS a_28110_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23631 a_6339_34863# a_5989_34863# a_6244_34863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23632 a_46182_63158# a_18162_63198# a_46274_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23633 a_4243_54991# a_3970_55311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23634 a_32218_58138# a_18546_58180# a_32126_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23635 a_8782_12559# a_8656_12675# a_8378_12691# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23636 VSS a_26283_42325# a_14497_42658# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23637 a_18235_34743# a_17113_34789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23638 VDD a_7658_71543# a_13183_72405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23639 a_6612_15797# a_3571_13627# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2364 a_6254_71017# a_6200_70919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X23640 a_11391_69831# a_11487_69653# a_11789_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23641 a_30610_9460# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23642 a_8105_7125# a_7939_7125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23643 a_37238_21540# a_18546_21538# a_37146_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23644 VDD nmat.rowon_n[10] a_49194_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23645 a_12069_38517# a_29023_38571# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X23646 a_7255_71829# a_6292_65479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23647 a_46674_10464# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23648 a_4345_34863# a_2563_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23649 a_15093_39638# a_13985_40229# a_15107_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X2365 a_45670_59504# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23650 a_19074_65166# a_18162_65206# a_19166_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23651 a_12521_28335# a_6830_22895# a_12437_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23652 a_6263_49373# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23653 a_23182_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23654 a_20078_60146# a_18162_60186# a_20170_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23655 VDD a_1923_53055# a_1643_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23656 a_29606_20504# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23657 VSS pmat.row_n[12] a_44570_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23658 a_29206_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23659 pmat.col_n[27] _1192_.A2 a_45557_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2366 VDD a_45019_38645# ANTENNA__1395__A2.DIODE VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.62e+12p ps=1.524e+07u w=1e+06u l=150000u M=4
X23660 a_8051_46607# a_8079_46519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23661 VDD a_1823_64213# a_3399_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23662 VDD a_17285_32117# nmat.rowoff_n[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23663 VSS a_19965_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23664 a_19566_12472# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23665 a_21082_23954# a_18162_23548# a_21174_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23666 VDD nmat.rowon_n[13] a_23090_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23667 a_2781_18377# a_1591_18005# a_2672_18377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23668 a_55610_40254# comp.adc_nor_latch_0.R VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23669 a_7467_63303# a_7131_64822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2367 VSS a_5232_72373# a_3956_72373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X23670 a_37146_63158# pmat.row_n[7] a_37638_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23671 a_34134_22950# a_18162_22544# a_34226_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23672 VDD a_2672_23817# a_2847_23743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23673 a_12020_39783# a_12235_39913# a_12162_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23674 a_21478_68218# pmat.rowon_n[12] a_21082_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23675 VSS pmat.row_n[3] a_47582_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23676 VDD pmat.rowon_n[8] a_44174_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23677 a_41654_61512# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23678 a_31214_19532# a_18546_19530# a_31122_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23679 a_51598_57174# pmat.rowon_n[1] a_51202_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2368 a_27560_36391# a_27605_37127# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X23680 a_26773_40955# a_26317_40726# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X23681 a_23083_47753# a_22733_47381# a_22988_47741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23682 a_26498_61190# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23683 a_39473_41605# a_39781_41245# a_31793_41570# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X23684 a_6339_34863# a_5823_34863# a_6244_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23685 VSS pmat.row_n[10] a_30514_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23686 VDD pmat.rowon_n[0] a_34134_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23687 a_4030_33231# a_2953_33237# a_3868_33609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23688 VDD a_1643_65301# a_1591_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23689 a_48586_55166# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2369 a_78165_40202# a_78261_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23690 a_45670_60508# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23691 VDD a_5779_71285# a_6749_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23692 a_39246_68178# a_18546_68220# a_39154_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23693 vcm a_18162_57174# a_31214_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23694 a_29079_47375# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23695 VSS a_5351_19913# a_9421_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23696 VSS a_3305_15823# a_13643_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23697 VDD a_8305_20871# a_11985_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23698 a_31518_14878# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23699 a_11530_77661# a_10772_77563# a_10967_77532# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X237 VSS a_14163_55295# a_14097_55369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X2370 VSS a_10515_13967# a_20776_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X23700 VDD a_2389_45859# a_5173_45993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23701 vcm a_18162_20536# a_36234_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23702 VDD a_7088_42479# a_7263_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23703 a_40158_57134# a_18162_57174# a_40250_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23704 a_12252_21583# a_12155_20719# a_11949_21237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23705 a_6853_55509# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23706 a_23090_67174# a_18162_67214# a_23182_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23707 a_28506_58178# pmat.rowon_n[2] a_28110_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23708 VDD pmat.rowon_n[4] a_22086_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23709 a_2289_29397# a_2422_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2371 a_33765_36965# a_33007_37683# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X23710 VSS a_6643_5724# a_6574_5853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23711 a_37238_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23712 VDD VDD a_37146_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23713 VSS _1187_.A2 pmat.col_n[22] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23714 a_2193_12342# a_1717_13647# a_1979_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23715 VDD a_7631_75895# a_6051_74183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X23716 VDD a_1591_74031# a_1899_76001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23717 a_12167_21263# a_12247_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23718 a_4174_26486# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23719 a_43566_7850# VDD a_43170_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2372 nmat.col[24] ANTENNA__1190__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=0p ps=0u w=650000u l=150000u M=4
X23720 a_21087_36649# a_19965_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23721 VSS a_18547_51565# a_19948_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23722 VSS pmat.row_n[11] a_20474_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23723 a_33567_30199# a_31339_31787# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23724 VSS pmat.row_n[0] a_50594_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23725 VDD a_6200_70919# a_6381_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23726 a_44174_15922# pmat.row_n[7] a_44666_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23727 a_19470_7850# VDD a_19074_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23728 VSS pmat.row_n[13] a_44570_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23729 a_47582_24918# VSS a_47186_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2373 vcm a_18162_8488# a_20170_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23730 VSS a_11444_55535# a_11711_56079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23731 a_31518_7850# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23732 a_6557_35105# a_6339_34863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23733 VSS a_12116_39783# a_24895_39605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23734 VSS pmat.row_n[10] a_33526_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23735 a_47678_57496# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23736 VDD VSS a_51202_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23737 VSS pmat.row_n[1] a_24490_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23738 VSS a_6179_69831# a_3936_70197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X23739 a_31614_23516# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2374 a_15210_51727# a_14452_51843# a_14647_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X23740 a_31214_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23741 VDD a_11337_25071# a_13798_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23742 a_30913_36603# a_29404_36165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X23743 a_37542_16886# nmat.rowon_n[7] a_37146_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23744 a_12049_66415# a_11797_60431# a_11977_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23745 a_10287_61127# a_10049_60663# a_10521_60975# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23746 a_2405_29967# a_2237_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23747 a_3141_38127# a_2935_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23748 a_5245_56053# a_5682_56311# a_5402_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23749 a_34226_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2375 VSS a_4461_26133# a_4395_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23750 VDD nmat.rowon_n[5] a_24094_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23751 a_19970_46287# a_19793_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23752 a_21574_15484# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23753 VSS pmat.row_n[4] a_47582_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23754 a_21478_21906# nmat.rowon_n[2] a_21082_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23755 a_51598_10862# nmat.rowon_n[13] a_51202_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23756 VDD cgen.enable_dlycontrol_in a_21815_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23757 a_38242_55126# a_18546_55168# a_38150_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23758 a_34626_14480# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23759 a_38642_59504# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2376 a_31518_12870# pmat.rowoff_n[4] a_31122_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23760 a_41335_52815# a_13091_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23761 a_32126_15922# a_18162_15516# a_32218_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23762 VSS a_5173_9839# a_5602_11791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23763 a_1643_56597# a_1846_56875# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23764 a_9369_58827# a_1769_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23765 a_4671_21629# a_4523_21276# a_4308_21495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23766 a_36538_63198# pmat.rowon_n[7] a_36142_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23767 a_22086_11906# pmat.row_n[3] a_22578_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23768 VDD a_24719_39605# a_14589_40726# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23769 vcm a_18162_9492# a_39246_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2377 a_43566_63198# pmat.rowon_n[7] a_43170_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23770 a_29206_24552# a_18546_24550# a_29114_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23771 a_28202_66170# a_18546_66212# a_28110_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23772 a_35138_10902# pmat.row_n[2] a_35630_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23773 a_50594_58178# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23774 VSS a_4976_16091# a_9749_19061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23775 VDD a_1923_69823# a_3476_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23776 VSS a_12003_52815# a_12353_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23777 a_6373_49249# a_6155_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23778 VDD pmat.rowon_n[12] a_32126_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23779 VDD _1224_.X a_24965_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2378 a_28110_55126# VDD a_28602_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23780 a_33526_68218# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23781 a_12292_44869# a_11133_44581# a_12196_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23782 VDD pmat.rowon_n[2] a_28110_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23783 a_6171_77661# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23784 a_49286_9492# a_18546_9490# a_49194_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23785 a_6853_55509# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23786 a_28506_11866# nmat.rowon_n[12] a_28110_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23787 a_35071_39913# a_33949_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23788 VDD a_2672_50095# a_2847_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23789 a_28245_44581# a_27789_44743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X2379 VDD a_3052_29967# a_3622_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23790 a_3484_58229# a_3938_58229# a_3876_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X23791 a_42322_47919# a_42292_47893# a_41663_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23792 a_20570_65528# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23793 a_46182_56130# pmat.row_n[0] a_46674_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23794 a_48190_70186# a_18162_70226# a_48282_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23795 vcm a_18162_62194# a_29206_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23796 VSS pmat.row_n[15] a_41558_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23797 a_29114_66170# pmat.row_n[10] a_29606_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23798 vcm a_18162_22544# a_51294_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23799 a_33222_60146# a_18546_60188# a_33130_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X238 VSS a_45019_38645# a_46863_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2380 a_19541_28879# a_19083_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X23800 a_33622_64524# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23801 a_32072_38567# a_30913_38779# a_31976_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23802 a_30118_61150# pmat.row_n[5] a_30610_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23803 vcm a_18162_12504# a_47278_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23804 a_4174_26159# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23805 VDD nmat.rowon_n[2] a_38150_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23806 a_51294_10496# a_18546_10494# a_51202_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23807 a_20170_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23808 a_24959_31055# a_25084_31287# a_25042_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23809 a_29772_40517# a_28613_40229# a_29676_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2381 VDD a_2847_41151# a_2834_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23810 a_17739_50871# a_18011_50729# a_17969_50755# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23811 a_30913_44219# a_29404_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X23812 a_38150_62154# a_18162_62194# a_38242_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23813 VSS pmat.row_n[12] a_20474_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23814 a_14301_27023# a_8861_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23815 a_42258_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23816 a_5809_51335# a_4399_51157# a_5972_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23817 a_23582_56492# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23818 a_1846_61651# a_2163_61761# a_2121_61885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23819 a_10838_30877# a_9761_30511# a_10676_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2382 a_40250_17524# a_18546_17522# a_40158_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X23820 a_2163_53057# a_1586_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23821 VSS a_28915_50959# a_46487_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23822 VSS pmat.row_n[14] a_45574_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23823 a_24186_12504# a_18546_12502# a_24094_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23824 a_34134_60146# pmat.row_n[4] a_34626_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23825 a_43262_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23826 a_40158_20942# a_18162_20536# a_40250_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23827 VSS a_7907_52031# a_7841_52105# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23828 vcm a_18162_68218# a_28202_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23829 a_39246_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2383 a_12069_10089# a_11501_10927# a_11987_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23830 VSS a_30489_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23831 VSS a_13909_39605# a_14328_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23832 a_6254_67753# a_5403_67655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23833 a_4308_21495# a_4523_21276# a_4450_21302# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23834 VSS pmat.row_n[6] a_35534_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23835 a_14491_51969# a_5363_33551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23836 VSS clk_dig a_7387_33231# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X23837 a_39013_42693# a_39321_42333# a_38737_41814# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X23838 VDD a_2325_17973# a_2215_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23839 VDD a_10781_42869# a_10725_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2384 a_2629_74031# a_2250_74397# a_2557_74031# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X23840 VSS pmat.row_n[5] a_48586_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23841 a_22482_70226# pmat.rowon_n[14] a_22086_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23842 a_45574_17890# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23843 a_50290_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23844 a_10071_17999# a_9820_18115# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X23845 a_36234_71190# a_18546_71232# a_36142_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23846 a_28202_11500# a_18546_11498# a_28110_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23847 vcm a_18162_8488# a_28202_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23848 a_39154_9898# a_18162_9492# a_39246_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23849 a_29206_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2385 vcm a_18162_21540# a_33222_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23850 a_40250_58138# a_18546_58180# a_40158_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23851 VDD pmat.rowon_n[7] a_36142_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23852 VSS a_9367_53511# a_7163_53333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X23853 a_22715_32521# a_22365_32149# a_22620_32509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23854 vcm a_18162_59182# a_49286_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23855 VSS a_2315_44124# a_4075_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23856 VSS nmat.sw a_5455_22057# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23857 a_6613_65577# a_5462_62215# a_6179_65479# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X23858 VDD a_25639_43957# a_12197_43746# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23859 a_25494_61190# pmat.rowon_n[5] a_25098_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2386 a_4985_74895# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X23860 a_49286_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23861 a_50198_58138# pmat.row_n[2] a_50690_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23862 a_28545_29423# a_16478_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23863 VSS pmat.row_n[9] a_22482_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23864 a_49590_16886# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23865 a_50594_11866# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23866 VDD a_33775_29111# a_33011_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X23867 a_6013_13103# a_5579_12394# a_5941_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23868 a_47186_10902# a_18162_10496# a_47278_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23869 a_37146_71190# pmat.row_n[15] a_37638_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2387 a_15048_35077# a_15144_35077# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X23870 a_34497_50959# a_30663_50087# a_34425_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23871 VDD a_5156_14025# a_5331_13951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23872 a_7648_9117# a_6872_8725# a_7040_8725# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23873 VDD VDD a_44174_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23874 a_33526_21906# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23875 a_30210_69182# a_18546_69224# a_30118_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23876 a_17224_47491# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23877 a_4298_69367# a_4583_68021# a_4529_68367# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23878 a_26194_59142# a_18546_59184# a_26102_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23879 vcm a_18162_56170# a_23182_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2388 VDD pmat.rowon_n[3] a_22086_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X23880 VDD a_6853_55509# a_6883_55862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23881 a_19622_49257# a_18547_51565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23882 a_29510_60186# pmat.rowon_n[4] a_29114_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23883 VSS pmat.row_n[8] a_26498_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23884 a_29510_19898# nmat.rowon_n[4] a_29114_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23885 a_23486_13874# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23886 a_28626_29423# a_27794_28879# a_28872_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.85e+11p pd=2.77e+06u as=0p ps=0u w=1e+06u l=150000u
X23887 a_14365_22351# a_13798_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23888 VDD a_4257_34319# a_4349_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23889 a_30514_14878# nmat.rowon_n[9] a_30118_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2389 a_41254_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23890 a_4075_68583# a_2389_45859# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23891 a_24186_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23892 VSS a_23455_32447# a_23389_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23893 a_43179_31599# a_42240_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23894 a_48586_63198# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23895 VSS pmat.row_n[13] a_38546_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23896 vcm a_18162_65206# a_31214_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23897 VDD a_32687_46607# a_33239_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23898 a_31122_69182# pmat.row_n[13] a_31614_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23899 a_42562_67214# pmat.rowon_n[11] a_42166_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X239 a_15839_49525# a_13091_52047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2390 a_13331_74953# a_12815_74581# a_13236_74941# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X23900 vcm a_18162_55166# a_27198_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23901 VDD a_4523_21276# a_13717_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23902 a_3175_59585# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23903 a_27106_59142# pmat.row_n[3] a_27598_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23904 a_1979_9334# a_2021_9563# a_1979_9661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23905 VDD a_5682_56311# a_6400_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23906 VSS a_4036_70741# a_3710_70455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X23907 VSS a_18975_40871# a_19925_41046# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23908 VDD a_32371_47349# a_31105_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23909 a_40158_65166# a_18162_65206# a_40250_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2391 a_37638_24520# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23910 a_39246_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23911 a_7393_68047# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X23912 a_10959_23983# a_10515_24233# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X23913 a_30645_29673# a_30603_29575# a_30561_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23914 a_29685_34954# clk_ena VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23915 VSS a_2263_43719# a_29233_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23916 a_2107_23817# a_1591_23445# a_2012_23805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23917 a_39550_65206# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23918 vcm a_18162_17524# a_22178_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23919 a_39646_17492# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2392 VSS a_19817_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23920 a_28202_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23921 a_47582_9858# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23922 a_15397_32509# a_11067_64015# a_15325_32509# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23923 a_6171_77661# a_5547_77295# a_6063_77295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23924 VDD pmat.rowoff_n[7] a_43170_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23925 a_37146_18934# a_18162_18528# a_37238_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23926 a_45005_32687# a_40837_46261# a_44923_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23927 VSS a_3883_65845# a_3814_65871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23928 a_5423_30485# a_5248_30511# a_5602_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23929 VDD a_2672_8585# a_2847_8511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2393 a_15383_44265# a_14261_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X23930 a_7013_40303# a_5823_40303# a_6904_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23931 VSS a_24719_38517# a_14773_39394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23932 a_26234_27497# a_16311_28327# a_25931_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23933 a_12047_14165# a_11872_14191# a_12226_14191# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23934 a_19470_68218# pmat.rowon_n[12] a_19074_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23935 a_8782_63695# a_8656_63811# a_8378_63827# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23936 vcm a_18162_16520# a_26194_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23937 a_49590_57174# pmat.rowon_n[1] a_49194_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23938 a_44174_66170# a_18162_66210# a_44266_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23939 a_30210_14512# a_18546_14510# a_30118_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2394 VDD nmat.rowon_n[1] a_41162_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X23940 a_30514_71230# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23941 a_12337_18005# a_12171_18005# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23942 VSS a_22357_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X23943 a_44666_11468# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23944 VSS pmat.row_n[8] a_29510_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23945 a_34724_44527# a_34547_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23946 a_10779_21583# a_10071_17999# a_10441_21263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23947 a_27598_21508# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23948 a_27198_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23949 VDD a_40951_31599# a_45287_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X2395 VDD pmat.rowon_n[7] pmat.rowoff_n[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X23950 VSS a_10751_72917# a_10699_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23951 a_22733_47381# a_22567_47381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23952 VSS a_5047_76983# a_4993_77071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23953 a_34226_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23954 VSS config_2_in[11] a_1591_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X23955 VSS a_6787_47607# a_6200_70919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23956 VSS pmat.row_n[0] a_19470_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23957 a_34530_9858# nmat.rowon_n[14] a_34134_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23958 a_51598_60186# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23959 a_21174_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2396 a_28506_10862# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23960 a_51598_19898# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23961 a_22357_43493# a_20848_41605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X23962 VSS a_1674_68047# a_2695_76757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23963 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23964 a_34530_70226# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23965 VDD nmat.rowon_n[12] a_21082_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23966 a_38242_63158# a_18546_63200# a_38150_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23967 VSS a_10864_68565# a_11433_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23968 a_38642_67536# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23969 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2397 pmat.rowon_n[12] a_14839_65871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23970 a_32126_23954# a_18162_23548# a_32218_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23971 VDD pmat.rowon_n[9] a_42166_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23972 a_28110_13914# a_18162_13508# a_28202_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23973 a_29051_37607# a_23821_35279# a_29225_37483# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23974 a_11867_64899# a_10921_64786# a_11795_64899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23975 VSS a_35382_34191# a_36203_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23976 a_30473_49871# a_10883_3303# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23977 a_48190_63158# pmat.row_n[7] a_48682_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23978 a_24490_62194# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23979 VSS a_14773_39394# a_13837_39069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X2398 a_9943_15645# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X23980 a_3415_9839# a_3142_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23981 a_11292_40719# a_11041_40948# a_11071_41046# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23982 a_31976_38567# a_30913_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23983 VSS pmat.row_n[14] a_38546_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23984 a_42562_20902# pmat.rowoff_n[12] a_42166_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23985 vcm a_18162_71230# a_25190_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23986 a_4241_7663# a_2972_9991# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23987 a_12270_32182# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23988 VDD pmat.rowon_n[0] a_45178_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23989 a_25590_24520# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2399 a_23823_47679# a_23648_47753# a_24002_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X23990 a_2107_16201# a_1757_15829# a_2012_16189# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23991 VDD pmat.rowon_n[10] a_28110_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23992 a_3797_14709# a_3579_15113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23993 a_40125_31029# a_39939_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23994 a_39469_43493# a_39013_43655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X23995 a_29308_44869# a_28245_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23996 a_10923_17782# a_10741_17782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23997 a_28202_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23998 VSS config_2_in[9] a_2603_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X23999 a_17900_41831# a_16837_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_34887_39095# a_34277_38550# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X240 a_12934_35823# a_12757_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2400 a_34530_65206# pmat.rowon_n[9] a_34134_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24000 vcm.sky130_fd_sc_hd__nand2_1_1.A vcm.sky130_fd_sc_hd__buf_4_0.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24001 a_9485_15279# a_9319_15279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24002 VDD a_1781_9308# a_2193_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24003 a_7995_54281# a_7645_53909# a_7900_54269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24004 vcm a_18162_70226# a_29206_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24005 VDD nmat.rowon_n[15] a_41162_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24006 a_4032_26311# a_4068_25615# a_4174_26486# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24007 VDD VSS a_49194_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24008 VDD a_1586_18231# a_1591_18005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24009 a_7367_31055# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2401 VSS a_45450_48695# a_44697_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.3585e+12p ps=1.328e+07u w=650000u l=150000u M=4
X24010 a_8309_49007# a_8267_49159# a_7578_48553# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24011 a_26102_20942# pmat.row_n[12] a_26594_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24012 a_33622_72556# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24013 a_41558_68218# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24014 a_26102_16926# a_18162_16520# a_26194_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24015 vcm a_18162_20536# a_47278_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24016 VSS a_3199_40455# a_3149_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24017 a_29606_62516# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24018 a_30210_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24019 a_27155_31599# a_20616_27791# a_26983_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X2402 a_2586_29967# a_2051_29973# a_2500_30345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X24020 VDD pmat.rowon_n[4] a_33130_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24021 a_5621_47081# a_4985_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24022 VSS a_2163_69821# a_2124_69947# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24023 a_35646_29967# a_35520_30083# a_35242_30099# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X24024 a_5935_46983# a_6637_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24025 a_14369_50095# a_11711_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24026 a_19470_21906# nmat.rowon_n[2] a_19074_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24027 a_49590_10862# nmat.rowon_n[13] a_49194_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24028 nmat.col_n[11] a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24029 a_20570_10464# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2403 VSS a_10287_61127# a_10195_59861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24030 a_23486_8854# nmat.rowon_n[15] a_23090_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24031 a_12075_24233# a_10959_23983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X24032 a_34895_31849# a_34243_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24033 a_7509_63401# a_7467_63303# a_7321_63151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24034 a_44570_59182# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24035 a_24186_20536# a_18546_20534# a_24094_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24036 a_38546_24918# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24037 a_28507_52245# a_18243_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24038 a_42166_16926# pmat.row_n[8] a_42658_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24039 a_27502_69222# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2404 vcm a_18162_13508# a_41254_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24040 VSS pmat.row_n[11] a_31518_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24041 a_14466_29199# a_13479_26935# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24042 VSS a_28704_29568# a_40969_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24043 VDD a_5687_71829# a_6749_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24044 a_28110_58138# a_18162_58178# a_28202_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24045 VSS pmat.row_n[3] a_21478_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24046 a_18660_47607# a_12263_50959# a_18891_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24047 VDD a_5087_19319# a_5087_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X24048 a_48586_16886# nmat.rowon_n[7] a_48190_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24049 vcm a_18162_68218# a_36234_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2405 a_3305_15823# a_2847_16127# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X24050 a_4525_44905# a_2983_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24051 a_28110_17930# pmat.row_n[9] a_28602_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24052 VDD pmat.rowon_n[15] a_36142_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24053 a_14365_68743# a_3615_71631# a_14528_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24054 a_32618_15484# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24055 vcm a_18162_67214# a_49286_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24056 a_36234_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24057 a_38242_8488# a_18546_8486# a_38150_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24058 vcm a_18162_62194# a_50290_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24059 a_29272_28111# ANTENNA__1190__A1.DIODE a_28969_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2406 a_32771_31599# a_9963_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X24060 a_50198_66170# pmat.row_n[10] a_50690_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24061 a_49286_55126# a_18546_55168# a_49194_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24062 a_19166_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24063 VSS a_6795_76989# a_9225_76207# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24064 a_49686_59504# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24065 VSS pmat.row_n[2] a_25494_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24066 a_22482_55166# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24067 VDD a_1923_61759# a_1643_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24068 a_27986_50095# a_22199_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24069 cgen.dlycontrol2_in[1] a_1591_38127# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2407 a_47582_64202# pmat.rowon_n[8] a_47186_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24070 a_26194_67174# a_18546_67216# a_26102_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24071 VDD a_20776_51959# a_19579_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X24072 a_1757_15829# a_1591_15829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24073 vcm a_18162_64202# a_23182_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24074 a_33130_11906# pmat.row_n[3] a_33622_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24075 a_19074_19938# pmat.row_n[11] a_19566_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24076 VSS a_2163_61761# a_2124_61635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24077 a_21621_40955# a_19409_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X24078 a_23090_68178# pmat.row_n[12] a_23582_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24079 a_6168_32687# a_5087_32687# a_5821_32929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2408 VDD pmat.sample a_18546_68220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X24080 VDD a_14504_37607# a_12513_36924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24081 VDD pmat.rowon_n[13] a_30118_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24082 a_44266_17524# a_18546_17522# a_44174_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24083 VSS a_1781_9308# a_2200_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24084 VDD pmat.rowon_n[3] a_26102_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24085 a_14471_27247# a_12987_26159# a_14471_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24086 a_38913_31055# a_25575_31055# a_38759_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24087 VSS a_2715_51969# a_2676_51843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24088 a_30210_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24089 VDD a_1674_57711# a_7847_56085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2409 a_38150_20942# pmat.row_n[12] a_38642_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24090 a_41558_21906# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24091 VDD a_16478_29423# a_28456_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24092 a_14648_64015# a_10055_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24093 a_44174_57134# pmat.row_n[1] a_44666_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24094 VDD config_2_in[2] a_1591_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X24095 a_2882_52815# a_2124_52931# a_2319_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24096 vcm a_18162_63198# a_27198_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24097 a_27106_67174# pmat.row_n[11] a_27598_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24098 a_38546_65206# pmat.rowon_n[9] a_38150_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24099 a_7165_13353# a_5173_9839# a_7093_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X241 a_4263_49007# a_2389_45859# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.5875e+11p pd=9.45e+06u as=0p ps=0u w=650000u l=150000u M=4
X2410 VDD a_7840_27247# a_18200_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.345e+12p ps=1.269e+07u w=1e+06u l=150000u M=4
X24100 a_31614_65528# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24101 a_48282_16520# a_18546_16518# a_48190_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24102 vcm a_18162_13508# a_45270_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24103 VSS a_40352_41831# a_39781_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X24104 a_31122_55126# a_18162_55166# a_31214_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24105 a_44570_12870# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24106 VSS a_10391_69653# a_10325_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24107 a_21574_57496# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24108 a_47861_27497# a_17139_30503# nmat.col_n[27] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X24109 a_27502_22910# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2411 VDD a_38851_28327# a_47731_36103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X24110 a_14558_3311# _1184_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24111 a_31122_14918# pmat.row_n[6] a_31614_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24112 VSS pmat.row_n[12] a_31518_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24113 a_11277_77295# a_10898_77661# a_11205_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24114 a_16837_40955# a_16171_40157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X24115 a_34626_56492# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24116 a_22178_13508# a_18546_13506# a_22086_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24117 a_14641_57711# a_14287_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24118 a_11138_50347# a_11455_50237# a_11413_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24119 a_23700_38567# a_22541_38779# a_23663_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X2412 a_38150_16926# a_18162_16520# a_38242_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24120 a_22537_36911# a_22111_36950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24121 a_27198_7484# a_18546_7482# a_27106_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24122 VSS a_10943_8903# a_10378_7637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24123 a_24765_28111# a_13459_28111# nmat.col_n[4] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24124 VDD a_7373_48695# a_5411_48695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X24125 a_13537_54447# a_11202_55687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24126 a_24490_15882# pmat.rowoff_n[7] a_24094_15922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24127 VSS pmat.row_n[4] a_21478_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24128 a_24955_30761# a_23933_32143# a_24737_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24129 a_12792_12937# a_11877_12565# a_12445_12533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2413 a_4144_15113# a_3063_14741# a_3797_14709# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X24130 a_5779_30006# a_4719_30287# a_5320_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24131 a_45325_38127# a_45047_38155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X24132 vcm a_18162_24552# a_26194_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24133 VSS pmat.row_n[6] a_46578_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24134 a_43566_18894# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24135 a_50594_60186# pmat.rowon_n[4] a_50198_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24136 a_10055_22671# a_6664_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24137 a_50594_19898# nmat.rowon_n[4] a_50198_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24138 VSS VDD a_29510_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24139 a_15657_52317# a_11435_58791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2414 VDD nmat.rowon_n[2] a_45178_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X24140 pmat.col[17] a_34705_51959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24141 a_12231_16367# a_11785_16367# a_12135_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24142 a_33526_70226# pmat.rowon_n[14] a_33130_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24143 a_25590_58500# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24144 a_47278_71190# a_18546_71232# a_47186_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24145 VSS pmat.row_n[3] a_25494_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24146 a_8915_6409# a_8565_6037# a_8820_6397# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X24147 a_14264_72777# a_13349_72405# a_13917_72373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24148 VDD VSS a_47186_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24149 VSS a_40951_31599# a_44933_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2415 a_2659_35015# a_5558_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X24150 a_51294_58138# a_18546_58180# a_51202_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24151 a_23486_62194# pmat.rowon_n[6] a_23090_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24152 a_17136_28995# a_16863_29239# a_17054_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24153 a_24586_9460# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24154 VSS a_10055_31591# a_14809_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24155 a_5205_37039# a_4257_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24156 a_35630_21508# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24157 a_35230_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24158 a_17690_47081# a_14653_53458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24159 a_48190_71190# pmat.row_n[15] a_48682_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2416 a_42258_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24160 a_48682_20504# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24161 a_19611_27247# a_7415_29397# a_19439_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X24162 a_48282_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24163 a_22086_70186# a_18162_70226# a_22178_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24164 a_44449_31029# a_43776_30287# a_44695_31393# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24165 a_17007_50613# a_17163_50857# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X24166 a_5738_10927# a_4865_12533# a_5012_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X24167 a_6800_44629# a_4257_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24168 VDD a_9075_28023# a_11409_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24169 vcm a_18162_12504# a_21174_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2417 a_48282_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24170 a_14533_39631# a_14107_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24171 a_38642_12472# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24172 VDD a_35540_46983# a_35068_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24173 a_36142_13914# a_18162_13508# a_36234_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24174 VDD nmat.rowon_n[13] a_42166_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24175 a_10943_8903# a_9583_10121# a_11117_8779# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24176 a_36538_8854# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24177 a_20855_36885# a_21031_37217# a_20983_37277# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24178 a_41964_29423# a_41237_28585# a_41703_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24179 VSS a_46817_27221# nmat.col[27] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2418 VSS a_46753_41935# a_41731_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.053e+12p ps=1.104e+07u w=650000u l=150000u M=12
X24180 VDD pmat.rowoff_n[12] a_25098_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24181 a_40554_68218# pmat.rowon_n[12] a_40158_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24182 a_6521_67753# a_6451_67655# a_6087_67655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24183 a_49194_12910# a_18162_12504# a_49286_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24184 a_50290_19532# a_18546_19530# a_50198_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24185 a_28202_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24186 a_25098_61150# a_18162_61190# a_25190_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24187 VSS pmat.row_n[13] a_49590_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24188 VSS pmat.row_n[0] a_46578_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24189 a_22357_43493# a_20848_41605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X2419 a_45178_62154# a_18162_62194# a_45270_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24190 a_2129_12559# a_1959_12559# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24191 a_20217_32509# a_20173_32117# a_20051_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X24192 a_2250_56989# a_2124_56891# a_1846_56875# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X24193 a_26102_24958# a_18162_24552# a_26194_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24194 a_29606_70548# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24195 vcm a_18162_18528# a_20170_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24196 a_30210_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24197 VDD a_1923_61759# a_2655_59317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24198 a_43566_59182# pmat.rowon_n[3] a_43170_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24199 a_37638_18496# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X242 a_15101_29423# a_14829_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2420 a_1828_25589# a_2007_25597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24200 a_26194_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24201 VDD nmat.rowon_n[7] a_41162_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24202 a_26498_69222# pmat.rowon_n[13] a_26102_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24203 a_29114_60146# a_18162_60186# a_29206_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24204 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24205 VDD a_27405_52245# pmat.col_n[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24206 a_25647_39783# a_21981_34191# a_25821_39659# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24207 vcm a_18162_17524# a_33222_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24208 VDD a_45187_38129# a_45047_38155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24209 a_48190_18934# a_18162_18528# a_48282_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2421 a_37542_56170# pmat.rowon_n[0] a_37146_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24210 VDD nmat.rowon_n[12] a_19074_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24211 VSS a_1923_31743# a_7521_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24212 VSS clk_vcm vcm.sky130_fd_sc_hd__inv_1_4.Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24213 a_12792_12937# a_11711_12565# a_12445_12533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24214 a_44976_47349# a_33423_47695# a_45196_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24215 VSS _1224_.X a_46027_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24216 a_42166_67174# a_18162_67214# a_42258_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24217 a_47582_58178# pmat.rowon_n[2] a_47186_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24218 VSS VDD a_44570_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24219 VSS a_12447_16143# a_16833_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2422 a_28110_72194# a_18162_72234# a_28202_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24220 VSS a_20616_27791# a_27167_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24221 a_48190_8894# a_18162_8488# a_48282_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24222 VDD a_15163_32375# a_14839_20871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24223 a_43170_7890# VDD a_43662_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24224 VSS pmat.row_n[9] a_27502_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24225 a_45368_47375# a_43315_48437# a_45113_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24226 a_21082_10902# a_18162_10496# a_21174_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24227 VSS a_12449_22895# a_14696_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24228 a_5550_34319# a_4792_34435# a_4987_34293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24229 a_19074_7890# VDD a_19566_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2423 a_30610_56492# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24230 a_13814_59663# a_10239_14183# a_13728_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24231 a_11941_47919# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24232 _1519_.A a_46804_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X24233 a_30485_31849# a_30412_31751# a_29635_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24234 VSS cgen.enable_dlycontrol_in a_23655_35279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24235 VDD a_8305_20871# a_8263_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24236 a_16478_29423# a_16131_29429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X24237 a_21478_55166# VSS a_21082_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24238 a_29606_7452# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24239 a_25494_7850# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2424 a_4913_40303# a_4705_39759# a_4831_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24240 VDD pmat.rowon_n[5] a_27106_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24241 VSS a_1739_47893# a_1775_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24242 a_32218_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24243 a_9368_9991# comp_latch a_9510_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24244 a_45405_30511# a_30663_50087# a_45321_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24245 VDD a_23648_47753# a_23823_47679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24246 a_25681_28879# a_25327_28992# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24247 vcm a_18162_70226# a_50290_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24248 a_49286_63158# a_18546_63200# a_49194_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24249 a_36789_52245# a_34705_51959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2425 VDD nmat.rowon_n[10] a_35138_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X24250 a_36142_58138# a_18162_58178# a_36234_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24251 a_50690_23516# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24252 VSS a_29797_51701# pmat.col_n[10] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24253 a_49686_67536# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24254 a_50290_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24255 a_12128_32375# a_7939_31591# a_12270_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24256 a_22482_63198# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24257 a_11829_53359# a_9463_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24258 a_19074_68178# a_18162_68218# a_19166_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24259 a_16607_36911# a_16430_36911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2426 a_32218_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24260 a_26317_40726# a_25393_41317# a_26456_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X24261 a_49194_57134# a_18162_57174# a_49286_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24262 a_36142_17930# pmat.row_n[9] a_36634_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24263 a_35534_62194# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24264 VSS pmat.row_n[15] a_36538_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24265 a_40650_15484# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24266 a_40554_21906# nmat.rowon_n[2] a_40158_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24267 vcm a_18162_72234# a_23182_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24268 VDD pmat.rowon_n[1] a_43170_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24269 VSS pmat.row_n[14] a_49590_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2427 a_10147_29415# a_36453_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X24270 a_20078_22950# pmat.row_n[14] a_20570_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24271 a_5173_9839# a_2972_9991# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24272 nmat.rowon_n[1] a_14195_7119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24273 VDD a_5423_30485# a_5410_30877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24274 VDD pmat.rowon_n[11] a_26102_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24275 a_51202_15922# a_18162_15516# a_51294_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24276 a_11258_18870# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24277 a_8201_67503# a_5363_70543# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24278 a_33222_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24279 a_26194_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2428 VDD a_34924_36165# a_34828_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X24280 a_43566_12870# pmat.rowoff_n[4] a_43170_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24281 a_8539_76181# a_9183_76359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24282 a_41162_11906# pmat.row_n[3] a_41654_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24283 a_27340_31055# a_15101_29423# a_27249_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24284 a_26498_64202# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24285 VDD a_33436_34191# a_33542_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24286 a_26498_22910# nmat.rowon_n[1] a_26102_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24287 a_24094_21946# pmat.row_n[13] a_24586_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24288 a_24094_17930# a_18162_17524# a_24186_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24289 vcm a_18162_21540# a_45270_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2429 VDD a_10967_77532# a_10898_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X24290 a_48282_24552# a_18546_24550# a_48190_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24291 VDD nmat.rowon_n[9] a_30118_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24292 VDD pmat.rowon_n[3] a_34134_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24293 a_27535_27497# a_10883_3303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24294 VSS a_4608_41909# a_4542_42313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X24295 a_82783_53524# _1519_.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24296 VDD a_13697_47349# a_12604_47080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24297 a_31122_63158# a_18162_63198# a_31214_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24298 nmat.rowon_n[9] a_13446_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24299 a_11071_41046# a_11041_40948# a_10999_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 VDD pmat.rowon_n[14] a_44174_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2430 VDD a_2727_58470# a_4259_65103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X24300 VDD pmat.rowon_n[2] a_47186_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24301 VSS a_37291_29397# a_47685_30517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24302 a_2847_43327# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24303 a_17499_38825# a_16377_38779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24304 a_47582_11866# nmat.rowon_n[12] a_47186_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24305 VDD a_11852_49783# a_11803_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24306 a_27106_12910# pmat.row_n[4] a_27598_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24307 VSS a_2007_76970# a_1823_77821# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X24308 VSS a_45251_53047# pmat.col[25] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24309 a_22178_21540# a_18546_21538# a_22086_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2431 a_31214_12504# a_18546_12502# a_31122_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X24310 a_8179_71689# a_7663_71317# a_8084_71677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24311 a_28267_50639# a_28131_50069# a_28049_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24312 a_31614_10464# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24313 a_10233_19881# a_10045_19677# a_10151_19637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24314 a_2944_65576# a_3609_65015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24315 VSS a_9963_13967# a_14458_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24316 VSS a_8767_16055# a_8767_15823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X24317 vcm a_18162_69222# a_43262_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24318 a_9393_17455# a_4976_16091# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24319 a_15420_41831# a_14261_42043# a_15324_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2432 a_4351_55527# a_4927_50613# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X24320 a_35077_50095# a_30571_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24321 a_36465_28879# a_31263_28309# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24322 VDD a_4461_46805# a_4491_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24323 a_2122_17455# a_1945_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24324 a_47186_9898# pmat.row_n[1] a_47678_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24325 a_40158_19938# pmat.row_n[11] a_40650_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24326 a_4333_7913# a_2972_9991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24327 VDD a_14773_39394# a_13837_39069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X24328 VDD a_3339_70759# a_6619_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24329 a_4675_54599# a_4025_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2433 VSS a_23741_42567# a_23939_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X24330 a_44266_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24331 a_6639_63927# a_6568_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24332 a_25190_62154# a_18546_62196# a_25098_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24333 a_6987_15279# a_6541_15279# a_6891_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24334 a_25590_66532# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24335 a_22086_63158# pmat.row_n[7] a_22578_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24336 a_17033_51183# a_16679_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24337 a_42258_9492# a_18546_9490# a_42166_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24338 a_4266_18365# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24339 VSS pmat.row_n[3] a_32522_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2434 VDD pmat.rowoff_n[4] a_48190_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X24340 a_43262_12504# a_18546_12502# a_43170_12910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24341 VSS a_2935_38279# a_3983_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24342 vcm a_18162_68218# a_47278_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24343 VDD a_1923_31743# a_1643_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24344 a_47278_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24345 a_46857_45199# a_43720_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24346 a_26102_62154# pmat.row_n[6] a_26594_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24347 a_42240_29423# a_41703_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X24348 a_30610_60508# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24349 a_33526_55166# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2435 vcm a_18162_19532# a_40250_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24350 a_19176_35279# a_18999_35279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24351 VDD nmat.rowon_n[14] a_34134_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24352 a_11258_18543# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24353 a_24186_68178# a_18546_68220# a_24094_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24354 a_48282_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24355 a_45178_21946# a_18162_21540# a_45270_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24356 a_5179_59663# a_3866_57399# a_5085_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24357 VSS a_25839_49783# a_25785_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24358 a_42258_18528# a_18546_18526# a_42166_18934# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24359 VSS a_18563_27791# a_37837_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2436 a_50290_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24360 VDD a_10839_11989# a_10471_12791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24361 vcm a_18162_20536# a_21174_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24362 VSS a_11892_21959# a_11897_21813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24363 a_44570_61190# pmat.rowon_n[5] a_44174_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24364 VSS a_43781_52245# pmat.col_n[24] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24365 VSS pmat.row_n[9] a_41558_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24366 VDD nmat.sw a_12191_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24367 VSS a_14947_26159# a_15749_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24368 VSS a_10515_61839# a_14287_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24369 a_12271_24233# a_7026_24527# a_12147_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X2437 VDD a_25997_42902# a_26272_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X24370 a_27502_71230# pmat.rowon_n[15] a_27106_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24371 VDD ANTENNA__1395__A1.DIODE a_37007_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24372 a_19595_47491# a_16800_47213# a_19523_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24373 a_22178_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24374 a_9135_49257# a_4719_30287# a_9217_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24375 a_8765_76725# a_8547_77129# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24376 VSS a_36617_37691# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X24377 a_17811_39605# a_13909_39605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24378 a_49194_20942# a_18162_20536# a_49286_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24379 a_7405_32441# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2438 VDD pmat.sample_n a_18162_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X24380 vcm a_18162_14512# a_43262_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24381 a_40969_30287# a_25575_31055# a_41053_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24382 a_45270_59142# a_18546_59184# a_45178_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24383 vcm a_18162_56170# a_42258_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24384 a_26475_34343# a_24833_34191# a_26649_34219# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24385 a_2163_67645# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24386 a_12705_10389# a_12539_10389# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24387 a_2012_41213# a_1895_41018# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24388 a_26767_46831# a_26321_46831# a_26671_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24389 a_12032_59887# a_5651_66975# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2439 a_46274_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24390 a_16671_39913# a_15549_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24391 VSS pmat.row_n[8] a_45574_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24392 a_42562_13874# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24393 a_43262_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24394 VSS a_33395_43455# a_33341_43777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24395 a_25494_23914# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24396 a_9090_73487# a_8013_73493# a_8928_73865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24397 VDD a_4312_74005# a_4048_74549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X24398 a_32522_24918# VSS a_32126_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24399 a_2157_14013# a_2122_13779# a_1687_13621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X244 vcm a_18162_69222# a_26194_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2440 vcm a_18162_68218# a_35230_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24400 a_19166_19532# a_18546_19530# a_19074_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24401 a_26194_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24402 a_11979_47068# a_11784_47099# a_12289_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24403 a_39472_47753# a_38557_47381# a_39125_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24404 a_37238_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24405 a_32618_57496# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24406 VDD a_43971_28487# a_27763_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X24407 a_42258_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24408 vcm a_18162_55166# a_46274_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24409 a_9834_6397# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2441 a_22178_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24410 a_5823_52521# a_5784_52423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24411 a_46182_59142# pmat.row_n[3] a_46674_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24412 a_22482_16886# nmat.rowon_n[7] a_22086_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24413 a_12557_30485# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24414 a_13439_8207# a_12815_8213# a_13331_8585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24415 a_14749_48285# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24416 VSS a_4383_7093# a_6559_6031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24417 VSS a_25695_28111# a_35717_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24418 a_28715_28879# a_28442_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24419 VSS a_36561_38780# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X2442 VDD a_2163_53057# a_2124_52931# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24420 VSS pmat.row_n[4] a_32522_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24421 VSS pmat.row_n[7] a_44570_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24422 a_7937_61519# a_5784_52423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24423 a_10593_15823# a_10423_15823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X24424 a_34530_69222# pmat.rowon_n[13] a_34134_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24425 vcm a_18162_57174# a_19166_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24426 vcm a_18162_17524# a_41254_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24427 a_23182_55126# a_18546_55168# a_23090_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24428 VSS a_82787_26133# nmat.col_n[26] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24429 a_23582_59504# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2443 VSS a_33719_44527# a_33825_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24430 VDD a_23280_32521# a_23455_32447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24431 a_19470_14878# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24432 a_1881_67503# a_1846_67755# a_1643_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24433 a_2244_26935# rst_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24434 a_38150_24958# VDD a_38642_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24435 a_42658_22512# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24436 a_37612_30663# a_37820_30485# a_37754_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24437 a_2369_41213# a_2325_40821# a_2203_41225# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24438 a_21478_63198# pmat.rowon_n[7] a_21082_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24439 a_1925_26935# a_2021_26677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2444 a_8491_47911# a_6787_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X24440 VSS pmat.row_n[9] a_35534_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24441 a_3517_11849# a_2327_11477# a_3408_11849# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24442 a_10751_72917# a_10954_73195# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24443 VDD nmat.rowon_n[6] a_35138_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24444 a_8581_73461# a_8363_73865# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X24445 VSS pmat.row_n[8] a_48586_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24446 a_9023_6031# a_8399_6037# a_8915_6409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24447 a_10979_42390# a_11021_42619# a_10979_42717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24448 VDD VDD a_39154_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24449 VSS VDD a_35534_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2445 VDD a_5417_11445# a_5223_11079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24450 a_46674_21508# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24451 a_43170_14918# a_18162_14512# a_43262_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24452 a_51202_7890# VDD a_51694_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24453 a_46274_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24454 VSS a_30765_37692# a_30457_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24455 a_38293_51727# _1184_.A2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24456 a_49194_65166# a_18162_65206# a_49286_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24457 VDD a_21981_34191# a_25647_37607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24458 a_40554_9858# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24459 a_50198_60146# a_18162_60186# a_50290_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2446 a_10885_64899# a_10423_64786# a_10789_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=2.43e+11p ps=2.66e+06u w=420000u l=150000u
X24460 VSS pmat.row_n[0] a_38546_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24461 a_45574_7850# VDD a_45178_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24462 a_31122_56130# pmat.row_n[0] a_31614_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24463 a_40250_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24464 a_33130_70186# a_18162_70226# a_33222_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24465 VDD nmat.rowon_n[7] a_39154_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24466 a_36634_13476# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24467 VDD nmat.rowon_n[12] a_40158_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24468 a_25494_64202# pmat.rowon_n[8] a_25098_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24469 a_19566_23516# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2447 VSS VDD a_25494_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X24470 vcm a_18162_12504# a_32218_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24471 a_19166_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24472 a_8378_12691# a_8695_12801# a_8653_12925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24473 a_51202_23954# a_18162_23548# a_51294_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24474 VSS a_2944_72104# a_2882_72221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24475 a_49686_12472# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24476 VDD nmat.rowon_n[2] a_23090_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24477 a_14426_72399# a_13349_72405# a_14264_72777# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24478 VSS a_2935_38279# a_4154_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24479 a_47186_13914# a_18162_13508# a_47278_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2448 a_10515_13967# a_21063_48723# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X24480 a_26194_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24481 a_23090_62154# a_18162_62194# a_23182_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24482 a_9258_50345# a_7373_49007# a_9176_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24483 VSS pmat.row_n[1] a_26498_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24484 a_44763_34293# a_44647_35520# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24485 a_51598_68218# pmat.rowon_n[12] a_51202_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24486 a_9579_26159# a_9135_26409# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X24487 a_26498_72234# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24488 a_45837_27791# a_16311_28327# nmat.col_n[25] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X24489 a_41876_52047# ANTENNA__1197__A.DIODE a_41573_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2449 a_44570_7850# VDD a_44174_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24490 VSS pmat.row_n[14] a_30514_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24491 VSS a_4124_28023# a_2283_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24492 a_37146_7890# a_18162_7484# a_37238_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24493 vcm a_18162_71230# a_44266_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24494 VDD pmat.rowon_n[11] a_34134_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24495 a_5857_74031# a_6051_74183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24496 VDD pmat.rowoff_n[4] a_26102_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24497 a_24186_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24498 a_39472_47753# a_38391_47381# a_39125_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24499 a_12981_74581# a_12815_74581# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X245 VSS a_10781_42364# a_11200_42717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2450 a_19423_37737# a_19817_37692# a_13597_37571# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X24500 VDD pmat.rowon_n[10] a_47186_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24501 a_44666_63520# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24502 VSS pmat.row_n[6] a_20474_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24503 a_9913_69679# a_9869_69921# a_9747_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24504 a_47278_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24505 a_36419_28023# a_26891_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24506 a_19470_55166# VSS a_19074_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24507 a_30015_51727# a_21739_29415# a_29797_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24508 VDD a_12020_39783# a_11565_39061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24509 a_2672_18377# a_1757_18005# a_2325_17973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2451 a_39757_50700# a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24510 a_34530_22910# nmat.rowon_n[1] a_34134_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24511 VSS pmat.row_n[5] a_33526_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24512 a_30514_17890# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24513 a_21174_71190# a_18546_71232# a_21082_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24514 VDD a_12449_40693# a_12479_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24515 a_38546_58178# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24516 a_40158_68178# a_18162_68218# a_40250_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24517 a_18597_31599# a_18243_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24518 VSS _1183_.A2 a_83092_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24519 VDD pmat.rowon_n[7] a_21082_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2452 a_20078_22950# a_18162_22544# a_20170_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24520 a_23090_8894# pmat.row_n[0] a_23582_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24521 a_48682_62516# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24522 a_16657_42567# a_16745_44581# a_17867_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24523 a_6087_70919# a_2879_57487# a_6432_70767# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X24524 vcm a_18162_59182# a_34226_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24525 VSS a_31412_43439# a_31518_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24526 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24527 a_46765_52815# ANTENNA__1197__A.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24528 a_34530_16886# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24529 a_25190_70186# a_18546_70228# a_25098_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2453 a_43262_71190# a_18546_71232# a_43170_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24530 a_32126_10902# a_18162_10496# a_32218_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24531 vcm a_18162_22544# a_39246_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24532 a_22086_71190# pmat.row_n[15] a_22578_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24533 a_43170_59142# a_18162_59182# a_43262_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24534 a_20051_32521# a_19605_32149# a_19955_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24535 a_37945_28879# a_18563_27791# a_28812_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24536 a_43262_20536# a_18546_20534# a_43170_20942# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24537 a_12265_49551# a_12002_49917# a_11852_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24538 VDD pmat.rowon_n[6] a_25098_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24539 VDD a_77882_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2454 VSS a_45119_32661# a_45673_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X24540 a_11797_65871# a_11883_62063# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24541 a_39246_10496# a_18546_10494# a_39154_10902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24542 VDD a_4123_16042# a_3367_14906# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X24543 a_46578_69222# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24544 VDD a_78802_40202# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_0.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24545 VSS pmat.row_n[11] a_50594_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24546 vcm.sky130_fd_sc_hd__nand2_1_0.Y clk_vcm a_79722_40050# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24547 VSS a_12967_58559# a_12901_58633# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X24548 a_12248_42583# a_12344_42325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24549 a_25647_38695# a_21981_34191# a_25821_38571# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2455 a_19166_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24550 a_26102_70186# pmat.row_n[14] a_26594_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24551 a_47186_58138# a_18162_58178# a_47278_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24552 VSS pmat.row_n[3] a_40554_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24553 a_12581_69135# a_12067_67279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24554 a_33526_63198# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24555 VSS pmat.row_n[13] a_23486_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24556 a_20474_66210# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24557 a_13086_4175# _1194_.B1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24558 a_47186_17930# pmat.row_n[9] a_47678_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24559 VSS pmat.row_n[15] a_47582_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2456 VDD a_21219_36885# a_22325_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24560 a_51694_15484# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24561 a_50290_9492# a_18546_9490# a_50198_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24562 a_51598_21906# nmat.rowon_n[2] a_51202_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24563 VSS a_35224_50613# pmat.col[16] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X24564 a_29829_51433# a_21739_29415# pmat.col[10] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X24565 a_24186_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24566 VDD a_8560_54281# a_8735_54207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24567 a_38242_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24568 a_10515_24233# a_10513_24135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24569 a_6619_41909# a_4128_46983# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2457 VDD a_5654_9527# a_3663_9269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X24570 VSS pmat.row_n[7] a_37542_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24571 a_41558_55166# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24572 a_41558_13874# nmat.rowon_n[10] a_41162_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24573 VDD a_11421_17455# a_11711_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X24574 a_24490_65206# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24575 VDD a_13988_55369# a_14163_55295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24576 VDD a_5779_71285# a_5718_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24577 a_24586_17492# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24578 VSS a_23707_34165# a_14589_35286# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24579 a_13719_43177# a_14113_43132# a_13779_43123# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2458 a_6628_77295# a_5713_77295# a_6281_77537# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X24580 VDD a_10697_75218# a_11823_74895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24581 a_22086_18934# a_18162_18528# a_22178_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24582 a_35306_46831# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24583 a_45270_67174# a_18546_67216# a_45178_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24584 vcm a_18162_64202# a_42258_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24585 a_6337_6825# a_5935_6575# a_6173_6575# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X24586 VSS a_30857_41245# a_30549_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24587 a_42166_68178# pmat.row_n[12] a_42658_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24588 a_4553_18297# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24589 a_5463_17027# a_5271_17271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2459 a_39246_61150# a_18546_61192# a_39154_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24590 VDD a_3331_72373# a_3262_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24591 a_2847_36799# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24592 a_35138_21946# pmat.row_n[13] a_35630_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24593 a_38150_58138# pmat.row_n[2] a_38642_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24594 VSS a_2791_57703# a_4511_71631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24595 a_35138_17930# a_18162_17524# a_35230_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24596 VSS vcm.sky130_fd_sc_hd__buf_4_2.A a_77428_38962# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24597 VDD a_6087_70919# a_4396_69109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X24598 VDD pmat.rowon_n[3] a_45178_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24599 VDD a_14379_6567# a_14839_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X246 VSS ANTENNA__1197__B.DIODE nmat.col_n[31] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2460 a_6823_58951# a_6559_57167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X24600 a_12077_20291# a_11803_20535# a_11995_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24601 a_38546_11866# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24602 a_27502_56170# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24603 VSS a_3305_27791# a_6564_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24604 VSS a_14365_68743# a_12789_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24605 VDD a_6557_40545# a_6447_40669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24606 a_28602_16488# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24607 a_25098_13914# pmat.row_n[5] a_25590_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24608 a_4395_26159# a_4068_25615# a_4032_26311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24609 a_26957_39867# a_26460_40517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X2461 VDD a_13335_31359# a_13479_26935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X24610 a_40678_31599# a_26479_32117# a_40509_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24611 vcm a_18162_63198# a_46274_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24612 a_6059_44905# a_2389_45859# a_5597_44807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24613 a_46182_67174# pmat.row_n[11] a_46674_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24614 a_50690_65528# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24615 a_20752_35077# a_19689_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24616 VSS a_4123_76181# a_4985_74895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24617 a_4031_53034# a_4123_52789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24618 a_28325_27221# a_27763_27221# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24619 vcm a_18162_65206# a_19166_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2462 nmat.col_n[7] a_14458_4399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24620 a_40650_57496# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24621 a_46578_22910# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24622 a_10979_42717# a_10725_42390# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24623 a_19074_69182# pmat.row_n[13] a_19566_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24624 a_23182_63158# a_18546_63200# a_23090_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24625 vcm a_18162_60186# a_20170_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24626 VSS pmat.row_n[12] a_50594_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24627 a_1846_61651# a_2124_61635# a_2080_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24628 a_23582_67536# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24629 a_20078_64162# pmat.row_n[8] a_20570_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2463 VDD a_31015_29111# a_30603_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X24630 vcm a_18162_15516# a_37238_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24631 a_41254_13508# a_18546_13506# a_41162_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24632 a_2295_45577# a_1849_45205# a_2199_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24633 a_4496_14013# a_4379_13818# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24634 a_33130_63158# pmat.row_n[7] a_33622_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24635 a_50290_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24636 VSS pmat.row_n[4] a_40554_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24637 VSS pmat.row_n[14] a_23486_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24638 VSS a_1586_18231# a_1591_23445# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24639 VDD a_28281_41245# a_27887_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2464 a_33130_21946# a_18162_21540# a_33222_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24640 VSS a_4032_26311# a_2191_25045# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24641 VDD pmat.rowon_n[0] a_30118_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24642 VDD a_13479_26935# a_13437_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24643 VSS VDD a_48586_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24644 a_9217_28879# a_2952_25045# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24645 a_31783_42689# a_24833_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24646 a_49590_9858# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24647 a_43170_22950# a_18162_22544# a_43262_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24648 VDD a_12559_51325# a_12520_51451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24649 a_2250_31965# a_2124_31867# a_1846_31851# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2465 VDD pmat.rowon_n[7] a_43170_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X24650 a_12967_12863# a_12792_12937# a_13146_12925# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24651 a_42562_62194# pmat.rowon_n[6] a_42166_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24652 VSS a_3484_58229# a_2944_59048# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X24653 a_25647_34343# a_25755_34343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24654 VDD a_12445_12533# a_12335_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24655 a_25494_72234# VDD a_25098_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24656 a_8928_73865# a_8013_73493# a_8581_73461# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24657 a_4542_42313# a_4149_41941# a_4432_42313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24658 VDD a_1923_69823# a_2464_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24659 vcm a_18162_20536# a_32218_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2466 a_7369_19407# a_3688_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X24660 a_2163_31741# a_2046_30184# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24661 vcm a_18162_10496# a_28202_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24662 a_1757_43029# a_1591_43029# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24663 VDD a_7299_58951# a_7257_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24664 vcm a_18162_57174# a_40250_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24665 a_2012_64061# a_1895_63866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24666 a_39550_60186# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24667 a_39550_19898# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24668 a_2834_23439# a_1757_23445# a_2672_23817# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24669 a_16295_43177# a_16689_43132# a_16355_43123# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2467 VDD a_16689_43132# a_16295_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X24670 a_41162_70186# a_18162_70226# a_41254_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24671 a_40554_14878# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24672 a_23486_24918# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24673 a_79368_40202# vcm.sky130_fd_sc_hd__nand2_1_0.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24674 a_4313_44111# a_2659_35015# a_4241_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24675 VDD a_25997_42902# a_25061_43132# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X24676 a_44666_71552# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24677 a_28591_36519# a_28431_34735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24678 a_12237_38772# a_12543_39126# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24679 VDD pmat.rowoff_n[12] a_44174_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2468 a_9217_49257# a_7373_49007# a_9135_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24680 a_2439_13889# a_3571_13627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24681 a_19470_63198# pmat.rowon_n[7] a_19074_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24682 a_41600_27247# ANTENNA__1395__A1.DIODE a_41297_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24683 a_44174_61150# a_18162_61190# a_44266_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24684 a_27106_71190# a_18162_71230# a_27198_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24685 VDD a_14347_69831# a_12719_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X24686 VSS pmat.row_n[10] a_29510_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24687 VDD pmat.rowoff_n[4] a_34134_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24688 a_33526_16886# nmat.rowon_n[7] a_33130_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24689 vcm a_18162_68218# a_21174_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2469 a_8996_63695# a_8782_63695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24690 a_9303_22351# a_8859_22467# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X24691 a_11681_35823# a_11255_35862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24692 VDD pmat.rowon_n[15] a_21082_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24693 a_48682_70548# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24694 vcm a_18162_67214# a_34226_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24695 VSS config_1_in[3] a_1591_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X24696 a_45270_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24697 a_19689_38053# a_19233_38215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X24698 a_21174_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24699 VSS a_3793_47479# a_3799_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X247 a_51598_63198# pmat.rowon_n[7] a_51202_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2470 a_7436_60039# a_5682_56311# a_7578_60214# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X24700 a_45574_69222# pmat.rowon_n[13] a_45178_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24701 VSS pmat.row_n[10] a_42562_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24702 a_34226_55126# a_18546_55168# a_34134_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24703 VSS a_36617_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X24704 VDD ANTENNA__1195__A1.DIODE a_45837_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24705 a_34626_59504# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24706 a_34816_34191# a_34639_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24707 VSS a_4520_60975# a_4220_62037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24708 VDD pmat.rowon_n[14] a_25098_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24709 a_18799_51843# a_13091_52047# a_18703_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2471 a_6835_14735# a_6853_14967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X24710 VDD nmat.rowon_n[15] a_43170_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24711 VSS a_4068_25615# a_9137_27253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24712 a_3175_72641# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24713 a_8206_26703# a_7840_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24714 a_25190_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24715 a_49590_68218# pmat.rowon_n[12] a_49194_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24716 VSS pmat.row_n[9] a_46578_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24717 VDD nmat.rowon_n[6] a_46182_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24718 VDD nmat.rowon_n[15] a_19074_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24719 VSS a_12447_16143# a_14287_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2472 VSS a_16025_29469# a_16131_29429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X24720 a_44266_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24721 a_11497_40719# a_11071_41046# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24722 a_31122_8894# pmat.row_n[0] a_31614_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24723 VSS a_31793_41570# a_30857_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X24724 a_30255_49783# ANTENNA__1187__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24725 a_25042_31055# a_25084_31287# a_25042_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24726 VSS pmat.row_n[1] a_36538_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24727 a_30549_41605# a_30857_41245# a_30523_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X24728 a_25494_8854# nmat.rowon_n[15] a_25098_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24729 a_40554_55166# VSS a_40158_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2473 VDD a_13561_42333# a_13167_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X24730 a_13185_2473# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24731 a_29367_35831# a_28245_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24732 VSS pmat.row_n[11] a_19470_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24733 vcm a_18162_18528# a_29206_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24734 a_23741_42567# a_22817_41317# a_23880_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X24735 a_23486_65206# pmat.rowon_n[9] a_23090_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24736 VSS pmat.row_n[0] a_49590_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24737 VSS a_11203_62037# a_11115_71285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24738 a_33222_16520# a_18546_16518# a_33130_16926# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24739 vcm a_18162_13508# a_30210_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2474 VSS pmat.row_n[1] a_25494_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X24740 a_51294_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24741 a_6904_40303# a_5989_40303# a_6557_40545# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24742 a_47678_13476# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24743 a_37238_66170# a_18546_66212# a_37146_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24744 VDD a_2672_33775# a_2847_33749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24745 VDD nmat.rowon_n[12] a_51202_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24746 VDD nmat.rowon_n[4] a_37146_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24747 VDD a_1957_43567# a_11848_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24748 a_10529_77295# a_10494_77547# a_10291_77269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24749 VDD pmat.rowon_n[12] a_41162_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2475 VDD a_11927_27399# a_14691_27399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X24750 a_12353_16609# a_12135_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24751 a_17141_52521# a_16800_47213# a_17046_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24752 a_8378_63827# a_8695_63937# a_8653_64061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24753 a_41558_63198# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24754 VSS a_5223_11079# a_5012_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X24755 VDD pmat.rowon_n[7] a_19074_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24756 a_26498_56170# pmat.rowon_n[0] a_26102_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24757 vcm a_18162_72234# a_42258_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24758 a_10379_8439# a_9668_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24759 a_34924_36165# a_33765_35877# a_34828_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2476 VSS a_2007_25597# a_22977_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X24760 vcm a_18162_62194# a_38242_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24761 VSS a_17739_50871# a_17163_50857# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X24762 a_38150_66170# pmat.row_n[10] a_38642_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24763 a_42258_60146# a_18546_60188# a_42166_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24764 VDD pmat.rowon_n[11] a_45178_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24765 a_42658_64524# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24766 a_32162_34191# a_31985_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24767 a_27198_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24768 a_22578_7452# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24769 a_45270_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2477 VSS a_11921_35286# a_10985_35516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X24770 VDD a_42769_50069# pmat.col_n[23] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24771 VSS pmat.row_n[6] a_31518_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24772 a_7578_59887# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24773 VDD a_8264_11703# a_7283_11484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24774 a_28202_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24775 a_40694_46287# a_40645_46519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24776 a_45574_22910# nmat.rowon_n[1] a_45178_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24777 a_2834_50461# a_1757_50095# a_2672_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24778 a_15749_28111# a_9963_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24779 a_30013_30761# a_29825_30557# a_29931_30517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2478 VDD a_5821_32929# a_5711_33053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X24780 a_32218_71190# a_18546_71232# a_32126_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24781 a_43170_60146# pmat.row_n[4] a_43662_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24782 VSS a_25209_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X24783 a_6155_49007# a_5805_49007# a_6060_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24784 VDD a_2595_13621# a_2526_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24785 VDD VSS a_32126_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24786 a_38041_30485# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24787 a_29217_41570# a_30913_42043# a_32035_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24788 VDD a_3866_57399# a_6613_65577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24789 a_11421_17455# a_10995_17782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2479 a_22527_27221# ANTENNA__1395__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X24790 a_36634_55488# pmat.en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24791 a_7385_51701# a_7167_52105# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24792 a_20078_72194# VDD a_20570_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24793 vcm a_18162_23548# a_37238_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24794 a_29825_52271# a_18243_28327# pmat.col_n[9] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24795 a_49590_21906# nmat.rowon_n[2] a_49194_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24796 a_12500_68021# a_12789_68021# a_12723_68367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24797 a_46182_12910# pmat.row_n[4] a_46674_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24798 a_20570_21508# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24799 a_19566_65528# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X248 a_30210_67174# a_18546_67216# a_30118_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2480 VDD a_31978_43439# a_33259_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24800 a_20170_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24801 a_41254_21540# a_18546_21538# a_41162_21946# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24802 VSS a_21279_48999# a_22015_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24803 VDD a_18751_53034# pmat.rowoff_n[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X24804 a_50690_10464# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24805 a_37238_11500# a_18546_11498# a_37146_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24806 a_29114_22950# pmat.row_n[14] a_29606_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24807 a_33130_71190# pmat.row_n[15] a_33622_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24808 a_19074_55126# a_18162_55166# a_19166_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24809 a_33622_20504# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2481 a_25398_47081# a_11067_64015# a_25090_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.25e+11p pd=2.65e+06u as=7.4e+11p ps=5.48e+06u w=1e+06u l=150000u
X24810 a_18143_38007# a_17021_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24811 a_33222_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24812 a_39550_13874# nmat.rowon_n[10] a_39154_13914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24813 a_34063_27791# a_24591_28327# a_33845_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24814 a_36946_34191# a_36769_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24815 VSS pmat.row_n[2] a_36538_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24816 VDD a_9463_53511# a_11834_52931# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24817 a_3514_40079# a_2839_38101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24818 VDD a_33467_46261# a_36532_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24819 a_19074_14918# pmat.row_n[6] a_19566_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2482 ANTENNA__1190__B1.DIODE a_47039_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=8
X24820 vcm a_18162_7484# a_43262_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24821 VSS pmat.row_n[12] a_19470_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24822 a_23582_12472# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24823 a_6750_70589# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24824 a_21082_13914# a_18162_13508# a_21174_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24825 a_27198_22544# a_18546_22542# a_27106_22950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24826 a_35242_30099# a_35559_30209# a_35517_30333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24827 a_41162_63158# pmat.row_n[7] a_41654_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24828 vcm a_18162_7484# a_19166_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24829 VSS pmat.row_n[3] a_51598_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2483 a_32522_61190# pmat.rowon_n[5] a_32126_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24830 a_45178_18934# pmat.row_n[10] a_45670_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24831 a_34134_12910# a_18162_12504# a_34226_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24832 a_5565_19605# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24833 a_6244_40303# a_6127_40516# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24834 VDD a_32162_34191# a_33259_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24835 VSS pmat.row_n[13] a_34530_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24836 a_29206_7484# a_18546_7482# a_29114_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24837 a_7059_64822# a_6877_64822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24838 a_10995_17782# a_9528_20407# a_10995_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24839 a_36234_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2484 a_2200_9661# a_1949_9308# a_1979_9334# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X24840 a_38546_60186# pmat.rowon_n[4] a_38150_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24841 a_6970_67191# a_7435_68021# a_7393_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24842 a_38546_19898# nmat.rowon_n[4] a_38150_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24843 a_14839_54599# a_14655_53359# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24844 VDD a_9112_65161# a_9287_65087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24845 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24846 a_49286_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24847 a_12047_14165# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24848 a_22578_18496# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24849 a_15163_32375# pmat.rowon_n[7] a_15397_32509# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2485 VSS pmat.row_n[2] a_37542_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X24850 a_40158_9898# pmat.row_n[1] a_40650_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24851 a_43262_68178# a_18546_68220# a_43170_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24852 vcm a_18162_65206# a_40250_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24853 a_12613_57141# a_13091_54447# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24854 VDD a_37497_38550# a_36561_38780# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X24855 a_35534_65206# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24856 VSS a_6975_34538# a_6127_35076# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X24857 a_35178_32182# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24858 a_40158_69182# pmat.row_n[13] a_40650_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24859 a_39246_58138# a_18546_58180# a_39154_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2486 a_11711_56079# a_10595_53361# a_11889_56399# VSS sky130_fd_pr__nfet_01v8 ad=5.07e+11p pd=5.46e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X24860 VDD a_25061_43132# a_24667_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24861 a_33130_18934# a_18162_18528# a_33222_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24862 a_4809_28577# a_4591_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24863 VSS a_3331_59317# a_3262_59343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24864 VDD a_77528_40202# a_77341_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24865 a_49194_19938# pmat.row_n[11] a_49686_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24866 VDD a_4257_34319# a_6732_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24867 VDD a_11337_25071# a_14558_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24868 VDD a_1586_33927# a_1591_38677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24869 a_25494_57174# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2487 a_25117_39141# a_23700_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X24870 vcm a_18162_10496# a_36234_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24871 a_32522_58178# pmat.rowon_n[2] a_32126_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24872 a_26594_9460# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24873 a_9485_17705# a_4976_16091# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24874 a_41254_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24875 VDD a_13804_65161# a_13979_65087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24876 a_29206_69182# a_18546_69224# a_29114_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24877 a_37238_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24878 VSS a_2957_58255# a_3484_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24879 a_26594_19500# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2488 a_44174_71190# pmat.row_n[15] a_44666_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24880 a_37739_36649# a_36617_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24881 a_7343_16042# a_7387_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24882 VDD a_4413_62037# a_4349_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24883 a_20547_47491# a_13091_52047# a_20451_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24884 VSS a_8491_47911# a_9217_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24885 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24886 VSS a_14261_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X24887 a_5221_45199# a_4745_45519# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.34e+11p pd=2.02e+06u as=0p ps=0u w=650000u l=150000u
X24888 a_44570_23914# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24889 a_6612_66933# a_3339_70759# a_7004_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X2489 a_36142_7890# a_18162_7484# a_36234_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24890 a_2215_26525# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24891 a_33309_41479# a_33489_42043# a_34611_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24892 a_38242_19532# a_18546_19530# a_38150_19938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24893 a_45270_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24894 a_4815_28879# a_3351_27249# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24895 a_12901_58633# a_11711_58261# a_12792_58633# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24896 a_51694_57496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24897 VSS a_11202_55687# a_12149_56399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24898 a_34226_63158# a_18546_63200# a_34134_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24899 VSS a_10878_58487# a_11793_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X249 VDD a_1923_53055# a_2464_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2490 VDD a_6579_29199# a_6981_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X24900 a_21082_58138# a_18162_58178# a_21174_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24901 a_34626_67536# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24902 vcm a_18162_15516# a_48282_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24903 VSS a_31339_31787# a_38759_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24904 a_10379_8439# a_9668_10651# a_10613_8573# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24905 a_1643_54965# a_1846_55123# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24906 VSS a_41475_31751# a_41427_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24907 VSS pmat.row_n[0] a_48586_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24908 a_6924_25731# a_2952_25045# a_6829_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24909 a_34134_57134# a_18162_57174# a_34226_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2491 VDD nmat.rowon_n[7] pmat.rowon_n[11] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X24910 VSS _1196_.B1 a_84028_9615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24911 a_38095_32143# a_37471_32149# a_37987_32521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24912 a_21082_17930# pmat.row_n[9] a_21574_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24913 VSS pmat.row_n[15] a_21478_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24914 VDD a_9581_56079# a_11743_55329# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24915 a_46848_52047# a_13459_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24916 VSS pmat.row_n[4] a_51598_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24917 VDD a_2289_29397# a_2237_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24918 VSS pmat.row_n[14] a_34530_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24919 a_43566_70226# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2492 VSS a_5173_9839# a_5627_12879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X24920 VDD a_2389_45859# a_4927_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X24921 VDD _1154_.X a_31117_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24922 VSS a_76962_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_5.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24923 VDD a_39125_47349# a_39015_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24924 VSS a_10985_44220# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X24925 VSS a_12693_38543# a_12228_39605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24926 a_23571_44265# a_22449_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24927 a_10995_17782# a_9441_20189# a_10923_17782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24928 a_4987_34293# a_4792_34435# a_5297_34685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24929 a_83092_13103# ANTENNA__1187__B1.DIODE a_82787_13077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X2493 VDD a_46753_41935# a_41731_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.62e+12p ps=1.524e+07u w=1e+06u l=150000u M=12
X24930 a_27502_17890# nmat.rowon_n[6] a_27106_17930# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24931 a_10058_60431# a_10049_60663# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24932 a_40554_63198# pmat.rowon_n[7] a_40158_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24933 a_25098_55126# VDD a_25590_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24934 a_25776_52271# ANTENNA__1395__A1.DIODE a_25473_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24935 nmat.col[13] a_10883_3303# a_14830_3087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24936 VSS a_5688_52423# a_4659_53738# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24937 a_11113_39747# a_33489_44219# a_34552_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X24938 a_33222_24552# a_18546_24550# a_33130_24958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24939 vcm a_18162_21540# a_30210_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2494 a_23512_44007# a_22449_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X24940 a_20535_40183# a_19413_40229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24941 VDD a_82787_26133# nmat.col_n[26] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X24942 a_29206_14512# a_18546_14510# a_29114_14918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24943 a_28202_56130# a_18546_56172# a_28110_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24944 VSS config_1_in[7] a_1591_4399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X24945 a_42617_47081# a_42024_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24946 a_11979_47068# a_11823_46973# a_12124_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24947 a_45178_7890# VDD a_45670_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24948 a_2747_74549# a_2950_74707# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24949 VDD pmat.rowon_n[2] a_32126_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2495 VDD a_27789_44743# a_28572_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X24950 VSS pmat.row_n[5] a_28506_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24951 a_25494_10862# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24952 a_2387_70483# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X24953 a_32522_11866# nmat.rowon_n[12] a_32126_11906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24954 a_47915_46506# a_47975_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X24955 VSS a_10781_42869# a_22963_42657# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24956 VDD pmat.rowon_n[15] a_19074_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24957 a_12147_24233# a_11897_21263# a_12075_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24958 a_37238_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24959 a_5361_72399# a_5521_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2496 a_48190_69182# a_18162_69222# a_48282_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24960 vcm a_18162_70226# a_38242_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24961 a_15144_35077# a_13985_34789# a_15107_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24962 a_44570_64202# pmat.rowon_n[8] a_44174_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24963 a_27502_7850# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24964 a_38642_23516# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24965 vcm a_18162_12504# a_51294_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24966 a_38242_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24967 a_42658_72556# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24968 VDD nmat.rowon_n[2] a_42166_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24969 a_9333_72105# a_9279_71829# a_8283_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2497 VDD pmat.rowon_n[6] a_47186_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X24970 a_44837_35951# a_43776_30287# a_44647_36201# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24971 a_45270_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24972 a_42166_62154# a_18162_62194# a_42258_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24973 a_34530_56170# pmat.rowon_n[0] a_34134_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24974 a_25098_72194# a_18162_72234# a_25190_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24975 VSS pmat.row_n[4] a_27502_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24976 VSS pmat.row_n[11] a_27502_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24977 a_2099_76725# a_1899_76001# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X24978 a_10955_55687# a_11743_55329# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X24979 VDD a_6619_56311# a_5730_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X2498 a_43442_30287# a_28336_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X24980 a_39154_15922# a_18162_15516# a_39246_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24981 VDD pmat.rowoff_n[4] a_45178_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24982 vcm a_18162_68218# a_32218_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24983 a_43262_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24984 VDD nmat.rowon_n[1] a_28110_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24985 a_22963_34165# a_11149_36924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24986 vcm a_18162_58178# a_28202_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24987 vcm a_18162_18528# a_50290_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24988 a_1761_11471# a_1591_11471# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X24989 a_24270_49783# a_19283_49783# a_24573_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2499 VDD a_10985_37692# a_10591_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X24990 a_32218_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24991 a_30610_7452# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24992 a_29711_47679# a_29536_47753# a_29890_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24993 a_40250_71190# a_18546_71232# a_40158_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24994 VSS a_2935_38279# a_2785_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24995 VDD a_18975_40871# a_19925_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X24996 VDD nmat.rowon_n[12] a_49194_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24997 a_36234_61150# a_18546_61192# a_36142_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24998 a_7048_23277# a_7479_22467# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X24999 VSS a_82783_53524# pmat.col[31] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X25 a_10018_47741# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X250 a_39169_48829# a_39125_48437# a_39003_48841# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2500 a_33222_59142# a_18546_59184# a_33130_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X25000 VDD pmat.rowon_n[12] a_39154_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X25001 a_19074_63158# a_18162_63198# a_19166_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X25002 a_33222_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X25003 a_10995_17455# a_10741_17782# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25004 a_30118_21946# a_18162_21540# a_30210_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X25005 a_27532_28995# a_20616_27791# a_27437_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25006 VDD pmat.rowon_n[7] a_40158_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X25007 a_29206_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X25008 a_6061_38377# a_5659_38127# a_5897_38127# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X25009 VDD a_12345_36924# a_12289_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2501 vcm a_18162_56170# a_30210_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X25010 a_13769_37782# a_13597_37571# a_13555_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25011 a_1846_56875# a_2163_56765# a_2121_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25012 a_42029_48169# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25013 a_12407_28853# a_12851_28853# a_12605_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X25014 a_3417_47919# a_3151_48285# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X25015 VSS a_7658_71543# a_7663_71317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X25016 a_19566_10464# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2502 a_46274_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2503 VDD a_7131_19407# a_7533_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2504 a_29510_18894# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2505 VDD a_2419_53351# a_3891_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X2506 VSS a_1674_57711# a_7847_56085# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2507 VSS pmat.row_n[8] a_33526_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2508 a_30514_13874# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2509 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X251 a_9827_8181# a_10047_8751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2510 a_44402_32259# a_42791_32375# a_44320_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2511 a_4789_34685# a_4227_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2512 VDD a_10515_61839# a_14655_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X2513 a_31214_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2514 a_38242_22544# a_18546_22542# a_38150_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2515 VSS a_29051_37607# a_13357_37429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2516 a_21574_71552# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2517 a_42258_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2518 a_9367_53511# a_9463_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X2519 VDD a_2499_13077# a_2199_13887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X252 a_15393_28879# a_14691_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2520 a_11885_27247# a_5351_19913# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.72e+11p pd=4.36e+06u as=0p ps=0u w=650000u l=150000u
X2521 a_21082_61150# a_18162_61190# a_21174_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2522 VSS pmat.row_n[13] a_45574_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2523 a_42562_66210# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2524 a_2944_52789# a_3111_53333# a_3069_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2525 a_11133_34427# a_10651_35507# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X2526 vcm a_18162_55166# a_34226_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2527 a_22086_8894# pmat.row_n[0] a_22578_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2528 a_40158_23954# pmat.row_n[15] a_40650_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2529 a_34134_59142# pmat.row_n[3] a_34626_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X253 a_9601_66665# a_9545_66567# a_8891_66964# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X2530 a_40158_19938# a_18162_19532# a_40250_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2531 a_37463_39095# a_37497_38550# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X2532 VDD a_4128_64391# a_8477_57141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X2533 VSS a_7109_29423# a_46043_43343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X2534 a_32618_8456# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2535 a_25590_70548# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2536 a_46274_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2537 a_43170_55126# a_18162_55166# a_43262_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2538 result_out[0] a_1644_53877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2539 VSS a_5731_58951# a_5731_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X254 VSS a_17441_40482# a_16505_40157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X2540 VSS pmat.row_n[7] a_32522_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2541 VDD a_16981_37462# a_16045_37692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X2542 a_29206_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2543 VSS a_7631_15253# a_4976_16091# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X2544 a_22482_69222# pmat.rowon_n[13] a_22086_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2545 a_2935_38279# a_2847_38975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X2546 a_46578_65206# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2547 VSS a_2195_51701# a_1823_58237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2548 a_46674_17492# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2549 a_46578_23914# pmat.rowoff_n[15] a_46182_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X255 a_26194_57134# a_18546_57176# a_26102_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2550 a_43170_14918# pmat.row_n[6] a_43662_14480# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2551 VDD a_3684_22729# a_3859_22655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2552 a_79368_40202# vcm.sky130_fd_sc_hd__nand2_1_0.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2553 VDD pmat.rowoff_n[7] a_50198_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2554 a_44174_18934# a_18162_18528# a_44266_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2555 a_2847_16127# a_2672_16201# a_3026_16189# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X2556 a_6277_32687# a_5087_32687# a_6168_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2557 a_2557_56623# a_1923_53055# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2558 a_36538_57174# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2559 VSS _1194_.A2 a_12250_4175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X256 a_6612_65845# a_3339_70759# a_7004_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2560 a_36538_15882# pmat.rowoff_n[7] a_36142_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2561 VSS VDD a_40554_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2562 a_29404_36165# a_28245_35877# a_29367_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2563 a_19470_67214# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2564 a_2080_54991# a_1643_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2565 a_45428_49007# a_45450_48695# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=0p ps=0u w=650000u l=150000u
X2566 VSS a_5043_57399# a_4720_58487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2567 a_12715_51420# a_12559_51325# a_12860_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2568 a_30155_42583# a_29627_43983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2569 a_14460_61225# a_11435_58791# a_14369_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X257 a_23090_58138# pmat.row_n[2] a_23582_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2570 a_40837_46261# a_46897_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X2571 VSS pmat.row_n[9] a_23486_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2572 a_49590_56170# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2573 a_8735_54207# a_8560_54281# a_8914_54269# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X2574 a_9037_22467# a_7693_22365# a_8941_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2575 a_51202_66170# a_18162_66210# a_51294_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2576 VDD nmat.rowon_n[6] a_23090_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2577 vcm a_18162_24552# a_38242_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2578 vcm a_18162_66210# a_37238_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2579 a_47186_13914# pmat.row_n[5] a_47678_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X258 a_25098_8894# pmat.row_n[0] a_25590_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2580 VDD a_2325_38645# a_2215_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2581 a_2199_45577# a_1849_45205# a_2104_45565# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X2582 a_21174_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2583 a_51694_11468# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2584 a_41254_64162# a_18546_64204# a_41162_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2585 a_41654_68540# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2586 a_34626_21508# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2587 a_38651_37737# a_39045_37692# a_38711_37683# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2588 a_37638_58500# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2589 a_34226_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X259 VDD pmat.rowon_n[3] a_30118_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2590 a_19746_28111# a_19611_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.035e+11p pd=9.28e+06u as=0p ps=0u w=650000u l=150000u M=2
X2591 a_14917_23983# a_14475_24233# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2592 a_9463_50877# a_9135_49257# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2593 VSS pmat.row_n[3] a_37542_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2594 VSS a_33949_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X2595 VDD _1179_.X a_36722_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X2596 VSS a_46487_47919# ANTENNA__1195__A1.DIODE VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X2597 a_29510_59182# pmat.rowon_n[3] a_29114_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2598 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2599 VSS pmat.row_n[0] a_26498_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X26 VSS pmat.row_n[8] a_30514_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X260 a_20173_32117# a_19955_32521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X2600 nmat.col[5] _1192_.A2 a_23763_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X2601 VDD a_1586_33927# a_1591_40853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2602 VDD nmat.rowon_n[7] a_27106_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2603 a_24586_13476# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2604 VSS a_12069_36341# a_24895_36341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2605 a_12543_39126# a_12585_39355# a_12543_39453# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2606 VDD nmat.rowon_n[7] pmat.rowon_n[10] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X2607 a_45270_63158# a_18546_63200# a_45178_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2608 vcm a_18162_60186# a_42258_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2609 a_45670_67536# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X261 VSS pmat.row_n[6] a_26498_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2610 VSS a_17306_28879# a_17830_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X2611 a_24937_43655# a_25209_44581# a_26331_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X2612 a_42166_64162# pmat.row_n[8] a_42658_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2613 vcm a_18162_8488# a_29206_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2614 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2615 VDD a_15420_41831# a_15324_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2616 a_35138_13914# a_18162_13508# a_35230_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2617 a_8481_10396# a_9195_7423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2618 a_3508_69135# a_3029_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X2619 a_22933_32117# a_22715_32521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X262 a_23486_11866# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2620 VSS a_8385_51727# a_10081_52299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2621 a_31518_62194# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2622 a_7436_60039# a_6175_60039# a_7578_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2623 a_11113_38659# a_13801_38779# a_14923_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2624 VSS pmat.row_n[14] a_45574_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2625 vcm a_18162_71230# a_32218_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2626 VDD pmat.rowon_n[11] a_22086_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2627 a_36234_15516# a_18546_15514# a_36142_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2628 vcm a_18162_61190# a_28202_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2629 a_17867_34473# a_16745_34427# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X263 a_12437_28585# a_12175_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u
X2630 a_18084_38341# a_18180_38341# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X2631 a_6179_65479# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X2632 a_23759_52521# _1194_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X2633 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top ctopn a_52398_39208# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=9.32e+06u as=0p ps=0u w=2e+06u l=150000u M=4
X2634 a_32618_63520# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2635 a_9375_72007# a_8919_71615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2636 a_38913_31055# a_38851_30761# a_38841_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2637 VSS a_78448_39738# a_78261_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2638 a_36142_55126# pmat.en_bit_n[0] a_36634_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2639 a_82818_69135# _1154_.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X264 a_40125_31029# a_38913_31055# a_40371_31393# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2640 a_22482_22910# nmat.rowon_n[1] a_22086_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2641 a_12128_30663# a_6927_30503# a_12270_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2642 VSS a_11837_68591# a_12500_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X2643 a_19074_65166# pmat.row_n[9] a_19566_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2644 vcm a_18162_21540# a_41254_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2645 vcm a_18162_11500# a_37238_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2646 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2647 a_17012_47349# a_16863_47428# a_17308_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2648 a_20078_60146# pmat.row_n[4] a_20570_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2649 a_9556_62973# a_6175_60039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X265 VSS a_11021_42619# a_15107_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2650 a_13804_65161# a_12723_64789# a_13457_64757# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X2651 a_12987_26159# a_8013_25615# a_12902_26159# VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X2652 a_47582_72234# VDD a_47186_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2653 a_6487_5629# a_1586_8439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2654 a_14335_16519# a_11067_16359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X2655 a_38150_24958# a_18162_24552# a_38242_24552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2656 a_5081_13103# a_2648_29397# a_4863_13077# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2657 a_36538_10862# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2658 a_42258_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2659 a_25473_52245# ANTENNA__1190__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X266 a_3267_74817# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2660 nmat.rowoff_n[2] a_14839_9295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2661 a_19470_20902# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2662 a_8477_57141# a_8749_57141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X2663 a_23479_35831# a_12309_36483# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X2664 VDD pmat.rowon_n[1] a_29114_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2665 vcm a_18162_22544# a_27198_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2666 VDD a_13917_72373# a_13807_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2667 VDD a_2007_21482# a_1895_20346# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2668 a_51598_59182# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2669 a_31214_20536# a_18546_20534# a_31122_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X267 vcm a_18162_63198# a_31214_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2670 a_45574_24918# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2671 a_44444_32233# a_44382_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X2672 a_51598_17890# nmat.rowon_n[6] a_51202_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2673 a_27198_10496# a_18546_10494# a_27106_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2674 pmat.row_n[1] a_22895_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X2675 a_34530_69222# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2676 VDD _1154_.X a_31761_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X2677 a_29510_12870# pmat.rowoff_n[4] a_29114_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2678 a_36142_72194# a_18162_72234# a_36234_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2679 VSS pmat.row_n[4] a_38546_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X268 VSS pmat.row_n[11] a_38546_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2680 VSS pmat.row_n[11] a_38546_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2681 a_26891_28327# a_44515_38645# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X2682 a_40250_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2683 a_20695_30485# a_20520_30511# a_20874_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X2684 a_7674_69135# a_7730_69109# a_7674_69455# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X2685 VDD a_13151_23957# a_11927_27399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X2686 a_35138_58138# a_18162_58178# a_35230_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2687 a_49194_71190# a_18162_71230# a_49286_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2688 VDD a_4144_15113# a_4319_15039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2689 a_48586_15882# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X269 VSS a_42462_48071# a_42322_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.2e+11p ps=2.9e+06u w=650000u l=150000u
X2690 a_22086_18934# pmat.row_n[10] a_22578_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2691 VSS VDD a_22482_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2692 a_10591_37737# a_10985_37692# a_10651_37683# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2693 a_19166_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2694 a_22332_37277# a_20605_40719# a_22111_36950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2695 a_7011_44905# a_4257_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2696 a_17902_43439# a_17725_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2697 a_33905_48463# a_33957_48437# a_20475_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X2698 VDD nmat.rowon_n[1] a_39154_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2699 a_46705_38671# a_46427_39009# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_11969_27497# a_11927_27399# a_11885_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X270 a_31122_67174# pmat.row_n[11] a_31614_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2700 vcm a_18162_58178# a_39246_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2701 VDD pmat.rowon_n[15] a_43170_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2702 a_35138_17930# pmat.row_n[9] a_35630_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2703 a_43262_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2704 VSS a_35290_44527# a_36111_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2705 a_26180_39429# a_25117_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2706 a_26194_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2707 a_5621_47081# a_5221_45199# a_5537_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X2708 a_28506_18894# nmat.rowon_n[5] a_28110_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2709 a_23191_37277# a_14712_37429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X271 a_42562_65206# pmat.rowon_n[9] a_42166_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2710 a_23759_52521# _1192_.A2 a_23541_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2711 a_20170_68178# a_18546_68220# a_20078_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2712 a_8385_51727# a_7907_52031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2713 a_2831_21807# a_2683_22089# a_2468_21959# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2714 VDD a_10814_29111# a_10763_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2715 a_41162_21946# a_18162_21540# a_41254_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2716 cgen.start_conv_in a_1591_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2717 a_39092_50639# _1183_.A2 a_38627_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2718 a_13985_40229# a_11773_39087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X2719 VDD pmat.rowon_n[14] a_47186_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X272 a_29827_39095# a_28705_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2720 vcm a_18162_69222# a_29206_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2721 a_37146_11906# a_18162_11500# a_37238_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2722 a_33222_67174# a_18546_67216# a_33130_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2723 vcm a_18162_64202# a_30210_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2724 a_26102_19938# pmat.row_n[11] a_26594_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2725 a_3300_19453# a_3183_19258# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X2726 a_30118_68178# pmat.row_n[12] a_30610_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2727 a_29206_57134# a_18546_57176# a_29114_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2728 a_41558_66210# pmat.rowon_n[10] a_41162_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2729 VSS pmat.row_n[0] a_39550_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X273 a_21032_44007# a_19873_44219# a_20995_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2730 a_37129_36130# a_36617_36603# a_37739_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2731 a_51294_17524# a_18546_17522# a_51202_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2732 VDD pmat.rowon_n[3] a_33130_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2733 a_9761_30511# a_9595_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2734 a_20425_49667# a_19584_52423# a_20353_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2735 VDD a_2319_54965# a_2250_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X2736 VSS pmat.row_n[6] a_29510_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2737 VSS comp.adc_inverter_1.out a_52398_39208# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u M=8
X2738 VDD a_11113_36483# a_20752_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2739 a_33715_48783# a_33685_48437# a_20475_49783# VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X274 a_12217_66389# a_13973_66933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X2740 VSS a_32162_34191# a_33259_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2741 a_17588_32463# a_11067_64015# a_17285_32117# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X2742 a_27519_42359# a_27913_42333# a_27329_42902# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2743 a_51202_57134# pmat.row_n[1] a_51694_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2744 a_5602_30511# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X2745 vcm a_18162_63198# a_34226_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2746 a_38546_64202# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2747 a_34134_67174# pmat.row_n[11] a_34626_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2748 a_2417_45173# a_2199_45577# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X2749 a_45574_65206# pmat.rowon_n[9] a_45178_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X275 VSS a_9195_7423# a_9129_7497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X2750 a_12226_14191# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X2751 a_21478_23914# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2752 a_82817_25935# _1224_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X2753 a_43170_63158# a_18162_63198# a_43262_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2754 a_6369_39215# a_5687_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2755 a_51598_12870# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2756 a_11071_39958# a_11041_39860# a_10999_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2757 a_35534_57174# pmat.rowon_n[1] a_35138_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2758 a_3514_57167# a_1591_56623# a_3431_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X2759 VDD a_6634_26133# a_6829_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X276 a_36453_29199# a_7717_14735# a_36465_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2760 a_8213_53877# a_7995_54281# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X2761 a_34530_22910# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2762 VDD a_1923_61759# a_3207_65845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2763 VDD a_2325_20149# a_2215_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2764 a_28202_18528# a_18546_18526# a_28110_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2765 a_4128_64391# a_6343_32661# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2766 a_3615_71631# a_11071_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X2767 a_4193_66237# a_3814_65871# a_4121_66237# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X2768 a_6541_15279# a_6375_15279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2769 vcm a_18162_15516# a_25190_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X277 VSS a_20316_47607# a_20267_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2770 VDD nmat.rowon_n[15] a_42166_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2771 a_14287_59887# a_10239_14183# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X2772 a_48586_56170# pmat.rowon_n[0] a_48190_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2773 VDD nmat.rowon_n[10] a_46182_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2774 a_6521_71017# a_3339_70759# a_6087_70919# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X2775 VDD a_3423_74549# a_3354_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X2776 VDD a_7896_11079# a_7276_11739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2777 a_5825_22901# nmat.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X2778 VSS pmat.row_n[7] a_40554_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2779 a_12429_62607# a_12081_62723# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X278 a_40158_63158# a_18162_63198# a_40250_63158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2780 a_46921_30761# a_43776_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2781 a_34887_41271# a_34924_41605# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X2782 nmat.col[23] _1154_.X a_41786_28111# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X2783 VSS a_30699_29397# a_29455_31293# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2784 VDD a_41731_49525# a_24407_31375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X2785 a_45505_31599# a_45119_32661# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X2786 a_20474_70226# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2787 a_8091_49192# a_7373_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2788 a_12135_16367# a_11785_16367# a_12040_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X2789 VSS a_34942_51701# a_37092_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X279 a_49686_23516# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2790 a_20572_40517# a_19413_40229# a_20535_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2791 a_24490_8854# nmat.rowon_n[15] a_24094_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2792 a_50594_18894# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2793 VSS a_9135_60967# a_9335_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X2794 vcm a_18162_14512# a_29206_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2795 a_2781_26159# a_1591_26159# a_2672_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2796 a_41254_72194# a_18546_72236# a_41162_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2797 a_14347_69831# a_3615_71631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2798 a_37238_62154# a_18546_62196# a_37146_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2799 VDD a_4339_27804# a_7803_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X28 a_18243_28327# a_45589_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u M=4
X280 a_49286_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2800 a_37638_66532# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2801 a_10286_60405# a_9135_60967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X2802 VDD pmat.rowon_n[8] a_41162_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2803 result_out[11] a_1644_70197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2804 a_45563_31055# a_30571_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X2805 VSS a_24719_35253# a_11921_35286# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2806 a_37146_56130# a_18162_56170# a_37238_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2807 a_23486_61190# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2808 a_40158_8894# a_18162_8488# a_40250_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2809 VDD a_4583_68021# a_9139_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X281 a_3408_11849# a_2493_11477# a_3061_11445# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X2810 a_30514_62194# pmat.rowon_n[6] a_30118_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2811 VDD cgen.dlycontrol3_in[3] a_25755_38695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2812 VSS a_8013_25615# a_14287_24349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X2813 VDD a_3983_43567# a_2315_44124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X2814 a_42166_72194# VDD a_42658_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2815 VSS a_4976_16091# a_10151_19637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X2816 a_8547_77129# a_8031_76757# a_8452_77117# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X2817 a_38150_62154# pmat.row_n[6] a_38642_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2818 a_44933_35951# a_43533_30761# a_44837_35951# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X2819 VDD a_14071_8511# a_14058_8207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X282 VSS a_12585_39355# a_27795_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2820 a_42658_60508# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2821 VSS a_9367_50871# a_9319_50639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2822 a_33684_32143# a_33205_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X2823 a_26194_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2824 a_27502_60186# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2825 a_27502_19898# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2826 a_21574_7452# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2827 VDD a_20503_48981# pmat.row_n[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2828 VSS a_3496_51701# a_3434_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X2829 VDD a_5363_33551# a_14287_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X283 a_31518_22910# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2830 a_2012_28157# a_1895_27962# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2831 VDD a_11142_64783# a_11019_71543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2832 a_9335_58575# a_9577_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X2833 VDD pmat.en_bit_n[2] a_35138_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2834 VSS a_12895_53359# a_13181_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X2835 VDD a_24895_43957# a_24719_43957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X2836 a_36234_23548# a_18546_23546# a_36142_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2837 a_28725_52271# a_18243_28327# a_28507_52245# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2838 a_45670_12472# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2839 VSS a_32256_44869# a_32219_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X284 VDD _1179_.X a_83178_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X2840 VDD VDD a_31122_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2841 a_45915_29941# a_46723_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2842 VSS a_1586_18231# a_4075_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2843 a_28602_22512# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2844 a_32618_71552# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2845 a_40554_67214# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2846 a_49286_22544# a_18546_22542# a_49194_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2847 a_18162_55166# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X2848 VDD pmat.rowoff_n[12] a_32126_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2849 VSS a_15049_42902# a_14113_43132# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X285 a_25190_18528# a_18546_18526# a_25098_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2850 a_40685_50639# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X2851 a_32126_61150# a_18162_61190# a_32218_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2852 a_35534_10862# nmat.rowon_n[13] a_35138_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2853 a_18243_31599# a_14691_27399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X2854 VDD pmat.rowoff_n[4] a_22086_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2855 VSS a_33765_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X2856 vcm a_18162_61190# a_36234_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2857 a_20170_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2858 VDD a_16083_50069# a_18583_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2859 a_40650_63520# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X286 a_26497_36603# a_26041_36374# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X2860 pmat.col_n[29] _1194_.A2 a_46109_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2861 a_29114_14918# a_18162_14512# a_29206_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2862 a_21377_27497# a_11927_27399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2863 a_28273_28879# a_15667_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X2864 a_30103_43447# a_28981_43493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2865 a_50594_59182# pmat.rowon_n[3] a_50198_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2866 a_1849_45205# a_1683_45205# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2867 a_18546_72236# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X2868 a_44666_18496# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2869 a_12471_36950# a_12289_36950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X287 vcm a_18162_15516# a_22178_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2870 a_33222_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2871 VDD a_39496_30199# a_39497_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2872 a_33526_69222# pmat.rowon_n[13] a_33130_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2873 VSS a_25695_28111# a_35621_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X2874 a_19074_10902# pmat.row_n[2] a_19566_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2875 a_13427_74953# a_12981_74581# a_13331_74953# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X2876 vcm a_18162_7484# a_42258_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2877 VSS a_78448_40202# a_78261_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2878 VDD a_42240_29423# a_43913_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2879 a_1642_20871# a_1738_20693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X288 a_4553_28089# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2880 a_3024_22717# a_2907_22522# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2881 a_28116_38567# a_26957_38779# a_28079_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X2882 a_47582_57174# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2883 VSS VDD a_51598_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X2884 VDD nmat.rowon_n[5] a_21082_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2885 a_36541_29673# a_36453_29199# a_36459_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=1.87e+12p ps=1.774e+07u w=1e+06u l=150000u
X2886 VSS a_1899_35051# a_6403_37252# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2887 a_45047_38155# a_44444_32233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2888 VSS pmat.row_n[9] a_34530_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2889 vcm a_18162_66210# a_48282_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X289 a_45574_56170# pmat.rowon_n[0] a_45178_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2890 VDD a_31469_40726# a_31976_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2891 a_32218_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2892 a_27789_36039# a_27049_35515# a_28171_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2893 a_28202_7484# a_18546_7482# a_28110_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2894 a_48682_19500# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2895 VDD a_7589_33749# a_7619_34102# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2896 a_38627_50613# a_38770_50755# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2897 VSS a_15439_48071# a_14528_48114# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X2898 VSS a_11149_36924# a_22963_34165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2899 a_22086_69182# a_18162_69222# a_22178_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X29 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u M=33
X290 a_39646_15484# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2900 VSS pmat.row_n[1] a_24490_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2901 a_35230_10496# a_18546_10494# a_35138_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2902 VDD a_40837_46261# a_46753_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X2903 vcm a_18162_9492# a_33222_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2904 a_11575_18870# a_5351_19913# a_11116_18695# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X2905 a_27605_37127# a_26497_36603# a_27560_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2906 a_20316_47607# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2907 a_7657_22467# a_4703_24527# a_7561_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2908 a_12081_62723# a_12199_62621# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2909 a_40158_65166# pmat.row_n[9] a_40650_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X291 a_24719_43957# a_24895_43957# a_24847_43983# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X2910 VSS a_5423_30485# a_5357_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2911 a_44855_45199# a_43720_32143# a_44737_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X2912 VDD nmat.rowon_n[4] a_25098_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2913 a_5749_30265# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2914 a_12981_8213# a_12815_8213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2915 a_26102_68178# a_18162_68218# a_26194_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2916 VSS a_12047_14165# a_11981_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X2917 VDD a_8013_25615# a_14287_24349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2918 a_1775_47375# a_1769_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X2919 VSS pmat.row_n[15] a_43566_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X292 VDD nmat.rowon_n[10] a_43170_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2920 VDD a_9368_9991# a_8472_11739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2921 a_40554_20902# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2922 a_25590_9460# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2923 vcm a_18162_72234# a_30210_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2924 a_43170_56130# pmat.row_n[0] a_43662_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2925 a_29206_65166# a_18546_65208# a_29114_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2926 VDD pmat.rowon_n[1] a_50198_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2927 a_29606_69544# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2928 a_20627_38825# a_19505_38779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2929 a_20170_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X293 a_28506_66210# pmat.rowon_n[10] a_28110_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2930 VDD a_14917_23983# a_18243_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2931 VDD pmat.rowon_n[11] a_33130_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2932 a_4041_61225# a_4081_61127# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X2933 a_47278_15516# a_18546_15514# a_47186_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2934 a_29114_59142# a_18162_59182# a_29206_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2935 VSS a_2835_13077# a_11569_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2936 a_33222_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2937 VDD a_1643_52789# a_1591_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2938 a_49590_17890# nmat.rowon_n[6] a_49194_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2939 a_20570_17492# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X294 VSS a_14287_70543# a_14839_69135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2940 a_20474_23914# pmat.rowoff_n[15] a_20078_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2941 VDD a_23329_37462# a_23788_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2942 a_11067_16359# a_18487_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X2943 a_2847_23743# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2944 VDD a_4037_69109# a_2944_69928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2945 a_50594_12870# pmat.rowoff_n[4] a_50198_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2946 VSS a_18869_46831# a_19474_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2947 a_38546_72234# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2948 a_47186_55126# VDD a_47678_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2949 VSS config_2_in[1] a_1591_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X295 VDD pmat.rowoff_n[15] a_26102_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2950 a_17559_51157# a_17033_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X2951 a_10141_60431# a_10286_60405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X2952 a_33526_22910# nmat.rowon_n[1] a_33130_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2953 VSS pmat.row_n[14] a_42562_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2954 a_31122_21946# pmat.row_n[13] a_31614_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2955 VDD a_43776_30287# a_44449_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2956 VDD a_43533_30761# a_46921_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2957 a_5253_11177# a_5363_12015# a_5445_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2958 a_31122_17930# a_18162_17524# a_31214_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2959 a_26957_39867# a_26460_40517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X296 VDD a_5597_44807# a_5566_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.35e+11p ps=2.67e+06u w=1e+06u l=150000u
X2960 a_6244_71829# a_3339_70759# a_6636_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2961 VDD a_15368_31599# a_15543_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2962 a_10379_8439# a_10378_7637# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X2963 vcm a_18162_11500# a_48282_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2964 a_5747_44655# a_5921_44629# VSS VSS sky130_fd_pr__nfet_01v8 ad=6.565e+11p pd=5.92e+06u as=0p ps=0u w=650000u l=150000u
X2965 VDD a_14113_36604# a_13719_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2966 VSS a_4553_18297# a_4487_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2967 a_10975_62313# a_10190_60663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X2968 VSS a_17139_30503# a_25505_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2969 VSS a_10515_13967# a_20175_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X297 a_39359_49172# a_38793_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2970 a_21082_13914# pmat.row_n[5] a_21574_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2971 a_47582_10862# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2972 a_4291_48169# a_3417_47919# a_4071_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X2973 a_24586_55488# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2974 vcm a_18162_23548# a_25190_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2975 VDD a_12447_16143# a_14011_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2976 a_34134_12910# pmat.row_n[4] a_34626_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2977 a_12715_51420# a_12520_51451# a_13025_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X2978 nmat.col_n[21] a_82787_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2979 a_33130_9898# a_18162_9492# a_33222_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X298 a_2672_28169# a_1591_27797# a_2325_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X2980 a_12020_40871# a_12228_40693# a_12162_40719# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2981 VSS a_27001_30511# a_27995_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.3585e+12p ps=1.328e+07u w=650000u l=150000u M=4
X2982 a_18546_10494# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X2983 VDD a_12449_39605# a_12479_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2984 a_7747_25731# a_7186_25615# a_7665_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2985 VSS a_1586_18231# a_1591_27797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2986 VDD a_25647_39783# a_11339_39319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X2987 a_4509_24643# a_3305_27791# a_4437_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2988 a_27502_13874# nmat.rowon_n[10] a_27106_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2989 VDD a_5047_76983# a_4951_76983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X299 VSS a_12147_24233# a_8583_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X2990 vcm a_18162_69222# a_50290_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2991 VSS pmat.row_n[2] a_24490_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2992 VSS a_11545_18517# a_11479_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2993 VDD a_2244_26935# a_2021_26677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2994 a_47186_72194# a_18162_72234# a_47278_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2995 VSS pmat.row_n[4] a_49590_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2996 a_6700_57863# a_4843_54826# a_6842_57711# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2997 a_11337_25071# a_5991_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=2
X2998 VSS pmat.row_n[11] a_49590_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2999 a_6323_26409# a_6634_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.96e+12p pd=1.792e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3 a_41162_71190# pmat.row_n[15] a_41654_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X30 VDD nmat.rowon_n[7] nmat.rowoff_n[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X300 a_41968_46831# a_41926_46983# a_41665_46805# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3000 a_51294_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3001 VSS a_29711_47679# a_29076_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3002 a_39550_66210# pmat.rowon_n[10] a_39154_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3003 a_4337_22351# a_3859_22655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3004 a_37238_70186# a_18546_70228# a_37146_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3005 VDD a_6830_22895# a_12461_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X3006 VDD a_1923_69823# a_1643_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3007 VDD pmat.rowoff_n[15] a_37146_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3008 a_50290_12504# a_18546_12502# a_50198_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3009 VDD VDD a_41162_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X301 a_5320_57863# a_5528_57685# a_5462_57711# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3010 a_33130_18934# pmat.row_n[10] a_33622_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3011 a_2080_67869# a_1643_67477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3012 a_13103_26703# a_12987_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X3013 a_49194_8894# a_18162_8488# a_49286_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3014 a_37146_64162# a_18162_64202# a_37238_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3015 a_44174_7890# VDD a_44666_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3016 a_41254_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3017 a_1687_13621# a_2122_13779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3018 a_26456_38341# a_26501_37462# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3019 a_24186_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X302 VSS pmat.row_n[6] a_50594_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3020 a_26498_60186# pmat.rowon_n[4] a_26102_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3021 VSS a_33489_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3022 a_38546_7850# VDD a_38150_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3023 a_26498_19898# nmat.rowon_n[4] a_26102_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3024 a_50594_7850# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3025 VSS a_25393_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3026 a_38150_70186# pmat.row_n[14] a_38642_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3027 a_38242_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3028 a_39111_38825# a_22153_37179# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X3029 a_26498_7850# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X303 vcm a_18162_14512# a_26194_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3030 a_41665_46805# a_13275_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3031 a_31214_68178# a_18546_68220# a_31122_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3032 a_18751_53034# a_18777_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3033 a_27198_58138# a_18546_58180# a_27106_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3034 VSS pmat.row_n[1] a_19470_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3035 a_3045_19093# a_2879_19093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3036 a_48190_11906# a_18162_11500# a_48282_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3037 a_11229_72943# a_10751_72917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3038 a_2957_58255# a_2603_58368# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3039 a_2122_19087# a_1945_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X304 a_49590_55166# VSS a_49194_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3040 a_27757_43439# a_11497_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3041 a_10149_57961# a_10090_58093# a_10054_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X3042 a_34425_50639# a_28915_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.95e+11p pd=5.19e+06u as=0p ps=0u w=1e+06u l=150000u
X3043 vcm a_18162_10496# a_24186_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3044 a_41637_31599# a_39939_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X3045 a_18162_63198# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X3046 VSS pmat.row_n[12] a_39550_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3047 vcm a_18162_19532# a_49286_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3048 VSS a_1687_13621# a_1717_13647# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3049 a_5065_63669# a_5357_62779# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X305 VSS a_11261_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3050 a_2557_31599# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X3051 a_40352_41831# a_39193_42043# a_40315_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3052 a_36571_44527# a_36394_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3053 vcm a_18162_14512# a_50290_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3054 a_11275_36950# a_11093_36950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X3055 a_2319_69916# a_2124_69947# a_2629_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X3056 VSS a_2129_12559# a_3158_13647# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3057 a_16339_43745# a_12069_38517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3058 VDD a_20695_30485# a_20682_30877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3059 a_21037_43658# cgen.start_conv_in VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X306 VSS VDD a_33526_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3060 a_8333_24847# a_6173_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X3061 VSS a_4719_30287# a_5465_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3062 a_10383_75637# a_9581_73487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3063 a_50290_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3064 a_40650_71552# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3065 a_32522_23914# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3066 a_11990_73309# a_11271_73085# a_11427_73180# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X3067 a_29114_22950# a_18162_22544# a_29206_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3068 VDD pmat.rowon_n[8] a_39154_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3069 a_36634_61512# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X307 a_12489_12925# a_12445_12533# a_12323_12937# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3070 a_26194_19532# a_18546_19530# a_26102_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3071 a_33222_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3072 a_44266_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3073 VDD a_2163_67645# a_2124_67771# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3074 vcm a_18162_16520# a_23182_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3075 VDD a_54790_39198# comp.adc_nor_latch_0.R VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u M=2
X3076 a_46578_57174# pmat.rowon_n[1] a_46182_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3077 a_30549_41605# a_30523_41245# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3078 a_2847_50069# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3079 a_44927_43567# a_7109_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=0p ps=0u w=650000u l=150000u
X308 a_46263_52245# _1194_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X3080 a_22482_15882# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3081 VSS pmat.row_n[10] a_25494_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3082 a_33341_43777# a_24833_40719# a_33255_43777# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3083 VDD a_5547_14735# a_2648_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X3084 a_13145_26935# a_13683_24847# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.654e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3085 VSS a_40837_46261# a_25879_31591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X3086 VSS a_46339_31029# _1194_.B1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=8
X3087 a_45719_36495# a_35244_32411# a_45625_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X3088 VSS pmat.row_n[7] a_51598_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3089 a_48282_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X309 VDD pmat.rowon_n[13] a_37146_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3090 VSS a_27877_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3091 vcm a_18162_57174# a_26194_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3092 VSS a_31879_34191# a_31985_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3093 a_30210_55126# a_18546_55168# a_30118_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3094 a_11711_60751# a_5651_66975# a_12155_60751# VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=1.6185e+12p ps=1.668e+07u w=650000u l=150000u M=4
X3095 VDD a_4227_34293# a_4257_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3096 VDD a_5363_70543# a_14749_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3097 a_30610_59504# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3098 VSS a_44444_32233# a_47685_30517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3099 a_26498_14878# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u M=887
X310 a_83839_9295# ANTENNA__1190__A1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X3100 a_12335_58255# a_11711_58261# a_12227_58633# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3101 a_45178_24958# VDD a_45670_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3102 a_13427_8585# a_12981_8213# a_13331_8585# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X3103 a_27687_34967# cgen.dlycontrol1_in[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3104 a_17702_29967# a_12461_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3105 VDD pmat.sample_n a_18162_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X3106 a_48190_56130# a_18162_56170# a_48282_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3107 a_23455_32447# a_2007_25597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3108 a_1644_70197# a_1591_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3109 a_29864_39429# a_28705_39141# a_29827_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X311 a_51294_71190# a_18546_71232# a_51202_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3110 VSS a_37497_38550# a_36561_38780# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X3111 a_11071_38870# a_11041_38772# a_10999_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3112 VDD nmat.rowon_n[6] a_42166_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3113 a_31303_27497# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X3114 a_40250_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3115 a_43262_9492# a_18546_9490# a_43170_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3116 a_24719_38517# a_24895_38517# a_24847_38543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X3117 a_22578_24520# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3118 a_49194_23954# pmat.row_n[15] a_49686_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3119 a_44571_32143# a_44320_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X312 a_27198_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3120 a_49194_19938# a_18162_19532# a_49286_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3121 VDD a_9427_50095# a_9367_50871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3122 a_50198_14918# a_18162_14512# a_50290_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3123 VSS a_16377_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3124 a_14441_57533# a_10515_13967# a_14369_57533# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3125 VDD a_13479_26935# a_14833_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X3126 VSS a_5123_52423# a_5081_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X3127 a_4259_70767# a_2727_58470# a_4165_70767# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X3128 a_39015_48463# a_38391_48469# a_38907_48841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3129 VSS pmat.row_n[0] a_45574_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X313 a_47278_61150# a_18546_61192# a_47186_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3130 a_39154_15922# pmat.row_n[7] a_39646_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3131 a_14648_4175# ANTENNA__1183__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3132 VSS pmat.row_n[13] a_39550_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3133 a_43662_13476# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3134 a_40158_10902# pmat.row_n[2] a_40650_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3135 VSS a_39045_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3136 VSS pmat.row_n[10] a_28506_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3137 VDD a_15839_49525# a_10515_15055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3138 VSS a_11261_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3139 a_28721_47081# a_11067_49871# a_28639_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X314 a_20474_61190# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3140 a_32522_64202# pmat.rowon_n[8] a_32126_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3141 VDD VSS a_46182_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3142 a_23090_20942# pmat.row_n[12] a_23582_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3143 a_26594_23516# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3144 a_26194_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3145 VSS a_25647_38695# a_18975_40871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3146 pmat.col[8] a_28131_50069# a_27903_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X3147 a_23090_16926# a_18162_16520# a_23182_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3148 a_47278_23548# a_18546_23546# a_47186_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3149 VSS a_21219_36885# a_22332_37277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X315 VDD pmat.rowon_n[7] a_51202_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3150 a_7289_37039# a_6099_37039# a_7180_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X3151 VDD nmat.rowon_n[2] a_30118_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3152 a_33222_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3153 a_30118_62154# a_18162_62194# a_30210_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3154 a_3092_59343# a_2655_59317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3155 a_29206_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3156 a_22482_56170# pmat.rowon_n[0] a_22086_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3157 VDD nmat.rowon_n[5] a_19074_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3158 VSS config_1_in[1] a_1591_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3159 a_12806_53359# a_12003_52815# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X316 nmat.rowoff_n[9] a_10515_15055# a_12990_13967# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X3160 a_5138_65479# a_5399_65479# a_5352_65577# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X3161 VSS cgen.enable_dlycontrol_in a_24667_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3162 VSS a_45019_38645# a_17139_30503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u M=8
X3163 VDD a_20855_36885# a_19233_38215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3164 a_4687_14025# a_4241_13653# a_4591_14025# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X3165 a_46578_10862# nmat.rowon_n[13] a_46182_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3166 VDD nmat.rowon_n[10] a_20078_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3167 a_6720_49007# a_5639_49007# a_6373_49249# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X3168 a_9287_65087# a_9112_65161# a_9466_65149# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3169 a_19647_48052# a_19441_47491# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X317 pmat.col[14] a_34705_51959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3170 a_29606_14480# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3171 VDD cgen.dlycontrol4_in[1] a_31095_42367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3172 vcm a_18162_71230# a_51294_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3173 VSS a_13909_39605# a_13853_39958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3174 a_9687_67075# a_9405_66627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3175 a_27106_15922# a_18162_15516# a_27198_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3176 VDD pmat.rowoff_n[4] a_33130_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3177 vcm a_18162_61190# a_47278_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3178 a_31214_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3179 VSS a_2897_21781# a_2831_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 VDD a_2944_61493# a_2882_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X3180 a_24407_31375# a_41731_49525# a_44423_36815# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X3181 a_51694_63520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3182 VSS a_4075_31591# a_14633_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X3183 VDD a_26475_34343# a_11057_35836# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X3184 vcm a_18162_8488# a_22178_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3185 a_4895_12559# a_4865_12533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3186 a_30957_48169# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3187 VSS a_82788_10357# nmat.col_n[24] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X3188 a_45574_58178# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3189 a_24186_61150# a_18546_61192# a_24094_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X319 VDD a_12245_21807# a_12271_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3190 ndecision_finish comp.adc_nor_latch_0.NOR_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3191 VDD a_1586_8439# a_6375_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3192 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3193 a_8649_18115# a_7644_16341# a_8577_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3194 VDD pmat.rowon_n[12] a_27106_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3195 a_28506_68218# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3196 a_32218_8488# a_18546_8486# a_32126_8894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3197 a_11785_16367# a_11619_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3198 a_4995_52815# a_2315_44124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3199 a_33685_48437# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X32 a_49194_9898# pmat.row_n[1] a_49686_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X320 VDD a_2411_43301# a_4984_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X3200 a_13979_65087# a_13804_65161# a_14158_65149# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3201 a_43262_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3202 a_2847_43327# a_2672_43401# a_3026_43389# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3203 a_18546_69224# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3204 VSS a_18243_28327# a_44268_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3205 VSS a_3615_71631# a_13966_71631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X3206 VDD a_20475_49783# a_20517_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3207 a_6564_24527# a_5991_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.225e+11p pd=3.9e+06u as=0p ps=0u w=650000u l=150000u
X3208 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3209 a_11071_38543# a_10817_38870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X321 pmat.rowon_n[14] a_14839_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3210 a_25879_31591# a_44763_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3211 VSS pmat.row_n[2] a_22482_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3212 VSS pmat.row_n[15] a_36538_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3213 pmat.rowon_n[8] nmat.rowon_n[7] a_13686_13967# VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=1.2675e+12p ps=1.3e+07u w=650000u l=150000u M=4
X3214 a_50198_59142# a_18162_59182# a_50290_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3215 vcm a_18162_22544# a_46274_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3216 a_28202_60146# a_18546_60188# a_28110_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3217 VDD a_10378_7637# a_10747_6727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3218 a_28602_64524# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3219 a_19615_41959# a_12658_42895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X322 a_1643_67477# a_1846_67755# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3220 a_25098_61150# pmat.row_n[5] a_25590_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3221 a_50290_20536# a_18546_20534# a_50198_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3222 a_5688_52423# a_5731_58951# a_5919_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3223 a_33130_69182# a_18162_69222# a_33222_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3224 VSS a_33765_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3225 VDD pmat.rowon_n[6] a_32126_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3226 a_46274_10496# a_18546_10494# a_46182_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3227 a_37238_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3228 a_9900_32143# a_9231_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3229 a_4855_32509# a_4707_32156# a_4492_32375# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X323 a_43605_29423# a_41949_30761# a_43533_29423# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3230 pmat.rowon_n[9] a_14734_64015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3231 VDD a_41949_30761# a_42701_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X3232 a_23182_22544# a_18546_22542# a_23090_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3233 a_19166_12504# a_18546_12502# a_19074_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3234 a_24524_30287# a_22628_30485# a_24404_30287# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X3235 a_41162_18934# pmat.row_n[10] a_41654_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3236 VSS VDD a_41558_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3237 VSS a_34277_37462# a_34887_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X3238 a_29114_60146# pmat.row_n[4] a_29606_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3239 a_38242_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X324 VDD a_9441_20189# a_12311_19783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3240 a_6173_22895# a_5825_22901# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3241 a_15107_41271# a_13985_41317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3242 a_20568_38567# a_19509_39638# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3243 VSS pmat.row_n[13] a_30514_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3244 a_14371_25071# a_9441_20189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3245 a_26239_39095# a_25117_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3246 a_1957_43567# a_1927_43541# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X3247 a_34530_60186# pmat.rowon_n[4] a_34134_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3248 a_8744_71689# a_7663_71317# a_8397_71285# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X3249 a_34530_19898# nmat.rowon_n[4] a_34134_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X325 a_38642_65528# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3250 a_18769_36965# a_18180_38341# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X3251 a_18325_31599# a_18241_31698# a_18243_31599# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3252 a_13575_68743# a_3615_71631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3253 a_31214_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3254 a_23700_44869# a_22541_44581# a_23604_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3255 a_45270_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3256 a_43191_49551# a_38851_28327# a_28131_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3257 VSS pmat.row_n[7] a_44570_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3258 a_47582_18894# nmat.rowon_n[5] a_47186_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3259 a_31767_47919# a_31152_48071# a_28901_48437# VSS sky130_fd_pr__nfet_01v8 ad=7.085e+11p pd=7.38e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X326 VSS nmat.sample a_18546_19530# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X3260 a_41558_9858# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3261 VDD a_4831_34561# a_4792_34435# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3262 a_31518_65206# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3263 a_4429_37039# a_3325_36495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X3264 a_35230_58138# a_18546_58180# a_35138_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3265 a_31614_17492# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3266 a_31518_23914# pmat.rowoff_n[15] a_31122_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3267 VSS a_5955_55223# a_5904_55311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3268 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3269 VSS pmat.row_n[1] a_51598_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X327 a_40256_42919# a_39013_43655# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3270 a_48282_57134# a_18546_57176# a_48190_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3271 a_45178_58138# pmat.row_n[2] a_45670_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3272 a_21478_57174# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3273 a_21478_15882# pmat.rowoff_n[7] a_21082_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3274 a_14163_55295# a_1957_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3275 VSS pmat.row_n[6] a_48586_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3276 a_45574_11866# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3277 VSS a_3577_70197# a_2944_72104# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3278 a_4912_41935# a_4432_42313# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X3279 a_34530_56170# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 VSS comp.adc_nor_latch_0.R ndecision_finish VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3280 VDD VDD a_39154_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3281 a_28506_21906# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3282 vcm a_18162_24552# a_23182_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3283 a_25190_69182# a_18546_69224# a_25098_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3284 a_6817_21807# a_6469_21813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3285 vcm a_18162_66210# a_22178_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3286 a_32126_13914# pmat.row_n[5] a_32618_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3287 VSS a_5012_10927# a_3576_17143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.64e+11p ps=3.72e+06u w=650000u l=150000u M=4
X3288 a_7302_33775# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3289 a_2685_58621# a_1591_58799# a_2603_58368# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X329 a_3234_40553# a_3199_40455# a_2931_40277# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X3290 a_44774_40821# a_46013_42997# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3291 a_16879_50345# pmat.rowon_n[7] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3292 a_22578_58500# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3293 a_3399_24787# a_3325_23439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X3294 a_6845_13103# a_5173_9839# a_6763_13103# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3295 a_25494_14878# nmat.rowon_n[9] a_25098_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3296 a_36919_31849# a_37143_31573# a_5179_31591# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3297 VSS pmat.row_n[3] a_22482_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3298 a_6829_57487# a_6835_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X3299 a_19166_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X33 VDD nmat.rowon_n[4] a_48190_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X330 a_48190_61150# pmat.row_n[5] a_48682_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3300 a_18546_9490# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3301 a_48282_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3302 a_5331_13951# a_5156_14025# a_5510_14013# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3303 a_7373_49007# a_6895_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3304 vcm a_18162_65206# a_26194_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3305 a_22216_30761# a_22186_30485# pmat.en_bit_n[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=1.8668e+12p pd=1.774e+07u as=8.2245e+11p ps=7.66e+06u w=1e+06u l=150000u M=4
X3306 a_2080_31965# a_1643_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3307 VSS a_2407_49289# a_5399_65479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3308 VDD nmat.rowon_n[15] a_36142_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3309 a_20811_34743# a_19689_34789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X331 a_24490_60186# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3310 a_26102_69182# pmat.row_n[13] a_26594_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3311 a_37542_67214# pmat.rowon_n[11] a_37146_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3312 a_30210_63158# a_18546_63200# a_30118_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3313 a_30610_67536# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3314 VDD a_10055_31591# a_14655_53359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X3315 vcm a_18162_15516# a_44266_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3316 a_2375_18708# a_2467_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3317 a_2283_39189# a_2743_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3318 VSS a_35244_32411# a_42307_31756# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X3319 a_24094_8894# pmat.row_n[0] a_24586_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X332 cgen.dlycontrol4_in[0] a_1626_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3320 VDD pmat.rowoff_n[15] a_48190_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3321 VSS a_28189_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3322 a_13966_71631# a_13158_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3323 a_48190_64162# a_18162_64202# a_48282_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3324 VSS pmat.row_n[14] a_30514_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3325 VSS a_2411_43301# a_5256_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3326 VDD a_4167_48463# a_4075_50087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X3327 a_30514_8854# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3328 a_34626_8456# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3329 VDD a_14457_15823# a_14747_7663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X333 a_24490_19898# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3330 VDD a_45251_53047# pmat.col[25] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X3331 a_21174_15516# a_18546_15514# a_21082_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3332 a_3668_6397# a_3551_6202# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3333 VDD a_4461_26133# a_4491_26486# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3334 VDD pmat.rowoff_n[7] a_38150_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3335 a_40969_30287# a_17842_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X3336 a_83276_12015# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X3337 a_10498_19631# a_10151_19637# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X3338 a_8406_11837# a_2021_11043# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3339 a_50198_22950# a_18162_22544# a_50290_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X334 a_8861_24527# a_7415_29397# a_9063_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=7.9e+11p ps=7.58e+06u w=1e+06u l=150000u M=2
X3340 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3341 a_36341_38053# a_34924_37253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X3342 a_49286_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3343 a_21082_55126# VDD a_21574_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3344 a_4859_31274# a_4951_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3345 a_18277_37620# ndecision_finish VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3346 a_43561_47893# a_30111_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X3347 a_42562_61190# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3348 a_19955_30511# a_19605_30511# a_19860_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X3349 a_22097_52815# _1196_.B1 pmat.col_n[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X335 a_23420_39429# a_22357_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X3350 a_39154_66170# a_18162_66210# a_39246_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3351 a_12265_49551# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X3352 a_25190_14512# a_18546_14510# a_25098_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3353 a_25494_71230# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3354 vcm a_18162_11500# a_22178_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3355 a_21269_28585# a_11927_27399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3356 a_39646_11468# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3357 a_32522_72234# VDD a_32126_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3358 a_9441_20189# a_13427_18303# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3359 a_23090_24958# a_18162_24552# a_23182_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X336 a_20217_30511# a_20173_30753# a_20051_30511# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3360 VDD a_40628_39429# a_40532_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X3361 VSS a_20645_42044# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3362 vcm a_18162_10496# a_35230_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3363 VDD a_21815_34191# a_21981_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3364 a_21478_10862# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3365 VDD a_4319_15039# a_3688_17179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3366 VDD _1154_.A a_40415_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3367 a_29206_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3368 a_11885_27247# a_11235_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3369 a_46578_60186# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X337 VSS pmat.row_n[12] a_38546_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3370 a_11397_76457# a_10995_76207# a_11233_76207# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3371 a_46578_19898# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3372 VDD a_1586_18231# a_5087_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3373 VDD a_2163_31741# a_2124_31867# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3374 a_29510_70226# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3375 a_30514_24918# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3376 VDD a_11067_30287# a_21891_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X3377 a_27106_23954# a_18162_23548# a_27198_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3378 a_6432_70767# a_6559_70223# a_6242_70767# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X3379 VDD pmat.rowon_n[9] a_37146_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X338 a_20517_50345# a_19584_52423# a_20445_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3380 vcm a_18162_59182# a_20170_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3381 VSS a_14943_26703# a_17054_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3382 a_51694_71552# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3383 VSS a_40628_39429# a_40591_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X3384 a_19470_62194# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3385 a_47678_61512# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3386 a_21082_72194# a_18162_72234# a_21174_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3387 VSS pmat.row_n[4] a_23486_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3388 a_29937_31055# a_29493_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3389 VSS pmat.row_n[11] a_23486_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X339 VSS a_33423_47695# a_36956_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X3390 a_12531_42583# nmat.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3391 a_20474_16886# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3392 VSS a_39413_40956# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3393 a_51202_61150# a_18162_61190# a_51294_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3394 VDD a_12700_16367# a_12875_16341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3395 a_46130_34319# a_46522_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3396 a_34134_71190# a_18162_71230# a_34226_71190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3397 a_37542_20902# pmat.rowoff_n[12] a_37146_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3398 a_7935_20969# a_6981_21263# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3399 a_33526_15882# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X34 a_35230_22544# a_18546_22542# a_35138_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X340 a_28202_72194# a_18546_72236# a_28110_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3400 VSS a_17113_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3401 VDD nmat.rowon_n[1] a_24094_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3402 vcm a_18162_58178# a_24186_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3403 a_1757_27797# a_1591_27797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3404 a_18103_31421# a_12851_28853# a_17740_31287# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X3405 a_6173_42479# a_6007_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3406 VDD a_30155_42583# a_12116_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X3407 a_3339_70759# a_4075_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3408 a_45471_27497# a_16311_28327# a_45253_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3409 VSS a_45915_29941# a_46395_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X341 VDD a_14533_39631# a_19143_41085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X3410 a_6723_47375# a_6082_46831# a_6641_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.8e+11p pd=2.76e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3411 a_3981_6005# a_3763_6409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X3412 VDD a_29937_31055# a_46797_45993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X3413 VSS a_1769_47919# a_3707_53903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3414 a_36538_68218# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3415 a_28602_72556# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3416 VDD pmat.rowon_n[14] a_32126_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3417 a_25190_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3418 a_22086_11906# a_18162_11500# a_22178_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3419 VDD nmat.rowon_n[5] a_40158_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X342 vcm a_18162_8488# a_31214_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3420 VDD pmat.rowon_n[4] a_28110_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3421 a_49590_67214# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3422 a_30663_50087# a_45107_34863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3423 VSS clk_dig a_12171_18005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3424 VSS a_4987_34293# a_4918_34319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X3425 a_51294_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3426 a_3123_27399# a_3351_27249# a_3297_27275# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3427 a_7824_31433# a_6909_31061# a_7477_31029# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3428 VSS a_4516_21531# a_6747_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3429 a_5718_71311# a_3866_57399# a_5415_71543# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X343 a_36538_71230# pmat.rowon_n[15] a_36142_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3430 a_27340_31055# a_22459_28879# a_27167_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X3431 VSS a_5455_22057# a_5899_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X3432 a_39550_59182# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3433 a_19166_20536# a_18546_20534# a_19074_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3434 a_14460_12265# nmat.rowon_n[7] a_14287_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X3435 a_41162_69182# a_18162_69222# a_41254_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3436 VSS pmat.row_n[1] a_43566_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3437 a_37146_16926# pmat.row_n[8] a_37638_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3438 a_3395_19465# a_2879_19093# a_3300_19453# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X3439 VSS pmat.row_n[11] a_26498_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X344 a_25590_22512# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3440 a_23486_64202# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3441 a_30514_65206# pmat.rowon_n[9] a_30118_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3442 VSS a_7865_59861# a_7799_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3443 VDD _1224_.X a_83677_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3444 a_2369_20541# a_2325_20149# a_2203_20553# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3445 a_6168_32687# a_5253_32687# a_5821_32929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3446 a_44266_66170# a_18546_66212# a_44174_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3447 VDD _1179_.X a_46566_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X3448 a_8996_12559# a_8782_12559# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3449 a_33049_27497# a_24407_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X345 a_35465_32441# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3450 VDD nmat.rowon_n[4] a_44174_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3451 a_23835_40719# a_12228_40693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X3452 a_1757_63701# a_1591_63701# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3453 a_12449_22895# a_12247_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X3454 a_2319_59036# a_2163_58941# a_2464_59165# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X3455 a_22823_32143# a_2007_25597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X3456 a_20474_57174# pmat.rowon_n[1] a_20078_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3457 a_19566_9460# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3458 VSS a_4955_40277# a_4913_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3459 VDD a_12147_24233# a_8583_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X346 a_46274_22544# a_18546_22542# a_46182_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3460 a_1586_50247# a_1683_46295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3461 a_33526_56170# pmat.rowon_n[0] a_33130_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3462 a_18162_13508# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3463 a_27598_15484# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3464 a_21174_7484# a_18546_7482# a_21082_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3465 VDD nmat.rowon_n[10] a_31122_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3466 a_6884_74183# a_7099_74313# a_7026_74358# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X3467 a_48282_65166# a_18546_65208# a_48190_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3468 VSS a_28336_29967# a_43451_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X3469 vcm a_18162_62194# a_45270_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X347 VDD a_2651_29098# a_2422_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3470 a_48682_69544# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3471 a_45178_66170# pmat.row_n[10] a_45670_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3472 VSS a_12557_30485# a_12491_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3473 VDD a_44870_48437# a_45238_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3474 VDD a_9287_77055# a_9274_76751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3475 a_10957_64899# a_10921_64786# a_10885_64899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3476 a_26899_30761# a_24861_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X3477 a_5307_67655# a_7435_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3478 a_20221_40835# a_33765_40229# a_34887_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3479 a_47035_27497# a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X348 VDD pmat.rowon_n[8] a_28110_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3480 a_28110_11906# pmat.row_n[3] a_28602_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3481 a_32256_44869# a_31097_44581# a_32160_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3482 a_22178_62154# a_18546_62196# a_22086_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3483 VDD pmat.rowon_n[13] a_25098_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3484 a_22578_66532# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3485 a_39246_17524# a_18546_17522# a_39154_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3486 a_49194_65166# pmat.row_n[9] a_49686_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3487 a_3484_15101# a_3367_14906# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X3488 a_26460_40517# a_25301_40229# a_26364_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3489 a_50198_60146# pmat.row_n[4] a_50690_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X349 a_2882_74397# a_2124_74299# a_2319_74268# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3490 a_25190_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3491 a_22086_56130# a_18162_56170# a_22178_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3492 VSS a_30111_47911# a_31767_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X3493 VSS a_6051_74183# a_6649_75983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3494 a_36538_21906# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3495 VDD config_2_in[6] a_1591_38127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3496 VSS a_9871_48463# a_6787_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X3497 a_14071_74879# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3498 a_7094_9117# a_6872_8725# a_6412_8725# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.66e+10p pd=1.3e+06u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X3499 a_7413_63151# a_7364_63303# a_7321_63151# VSS sky130_fd_pr__nfet_01v8 ad=3.9e+11p pd=3.8e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X35 VDD a_23455_32447# a_23933_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X350 a_22628_30485# a_20616_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X3500 a_39154_57134# pmat.row_n[1] a_39646_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3501 VSS a_7939_29967# a_4075_31591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X3502 a_43662_55488# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3503 a_30860_48783# a_29076_48695# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=0p ps=0u w=650000u l=150000u M=2
X3504 a_49590_20902# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3505 vcm a_18162_23548# a_44266_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3506 a_38851_28327# a_47499_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3507 a_26594_65528# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3508 a_23090_62154# pmat.row_n[6] a_23582_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3509 VSS pmat.row_n[15] a_47582_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X351 VSS a_5320_30199# a_4951_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3510 a_44266_11500# a_18546_11498# a_44174_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3511 a_13146_12925# a_2835_13077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X3512 a_26102_55126# a_18162_55166# a_26194_55126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3513 a_43720_32143# a_43543_32151# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3514 a_13289_54697# a_12895_53359# a_13091_54447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3515 a_39550_12870# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3516 a_21239_50613# a_21395_50857# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X3517 VSS pmat.row_n[2] a_43566_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3518 nmat.col[18] ANTENNA__1183__B1.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3519 ANTENNA__1183__B1.DIODE a_45405_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X352 VSS a_11261_41245# a_10953_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X3520 VDD a_44444_32233# a_44402_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3521 VSS a_13985_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3522 VDD a_40047_47919# a_33467_46261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3523 VDD pmat.en_C0_n a_20078_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3524 a_26102_14918# pmat.row_n[6] a_26594_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3525 VSS pmat.row_n[12] a_26498_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3526 a_29510_23914# pmat.rowoff_n[15] a_29114_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3527 a_11711_62313# a_10049_60663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X3528 a_21174_23548# a_18546_23546# a_21082_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3529 a_35495_32182# a_35244_32411# a_35036_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X353 a_50594_66210# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3530 VSS nmat.sw a_6469_21813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3531 a_41558_61190# pmat.rowon_n[5] a_41162_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3532 a_30610_12472# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3533 VDD a_5595_65301# a_5553_65577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3534 a_29606_56492# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3535 VSS a_45277_32687# a_47039_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u M=3
X3536 a_34226_22544# a_18546_22542# a_34134_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3537 VSS pmat.row_n[0] a_40554_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3538 VDD nmat.rowon_n[15] a_44174_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3539 VDD a_7072_62037# a_5595_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X354 VDD a_4768_16055# a_4215_15797# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3540 VDD a_9427_50095# a_10233_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X3541 a_19470_15882# pmat.rowoff_n[7] a_19074_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3542 a_38150_7890# VDD a_38642_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3543 a_49286_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3544 a_20474_10862# nmat.rowon_n[13] a_20078_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3545 a_42258_59142# a_18546_59184# a_42166_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3546 VDD a_43548_30287# a_43776_30287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X3547 a_50594_8854# nmat.rowon_n[15] a_50198_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3548 a_38546_18894# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3549 a_43262_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X355 a_47858_53135# ANTENNA__1395__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X3550 pmat.rowoff_n[9] a_14460_61225# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3551 a_45574_60186# pmat.rowon_n[4] a_45178_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3552 vcm a_18162_61190# a_21174_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3553 VSS pmat.row_n[8] a_42562_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3554 a_45574_19898# nmat.rowon_n[4] a_45178_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3555 VSS a_2683_22089# a_9137_27253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3556 VSS a_6564_24527# a_7026_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3557 a_3429_76725# a_3211_77129# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X3558 nmat.col_n[18] a_82787_14709# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3559 a_33033_38567# a_33341_38780# a_33007_38771# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X356 a_2802_51727# a_2676_51843# a_2398_51859# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X3560 a_28506_70226# pmat.rowon_n[14] a_28110_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3561 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3562 VDD a_23063_36885# a_16981_37462# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3563 a_5341_59317# a_4719_58255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3564 a_35729_27497# a_25695_28111# nmat.col[16] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X3565 VDD a_4128_46983# a_6649_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X3566 VSS a_5779_13255# a_5131_13255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3567 VSS a_14287_17455# a_10239_14183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3568 a_50290_68178# a_18546_68220# a_50198_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3569 a_15655_50613# a_12263_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X357 a_5651_66975# a_10703_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3570 a_46274_58138# a_18546_58180# a_46182_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3571 vcm a_18162_55166# a_43262_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3572 VDD a_4025_54965# a_6583_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X3573 a_43170_59142# pmat.row_n[3] a_43662_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3574 a_42166_8894# a_18162_8488# a_42258_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3575 a_5271_35407# a_4601_35727# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3576 a_32522_57174# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3577 VSS a_6087_67655# a_4396_66933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3578 vcm a_18162_67214# a_20170_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3579 a_17187_49783# a_17459_49641# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X358 a_3337_22325# a_3119_22729# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X3580 a_19551_34191# a_19374_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3581 a_6817_21583# a_3351_27249# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X3582 VSS a_11435_58791# a_14441_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3583 vcm a_18162_66210# a_33222_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3584 a_44266_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3585 VSS a_1923_61759# a_2893_59709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3586 VSS a_27913_42333# a_27605_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3587 a_11693_70767# a_11345_70773# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3588 a_33622_19500# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3589 VSS a_7779_22583# a_8031_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 a_29114_72194# VDD a_29606_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3590 VSS comp.adc_inverter_1.in comp.adc_comp_circuit_0.adc_comp_buffer_0.in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3591 a_44806_48783# a_44774_48695# a_44697_48783# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X3592 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3593 a_28202_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3594 VDD a_1644_57141# a_1586_63927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3595 a_20170_10496# a_18546_10494# a_20078_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3596 a_23582_7452# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3597 a_27605_37127# a_26497_36603# a_27619_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3598 VDD nmat.rowon_n[13] a_37146_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3599 a_51598_23914# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_39949_50959# a_39757_50700# pmat.col_n[19] VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X360 a_9427_50095# a_9176_50345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3600 pmat.row_n[3] a_18203_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3601 a_8103_53903# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3602 a_35534_68218# pmat.rowon_n[12] a_35138_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3603 VSS a_2939_45503# a_2389_45859# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3604 vcm a_18162_16520# a_42258_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3605 VDD VDD a_33130_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3606 a_45270_19532# a_18546_19530# a_45178_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3607 VDD a_10595_53361# a_10455_53387# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3608 VDD a_29493_31375# a_29937_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3609 a_17996_35303# a_16837_35515# a_17900_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X361 a_33622_70548# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3610 VDD a_1923_53055# a_1643_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3611 a_14011_14735# a_10515_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X3612 VDD a_2983_48071# a_4985_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X3613 a_10409_53903# a_9871_53903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3614 a_48586_67214# pmat.rowon_n[11] a_48190_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3615 VSS a_11611_50332# a_11542_50461# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X3616 a_3158_13647# a_2400_13763# a_2595_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3617 a_41558_15882# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3618 a_3846_22351# a_2769_22357# a_3684_22729# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3619 a_45222_43567# a_40105_47375# a_44927_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 a_26102_14918# a_18162_14512# a_26194_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3620 VDD a_31535_49525# pmat.col_n[12] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X3621 a_25190_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3622 VSS a_9231_32117# a_9135_60967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3623 a_77882_40202# a_77978_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3624 VDD a_6051_74183# a_6607_75895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3625 a_38546_59182# pmat.rowon_n[3] a_38150_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3626 VDD a_6373_49249# a_6263_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X3627 a_4338_9839# a_1717_13647# a_4169_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X3628 a_22216_30761# a_22628_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3629 VDD nmat.rowon_n[7] a_36142_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X363 VDD a_6720_49007# a_6895_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3630 a_13257_4175# a_10883_3303# nmat.col[3] VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X3631 a_19689_34789# a_17996_35303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X3632 a_9139_68841# a_4583_68021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X3633 a_28336_29967# a_23021_29199# a_28078_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.53e+07u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u M=4
X3634 a_50594_70226# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3635 a_7674_69455# a_4991_69831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3636 vcm a_18162_17524# a_28202_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3637 VSS a_22199_30287# a_42795_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X3638 a_32218_15516# a_18546_15514# a_32126_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3639 a_17403_31599# a_11067_64015# nmat.rowon_n[5] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X364 a_41654_18496# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3640 VDD a_17441_40482# a_16505_40157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X3641 a_13441_70767# a_12809_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3642 a_40554_62194# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3643 a_37146_67174# a_18162_67214# a_37238_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3644 VSS a_10515_15055# a_14195_11791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3645 VSS a_20475_49783# a_22015_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X3646 VSS VDD a_39550_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3647 a_32126_55126# VDD a_32618_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3648 vcm a_18162_7484# a_44266_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3649 a_23486_72234# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X365 a_41558_24918# VSS a_41162_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3650 VSS a_34030_47893# a_13643_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X3651 VDD a_1927_43541# a_1957_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X3652 a_2951_11471# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3653 a_37238_9492# a_18546_9490# a_37146_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3654 vcm a_18162_11500# a_33222_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3655 VDD a_4505_74005# a_4441_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X3656 VDD a_12375_42895# a_12481_42895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3657 a_7212_62607# a_6583_62607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3658 a_41654_24520# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3659 VDD a_13102_71311# a_6451_67655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X366 a_29606_60508# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3660 VDD a_11339_39319# a_12289_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3661 VSS a_26891_28327# a_34948_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3662 VDD a_6564_24527# a_7026_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3663 a_32522_10862# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3664 VDD a_3859_23699# a_2411_16101# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X3665 a_2672_26159# a_1757_26159# a_2325_26401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3666 a_44266_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3667 VSS a_33489_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3668 VDD a_13327_70741# a_13203_70767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3669 a_10226_67503# a_5363_70543# a_10140_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X367 a_30210_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3670 a_27198_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3671 vcm a_18162_9492# a_35230_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3672 a_20016_43781# a_19233_41479# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3673 VDD a_29189_47349# a_29079_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X3674 VDD a_28715_28879# a_28336_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3675 nmat.col_n[12] a_12066_3087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3676 vcm a_18162_70226# a_45270_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3677 VSS config_1_in[10] a_1626_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3678 VDD a_43720_32143# a_46109_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3679 a_45670_23516# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X368 VSS a_10515_75895# a_10853_75119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3680 a_42166_20942# pmat.row_n[12] a_42658_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3681 a_15107_34743# a_15144_35077# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X3682 a_42166_16926# a_18162_16520# a_42258_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3683 a_41162_9898# pmat.row_n[1] a_41654_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3684 a_45270_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3685 cgen.dlycontrol3_in[0] a_1591_44655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3686 VDD pmat.rowon_n[9] a_48190_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3687 a_29159_37607# cgen.dlycontrol2_in[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3688 a_48282_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3689 a_5541_14191# a_5271_14557# a_5451_14557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X369 a_9961_19203# a_3688_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3690 a_51694_9460# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3691 a_32126_72194# a_18162_72234# a_32218_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3692 a_35630_15484# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3693 a_35534_21906# nmat.rowon_n[2] a_35138_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3694 VSS pmat.row_n[4] a_34530_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3695 a_27155_31599# a_23933_32143# a_27066_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X3696 VSS pmat.row_n[11] a_34530_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3697 VSS a_17113_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3698 a_19233_41479# a_18953_43493# a_20075_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3699 a_24490_66210# pmat.rowon_n[10] a_24094_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X37 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u M=325
X370 a_30514_69222# pmat.rowon_n[13] a_30118_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3700 VDD pmat.rowon_n[1] a_38150_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3701 a_22178_70186# a_18546_70228# a_22086_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3702 _1179_.X a_82787_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X3703 a_48682_14480# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3704 a_48586_20902# pmat.rowoff_n[12] a_48190_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3705 VDD pmat.rowoff_n[15] a_22086_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3706 a_13632_47919# pmat.rowon_n[7] a_13329_47893# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3707 a_46182_15922# a_18162_15516# a_46274_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3708 a_32785_47081# a_31675_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3709 VSS a_3052_29967# a_3622_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X371 a_14335_23439# a_9528_20407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3710 a_22086_64162# a_18162_64202# a_22178_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3711 nmat.col_n[19] a_82788_9991# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X3712 a_3211_77129# a_2861_76757# a_3116_77117# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X3713 a_50290_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3714 a_43566_69222# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3715 vcm a_18162_58178# a_35230_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3716 VDD a_39981_37462# a_40532_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X3717 VSS a_12053_27497# a_22792_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3718 VSS ANTENNA__1190__B1.DIODE a_44453_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3719 a_14427_46519# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X372 VDD a_7436_58487# a_7299_58951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3720 a_14347_69831# a_13327_70741# a_14521_69707# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3721 a_38546_12870# pmat.rowoff_n[4] a_38150_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3722 a_36142_11906# pmat.row_n[3] a_36634_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3723 VDD a_9155_17455# a_9557_17705# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3724 a_19074_21946# pmat.row_n[13] a_19566_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3725 a_19074_17930# a_18162_17524# a_19166_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3726 VDD a_46523_39733# a_45019_38645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=8
X3727 a_23090_70186# pmat.row_n[14] a_23582_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3728 VDD nmat.rowon_n[9] a_25098_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3729 a_49194_10902# pmat.row_n[2] a_49686_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X373 a_10195_30186# a_10287_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3730 VDD _1154_.A a_39092_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3731 a_22085_38550# a_22357_39141# a_23479_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3732 a_23182_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3733 a_20078_12910# a_18162_12504# a_20170_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3734 a_43262_61150# a_18546_61192# a_43170_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3735 a_26102_63158# a_18162_63198# a_26194_63158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3736 a_24719_36341# a_12237_36596# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3737 a_47582_68218# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3738 a_37238_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3739 a_36801_42405# a_36345_42567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X374 VDD a_15144_36165# a_15048_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X3740 a_33130_11906# a_18162_11500# a_33222_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3741 VDD a_2847_18303# a_2834_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3742 VDD nmat.rowon_n[5] a_51202_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3743 a_33489_44219# a_32256_44869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X3744 a_4328_6409# a_3247_6037# a_3981_6005# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X3745 a_13349_72405# a_13183_72405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3746 VDD a_24719_37429# a_14773_38306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3747 VDD nmat.rowon_n[10] a_29114_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3748 a_26594_10464# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3749 VSS pmat.row_n[2] a_41558_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X375 a_13459_28111# a_41731_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3750 a_13015_62927# a_13432_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=0p ps=0u w=650000u l=150000u M=2
X3751 a_22195_52521# ANTENNA__1196__A2.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X3752 VSS pmat.row_n[12] a_24490_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3753 a_44174_61150# pmat.row_n[5] a_44666_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3754 a_33501_31599# a_30278_30511# a_33413_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X3755 VDD a_20695_32447# a_18241_31698# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3756 a_15144_36165# a_13985_35877# a_15048_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3757 a_35138_9898# a_18162_9492# a_35230_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3758 vcm a_18162_19532# a_34226_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3759 VDD a_41663_47893# a_13091_52047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X376 a_52398_39208# ctopp comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top VSS sky130_fd_pr__nfet_01v8_lvt ad=4.025e+12p pd=3.144e+07u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u M=4
X3760 vcm a_18162_69222# a_38242_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3761 a_48190_16926# pmat.row_n[8] a_48682_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3762 a_4809_64015# a_4583_68021# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X3763 VSS a_17139_30503# a_24033_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X3764 a_42258_67174# a_18546_67216# a_42166_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3765 a_10239_20291# a_4976_16091# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X3766 a_44573_45173# a_44739_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3767 a_2121_65327# a_1643_65301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3768 VDD a_7355_37013# a_7342_37405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3769 VDD a_7693_22365# a_11241_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X377 a_45284_48169# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.3e+11p pd=5.26e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3770 VDD a_25802_48169# a_25850_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X3771 VSS a_4037_66933# a_2944_67752# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3772 a_39246_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3773 VDD a_3746_58487# a_8051_46607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3774 VDD a_2411_33749# a_4227_34293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3775 a_3267_74817# a_1674_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3776 VSS a_26773_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3777 VSS pmat.row_n[3] a_27502_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3778 VDD pmat.rowon_n[8] a_24094_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3779 a_21574_61512# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X378 a_44570_57174# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3780 a_38242_12504# a_18546_12502# a_38150_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3781 VDD a_18597_31599# a_43543_32151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3782 a_24937_36039# a_24565_34789# a_25687_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3783 a_31518_57174# pmat.rowon_n[1] a_31122_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3784 vcm a_18162_63198# a_43262_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3785 VDD a_6559_70223# a_6521_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3786 a_43170_67174# pmat.row_n[11] a_43662_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3787 a_46182_7890# VDD a_46674_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3788 a_50290_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3789 a_20619_49551# a_20175_49667# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X379 a_23604_44869# a_22541_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X3790 VDD a_17927_47349# pmat.row_n[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3791 a_2882_65693# a_2163_65469# a_2319_65564# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X3792 a_25590_60508# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3793 a_28506_55166# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3794 a_33222_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3795 a_19166_68178# a_18546_68220# a_19074_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3796 a_25260_42693# a_24197_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X3797 a_43566_22910# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3798 a_18546_56172# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3799 a_31701_37462# a_30913_38053# a_31976_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X38 a_24895_35253# a_10873_36341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X380 a_5921_44629# a_4399_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3800 a_50690_17492# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3801 a_50594_23914# pmat.rowoff_n[15] a_50198_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3802 a_37238_18528# a_18546_18526# a_37146_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3803 a_9577_28335# a_5351_19913# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3804 a_30118_24958# VDD a_30610_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3805 a_10873_26409# a_9579_26159# a_10791_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3806 a_20078_57134# a_18162_57174# a_20170_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3807 a_39550_61190# pmat.rowon_n[5] a_39154_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3808 VSS pmat.row_n[9] a_36538_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3809 VSS a_5931_74183# a_5857_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X381 a_8452_77117# a_6292_69831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3810 VSS a_34949_52245# pmat.col_n[14] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3811 a_23707_34165# a_23883_34165# a_23835_34191# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X3812 a_18777_51183# a_18429_51189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3813 a_40554_15882# pmat.rowoff_n[7] a_40158_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3814 VSS a_12449_40693# a_12383_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3815 a_33130_56130# a_18162_56170# a_33222_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3816 a_8481_75663# a_6795_76989# a_7092_74005# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3817 VSS a_22541_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3818 a_47582_21906# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3819 vcm a_18162_24552# a_42258_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X382 a_18546_63200# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X3820 vcm a_18162_66210# a_41254_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3821 a_51202_13914# pmat.row_n[5] a_51694_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3822 vcm a_18162_14512# a_38242_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3823 a_34887_36919# a_34924_37253# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X3824 vcm a_18162_56170# a_37238_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3825 a_3142_9839# a_2021_11043# a_2973_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X3826 a_17842_27497# a_7415_29397# a_18200_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3827 a_34134_23954# pmat.row_n[15] a_34626_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3828 a_34134_19938# a_18162_19532# a_34226_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3829 a_41654_58500# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X383 a_22178_7484# a_18546_7482# a_22086_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3830 a_37542_13874# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3831 a_18546_21538# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3832 a_12311_19783# a_9441_20189# a_12709_19631# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X3833 VSS a_13985_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3834 a_44570_14878# nmat.rowon_n[9] a_44174_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3835 VSS pmat.row_n[3] a_41558_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3836 a_38242_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3837 VSS a_2651_29098# a_2422_29575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3838 a_2012_8573# a_1895_8378# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X3839 VSS config_1_in[9] a_1591_7119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X384 a_27502_67214# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3840 VSS pmat.row_n[0] a_30514_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3841 VSS a_10781_42869# a_10725_43222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3842 a_24094_15922# pmat.row_n[7] a_24586_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3843 VSS pmat.row_n[13] a_24490_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3844 a_27502_24918# VSS a_27106_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3845 VDD a_4031_40455# a_3199_40455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3846 a_35447_50959# a_30663_50087# a_35353_50959# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X3847 a_27598_57496# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3848 a_47211_50069# _1154_.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3849 VDD VSS a_31122_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X385 a_18162_17524# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3850 a_6559_33767# a_7079_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3851 a_32218_23548# a_18546_23546# a_32126_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3852 VSS pmat.row_n[1] a_20474_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3853 a_8456_69135# a_7730_69109# a_4583_68021# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X3854 a_6334_69679# a_6292_69831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3855 VDD a_30663_50087# a_35077_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X3856 a_8809_65149# a_8765_64757# a_8643_65161# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3857 VDD a_3571_13627# a_12815_8213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3858 VDD a_11149_40188# a_11093_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3859 a_4520_60975# a_4041_61225# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X386 VSS pmat.row_n[9] a_31518_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3860 VSS pmat.row_n[4] a_27502_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3861 VSS pmat.row_n[7] a_39550_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3862 a_30514_9858# nmat.rowon_n[14] a_30118_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3863 VDD a_4003_7663# a_4254_7351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3864 a_31518_10862# nmat.rowon_n[13] a_31122_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3865 vcm a_18162_17524# a_36234_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3866 VDD config_2_in[5] a_1591_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3867 VSS a_4257_34319# a_4700_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.1125e+11p ps=1.95e+06u w=650000u l=150000u
X3868 a_40250_15516# a_18546_15514# a_40158_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3869 a_41418_53135# a_18243_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X387 VDD nmat.rowon_n[6] a_31122_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3870 a_21365_27247# a_12061_26703# a_21377_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3871 vcm a_18162_61190# a_32218_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3872 a_2107_39049# a_1591_38677# a_2012_39037# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X3873 a_41254_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3874 a_12543_36950# a_12513_36924# a_12471_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X3875 a_37638_22512# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3876 pmat.sample a_21815_42351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3877 a_6141_44629# a_6732_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3878 VDD pmat.rowoff_n[12] a_41162_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3879 a_23815_50069# a_23971_50228# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X388 VSS a_40415_49551# a_13091_28327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3880 a_45629_35773# a_44763_34293# a_45557_35773# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3881 a_44266_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3882 a_7648_9117# a_6956_8965# a_7040_8725# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3883 VSS a_4259_73807# a_5736_56399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X3884 a_11004_55535# a_10955_55687# a_10913_55535# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X3885 a_1757_8213# a_1591_8213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3886 a_35559_30209# a_6283_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3887 a_37654_47081# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X3888 a_30514_58178# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3889 a_44570_71230# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X389 a_48282_69182# a_18546_69224# a_48190_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3890 VSS a_2840_55509# a_2787_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X3891 vcm a_18162_11500# a_41254_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3892 a_36663_34191# a_36486_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3893 a_2882_52815# a_2163_53057# a_2319_52789# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X3894 VDD a_5351_19913# a_13549_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3895 a_42166_24958# a_18162_24552# a_42258_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3896 a_38150_14918# a_18162_14512# a_38242_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3897 VSS a_3305_27791# a_4443_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3898 a_42258_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3899 a_45270_9492# a_18546_9490# a_45178_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X39 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u M=466
X390 vcm a_18162_66210# a_45270_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3900 a_10391_69653# a_10216_69679# a_10570_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3901 a_29890_47741# a_2263_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X3902 a_48282_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3903 a_45178_60146# a_18162_60186# a_45270_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3904 a_23191_47375# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X3905 VDD a_2219_4943# a_2695_4943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3906 a_26102_56130# pmat.row_n[0] a_26594_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3907 VDD a_7079_40277# a_7066_40669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3908 a_35230_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3909 a_28110_70186# a_18162_70226# a_28202_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X391 a_9485_27247# a_9137_27253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3910 VSS pmat.row_n[15] a_21478_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3911 VDD a_8356_23671# a_8307_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X3912 VDD nmat.rowon_n[12] a_35138_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3913 VDD a_11545_18517# a_11575_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3914 vcm a_18162_22544# a_31214_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3915 a_24941_49257# a_21371_50087# a_24869_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3916 vcm a_18162_12504# a_27198_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3917 a_46182_23954# a_18162_23548# a_46274_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3918 a_46386_33231# a_45829_35407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3919 a_4535_50639# a_2315_44124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X392 a_45670_19500# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3920 a_31214_10496# a_18546_10494# a_31122_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3921 VSS a_26957_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3922 VDD nmat.rowon_n[13] a_48190_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3923 VDD pmat.sample_n a_18162_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X3924 VDD a_2727_58470# a_3801_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X3925 a_46811_33927# a_44444_32233# a_47045_33775# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3926 a_22178_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3927 a_46578_68218# pmat.rowon_n[12] a_46182_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3928 a_14725_26703# a_13479_26935# a_14301_27023# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3929 VSS pmat.row_n[14] a_25494_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X393 a_4241_28335# a_4075_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3930 a_46779_35113# a_43720_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3931 VSS a_40352_41831# a_40315_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X3932 vcm a_18162_71230# a_39246_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3933 a_10515_75895# a_11014_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3934 VDD a_9480_6409# a_9655_6335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3935 a_23182_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3936 a_20078_20942# a_18162_20536# a_20170_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3937 a_19166_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3938 VSS a_17191_48981# pmat.row_n[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X3939 VSS a_1923_69823# a_8441_71677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X394 VSS a_21215_48071# a_24638_49159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X3940 a_39646_63520# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3941 a_11202_55687# a_14163_55295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3942 VDD pmat.rowon_n[5] a_43170_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3943 a_8406_11510# a_2021_11043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3944 VSS pmat.row_n[5] a_28506_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3945 a_31041_42689# a_24833_40719# a_30955_42689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3946 VDD a_5687_71829# a_7044_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3947 a_25494_17890# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3948 a_30210_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3949 a_9023_6031# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X395 VSS pmat.row_n[1] a_21478_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3950 a_32522_18894# nmat.rowon_n[5] a_32126_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3951 VSS a_19689_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X3952 a_17525_36911# a_17459_37143# a_12228_39605# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3953 vcm a_18162_8488# a_24186_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3954 a_20170_58138# a_18546_58180# a_20078_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3955 a_41162_11906# a_18162_11500# a_41254_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3956 a_5711_33053# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3957 a_48190_67174# a_18162_67214# a_48282_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3958 VDD pmat.rowon_n[4] a_47186_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3959 vcm a_18162_59182# a_29206_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X396 a_4340_69455# a_4298_69367# a_4037_69109# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3960 VDD a_2319_56860# a_2250_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X3961 a_41237_28335# a_24747_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3962 a_4032_46983# a_2315_44124# a_4174_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3963 a_33222_57134# a_18546_57176# a_33130_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3964 VSS a_4991_69831# a_11645_68619# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3965 a_34226_8488# a_18546_8486# a_34134_8894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3966 a_30118_58138# pmat.row_n[2] a_30610_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3967 VSS a_19283_49783# a_21970_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X3968 a_29510_16886# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3969 a_45270_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X397 a_6750_70262# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3970 a_27509_44219# a_26552_43781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X3971 VSS pmat.row_n[6] a_33526_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3972 a_30514_11866# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3973 a_27106_10902# a_18162_10496# a_27198_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3974 a_38150_59142# a_18162_59182# a_38242_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3975 a_31976_38341# a_30913_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3976 VSS a_11803_49551# a_12174_50461# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X3977 VDD VDD a_24094_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3978 a_42258_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3979 a_38242_20536# a_18546_20534# a_38150_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X398 a_48586_14878# nmat.rowon_n[9] a_48190_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3980 a_3622_16950# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3981 pmat.rowoff_n[6] a_14458_58799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3982 a_11987_10089# a_11501_10927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3983 a_25180_46831# clk_ena a_25090_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X3984 VSS pmat.row_n[11] a_45574_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3985 a_42562_64202# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3986 a_17308_47491# a_16800_47213# a_17224_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3987 a_40158_21946# pmat.row_n[13] a_40650_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3988 a_6447_35229# a_5823_34863# a_6339_34863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3989 a_8363_56457# a_7847_56085# a_8268_56445# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X399 a_40707_48783# a_40677_48437# a_11711_50959# VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X3990 a_35860_29967# a_35646_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3991 a_13360_14191# a_10239_14183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3992 VDD a_10515_13967# a_14335_16519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3993 a_40158_17930# a_18162_17524# a_40250_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3994 a_5211_57172# a_7067_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3995 a_29187_27791# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X3996 a_7999_31359# a_7824_31433# a_8178_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3997 VDD a_28915_50959# a_46211_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3998 VSS pmat.row_n[3] a_35534_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3999 VDD a_3267_74817# a_3228_74691# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_9741_28585# a_9339_28335# a_9577_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X40 a_22178_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.94708e+14p ps=2.63924e+09u w=800000u l=150000u
X400 VSS pmat.row_n[0] a_34530_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4000 a_28506_63198# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4001 a_2897_21781# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4002 VDD a_7477_31029# a_7367_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4003 VSS a_11113_36483# a_20811_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4004 a_22482_67214# pmat.rowon_n[11] a_22086_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4005 VDD a_13252_18377# a_13427_18303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4006 a_2858_72531# a_3175_72641# a_3133_72765# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X4007 VDD nmat.rowon_n[5] a_49194_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4008 a_46674_15484# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4009 a_43170_12910# pmat.row_n[4] a_43662_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X401 a_28110_15922# pmat.row_n[7] a_28602_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4010 a_46578_21906# nmat.rowon_n[2] a_46182_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4011 a_3016_51727# a_2802_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X4012 VDD nmat.rowon_n[10] a_50198_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4013 VSS a_33341_38780# a_33033_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4014 VDD a_11949_21237# a_11897_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4015 a_20078_65166# a_18162_65206# a_20170_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4016 a_19166_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4017 VDD pmat.rowoff_n[15] a_33130_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4018 a_8013_73493# a_7847_73493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4019 a_36538_13874# nmat.rowon_n[10] a_36142_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X402 a_27605_42693# a_27329_42902# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X4020 VDD a_10423_16055# a_10423_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4021 a_9291_27497# a_4516_21531# a_9219_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4022 a_33130_64162# a_18162_64202# a_33222_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4023 a_23884_40517# a_22725_40229# a_23788_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4024 VSS a_36227_38771# a_36167_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4025 a_44382_40847# a_35312_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X4026 a_4255_66959# a_3983_67503# a_4037_66933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4027 a_19470_65206# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4028 a_19566_17492# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4029 VDD pmat.rowoff_n[7] a_23090_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X403 VSS a_38905_28853# a_40954_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4030 vcm a_18162_64202# a_37238_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4031 a_47186_11906# pmat.row_n[3] a_47678_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4032 VSS a_10589_22351# a_14287_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4033 VSS a_41731_49525# a_34705_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X4034 a_4319_15039# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4035 a_37146_68178# pmat.row_n[12] a_37638_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4036 a_41254_62154# a_18546_62196# a_41162_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4037 VDD pmat.rowon_n[13] a_44174_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4038 a_41654_66532# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4039 VDD a_1586_63927# a_8031_64789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X404 VSS a_16505_40157# a_16197_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X4040 a_23191_47375# a_22567_47381# a_23083_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4041 a_9740_15279# a_8937_15823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X4042 a_34226_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4043 a_11292_38543# a_11041_38772# a_11071_38870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X4044 a_41162_56130# a_18162_56170# a_41254_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4045 VSS a_21279_31599# a_11067_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X4046 a_24094_66170# a_18162_66210# a_24186_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4047 a_29510_57174# pmat.rowon_n[1] a_29114_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4048 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot vcm.sky130_fd_sc_hd__buf_4_0.X VSS VSS sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=4.74e+06u as=0p ps=0u w=500000u l=500000u M=2
X4049 a_11142_64783# a_10707_64783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X405 a_22178_66170# a_18546_66212# a_22086_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4050 a_24586_11468# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4051 VSS a_19948_51959# a_19831_51316# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4052 VDD comp_latch a_7419_14379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4053 a_2683_22089# a_4811_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4054 a_45670_65528# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4055 a_42166_62154# pmat.row_n[6] a_42658_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4056 a_7001_15055# a_3576_17143# a_6917_15055# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4057 VSS a_11067_16359# pmat.rowon_n[5] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4058 VSS ANTENNA__1190__A2.DIODE a_14729_5263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X4059 a_2121_58799# a_1643_58773# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X406 VSS pmat.sample a_18546_64204# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X4060 a_11347_36950# a_11317_36924# a_11275_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X4061 VDD a_33382_46983# a_31152_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X4062 a_31518_60186# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4063 a_31518_19898# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4064 VDD a_22361_41479# a_23420_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4065 a_35630_57496# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4066 VSS a_2046_30184# a_9595_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4067 a_32947_37737# a_33341_37692# a_33007_37683# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X4068 VSS pmat.row_n[12] a_45574_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4069 a_13151_23957# a_12463_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X407 a_32618_13476# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4070 VSS a_29711_47679# a_29645_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X4071 a_40250_23548# a_18546_23546# a_40158_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4072 ANTENNA__1187__B1.DIODE a_46636_36469# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4073 VDD pmat.rowon_n[9] a_22086_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4074 a_48682_56492# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4075 a_36234_13508# a_18546_13506# a_36142_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4076 a_43566_71230# pmat.rowon_n[15] a_43170_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4077 a_11789_69679# a_10864_68565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X4078 VDD nmat.rowon_n[15] a_38150_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4079 a_50198_8894# pmat.row_n[0] a_50690_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X408 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4080 a_28110_63158# pmat.row_n[7] a_28602_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4081 a_32618_61512# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4082 a_49286_12504# a_18546_12502# a_49194_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4083 VSS pmat.row_n[4] a_35534_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4084 a_4383_7093# a_4871_17429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4085 VDD a_14691_27399# a_14471_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.6e+11p ps=7.92e+06u w=1e+06u l=150000u
X4086 a_10497_64489# a_9405_66627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4087 a_10740_68841# a_4991_69831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4088 a_13919_65871# a_13432_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4089 a_26102_8894# pmat.row_n[0] a_26594_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X409 VDD a_3305_17999# a_6579_21583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4090 a_2882_59165# a_2163_58941# a_2319_59036# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X4091 a_22482_20902# pmat.rowoff_n[12] a_22086_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4092 a_5541_71855# a_5687_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X4093 a_19675_51157# a_19831_51316# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X4094 VDD pmat.rowon_n[0] a_25098_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4095 a_33489_43131# a_32072_42919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4096 a_2847_33749# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4097 _1154_.X a_82818_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u M=16
X4098 a_15753_28879# a_15299_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4099 a_47582_70226# pmat.rowon_n[14] a_47186_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X41 vcm a_18162_7484# a_51294_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X410 vcm a_18162_65206# a_49286_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4100 a_32522_8854# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4101 a_6829_26703# a_5320_27023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4102 a_38150_22950# a_18162_22544# a_38242_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4103 a_42258_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4104 VSS a_18953_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X4105 VSS a_1586_8439# a_6375_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4106 VSS a_10515_15055# a_14287_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4107 VDD a_38913_31055# a_40125_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4108 a_6817_29199# a_4516_21531# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X4109 a_37542_62194# pmat.rowon_n[6] a_37146_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X411 a_49194_69182# pmat.row_n[13] a_49686_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4110 a_6830_8751# a_6548_8751# a_6754_8751# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=9.66e+10p ps=1.3e+06u w=420000u l=150000u
X4111 a_9004_47741# a_8453_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4112 a_10129_19203# a_7644_16341# a_10057_19203# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4113 VSS a_12263_50959# a_16403_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4114 VDD VSS a_29114_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4115 VSS a_3351_27249# a_5825_22901# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4116 a_37927_52521# _1184_.A2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4117 a_7523_33775# a_6007_33767# a_7160_33927# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X4118 a_21478_68218# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4119 vcm a_18162_20536# a_27198_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X412 VDD nmat.rowon_n[4] a_22086_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4120 VSS pmat.row_n[9] a_47582_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4121 a_51598_57174# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4122 a_1757_18005# a_1591_18005# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4123 a_51598_15882# pmat.rowoff_n[7] a_51202_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4124 a_6800_44629# a_4128_46983# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X4125 a_34530_67214# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4126 a_44757_37289# a_44811_36469# a_17139_30503# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.44e+12p pd=2.288e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=8
X4127 VSS a_2263_43719# a_23345_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4128 VDD a_31323_29967# a_31399_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4129 VSS a_4068_25615# a_9323_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.225e+11p ps=3.9e+06u w=650000u l=150000u
X413 vcm a_18162_60186# a_50290_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4130 a_29510_10862# nmat.rowon_n[13] a_29114_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4131 a_36142_70186# a_18162_70226# a_36234_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4132 a_1644_53877# a_1591_52815# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4133 vcm a_18162_56170# a_48282_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4134 a_25681_46831# a_25090_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4135 a_24490_59182# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4136 a_48586_13874# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4137 a_22086_16926# pmat.row_n[8] a_22578_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4138 VSS a_4811_22351# a_2683_22089# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X4139 VDD a_44774_40821# a_44382_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X414 a_50198_64162# pmat.row_n[8] a_50690_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4140 VSS a_9919_57863# a_9577_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4141 a_49286_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4142 a_39646_71552# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4143 a_18235_42359# a_17113_42405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4144 VDD a_1781_9308# a_28721_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4145 VDD pmat.rowoff_n[12] a_39154_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4146 a_35138_15922# pmat.row_n[7] a_35630_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4147 a_39154_61150# a_18162_61190# a_39246_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4148 a_20659_49140# a_20267_50345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4149 a_10151_19637# a_8305_20871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X415 VDD nmat.sample a_18546_11498# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X4150 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4151 a_5423_69367# a_5363_70543# a_5597_69473# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4152 a_22522_50247# a_19283_49783# a_22825_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4153 a_40969_30287# a_25575_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4154 a_17113_34789# a_15144_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X4155 a_22138_27907# a_12061_26703# a_22056_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4156 a_28506_16886# nmat.rowon_n[7] a_28110_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4157 VDD a_11793_71311# a_11893_71427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X4158 VSS a_9528_20407# a_12353_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4159 VSS a_7160_33927# a_7067_34293# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X416 VDD _1154_.X a_33049_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X4160 a_7105_27907# a_6917_27907# a_7023_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4161 VSS a_6283_31591# a_26155_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4162 result_out[13] a_1644_72917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4163 VSS a_6917_27907# a_7023_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4164 VSS a_12128_32375# a_11299_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4165 a_2325_40821# a_2107_41225# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X4166 vcm a_18162_67214# a_29206_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4167 a_8627_11837# a_8479_11484# a_8264_11703# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X4168 VDD a_24861_29673# a_26983_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X4169 a_12860_51549# a_12646_51549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X417 VSS a_9103_56383# a_9581_56079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4170 a_33222_65166# a_18546_65208# a_33130_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4171 VSS pmat.row_n[10] a_37542_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4172 vcm a_18162_62194# a_30210_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4173 a_21174_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4174 a_31217_29429# a_19405_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X4175 a_33622_69544# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4176 vcm a_18162_17524# a_47278_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4177 a_30118_66170# pmat.row_n[10] a_30610_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4178 a_2791_57703# a_5692_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4179 a_29206_55126# a_18546_55168# a_29114_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X418 VDD a_3399_24787# a_2952_25045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X4180 a_41558_64202# pmat.rowon_n[8] a_41162_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4181 a_29606_59504# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4182 a_51294_15516# a_18546_15514# a_51202_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4183 a_11793_75663# a_11397_76457# a_6200_70919# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4184 a_8417_24527# a_6173_22895# a_8607_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u M=2
X4185 VSS a_39413_40956# a_39105_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X4186 a_34887_35831# a_34924_36165# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X4187 a_27895_41001# a_26773_40955# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X4188 a_6641_39759# a_5233_40553# a_6127_40516# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4189 a_12067_67279# a_11797_60431# a_11978_67279# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X419 a_6637_69367# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4190 a_11337_28585# a_10814_29111# a_11241_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4191 a_42258_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4192 a_39981_37462# a_39469_38053# a_40591_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4193 a_31085_27221# a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4194 vcm a_18162_7484# a_38242_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4195 a_12960_10749# a_11987_10089# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4196 VSS a_22085_36374# a_22743_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X4197 a_51202_55126# VDD a_51694_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4198 a_42562_72234# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4199 a_5725_24233# a_4068_25615# a_5629_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X42 a_49194_68178# a_18162_68218# a_49286_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X420 VDD a_31701_37462# a_31976_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4200 a_24186_17524# a_18546_17522# a_24094_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4201 a_34134_65166# pmat.row_n[9] a_34626_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4202 a_39246_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4203 a_21478_21906# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4204 VDD a_9521_31353# a_9551_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4205 a_28116_37479# a_26957_37691# a_28020_37479# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4206 a_2715_51969# a_1586_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4207 a_35786_47893# a_30111_47911# a_36956_47919# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X4208 a_51598_10862# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4209 VDD a_79368_40202# a_79181_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X421 a_20995_44265# a_19873_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4210 a_24094_57134# pmat.row_n[1] a_24586_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4211 VSS a_1586_18231# a_2879_19093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4212 a_8643_65161# a_8197_64789# a_8547_65161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4213 a_35534_55166# pmat.en_bit_n[2] a_35138_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4214 a_10991_68591# a_10740_68841# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4215 a_21999_37737# a_22393_37692# a_22059_37683# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X4216 a_34530_20902# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4217 a_3579_15113# a_3063_14741# a_3484_15101# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X4218 VDD a_19332_41959# a_19145_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4219 a_4525_44905# a_2659_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.95e+11p pd=5.19e+06u as=0p ps=0u w=1e+06u l=150000u
X422 VSS pmat.row_n[15] a_40554_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4220 a_4496_28335# a_4379_28548# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X4221 vcm a_18162_13508# a_25190_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4222 a_28202_16520# a_18546_16518# a_28110_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4223 a_46274_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4224 VSS pmat.row_n[15] a_32522_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4225 a_2557_67503# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4226 a_6601_40303# a_6557_40545# a_6435_40303# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X4227 a_28245_44581# a_27789_44743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4228 VDD nmat.rowon_n[12] a_46182_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4229 VDD pmat.rowon_n[12] a_36142_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X423 a_25481_29245# a_22307_27791# a_25409_29245# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4230 a_22823_32143# a_22199_32149# a_22715_32521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4231 a_24490_12870# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4232 vcm.sky130_fd_sc_hd__buf_4_3.A vcm.sky130_fd_sc_hd__buf_4_2.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4233 a_36538_63198# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4234 VDD a_6200_70919# a_11530_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4235 a_20310_28029# a_20695_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4236 vcm a_18162_59182# a_50290_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4237 a_7345_64822# a_6451_67655# a_7131_64822# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4238 a_35167_52521# a_34705_51959# a_34949_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4239 a_49590_62194# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X424 a_5420_62313# a_4985_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4240 a_8264_11703# a_8479_11484# a_8406_11510# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X4241 VDD a_24895_38517# a_24719_38517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4242 a_13547_48169# a_13688_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X4243 a_51202_72194# a_18162_72234# a_51294_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4244 vcm a_18162_72234# a_37238_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4245 a_32305_51335# _1196_.B1 a_32468_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4246 a_50594_16886# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4247 a_22541_43131# a_22085_42902# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4248 VSS a_16552_46805# a_13091_7655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4249 a_41254_70186# a_18546_70228# a_41162_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X425 VSS a_1642_26935# a_1591_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4250 a_40897_48463# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4251 a_13335_65161# a_12889_64789# a_13239_65161# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X4252 a_37238_60146# a_18546_60188# a_37146_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4253 VDD a_46027_44905# a_46797_45993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X4254 a_37638_64524# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4255 VSS a_3331_72373# a_3262_72399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X4256 a_34226_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4257 a_12985_62581# a_12429_62607# a_13656_62927# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X4258 a_23182_7484# a_18546_7482# a_23090_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4259 VDD a_10883_3303# a_13283_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X426 VSS a_39781_40157# a_39473_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X4260 VDD pmat.rowon_n[6] a_41162_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4261 a_41162_64162# a_18162_64202# a_41254_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4262 VDD a_16355_43123# a_16381_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4263 VSS a_17139_30503# a_24765_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4264 a_18397_31599# a_14691_27399# a_18325_31599# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4265 a_46815_37013# a_35244_32411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4266 VDD a_1642_20871# a_1591_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4267 a_38933_30761# a_17842_27497# a_38851_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4268 VSS pmat.sample_n a_18162_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X4269 VSS pmat.row_n[6] a_26498_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X427 a_5085_59663# a_5053_59575# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X4270 a_23486_18894# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4271 a_30514_60186# pmat.rowon_n[4] a_30118_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4272 VSS ANTENNA__1395__A2.DIODE a_83827_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X4273 a_30514_19898# nmat.rowon_n[4] a_30118_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4274 a_6467_29415# a_3576_17143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X4275 VSS a_3305_15823# a_7489_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X4276 a_38927_42359# a_39321_42333# a_38737_41814# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X4277 a_30913_44219# a_29404_44869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4278 VSS a_17619_43439# a_17725_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4279 a_42166_70186# pmat.row_n[14] a_42658_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X428 a_25143_28585# a_22307_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X4280 VDD nmat.rowon_n[9] a_44174_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4281 a_36617_37691# a_36161_37462# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4282 VSS a_1769_13103# a_1775_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4283 a_27198_71190# a_18546_71232# a_27106_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4284 a_38150_60146# pmat.row_n[4] a_38642_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4285 VDD VSS a_27106_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4286 a_4165_70767# a_2791_57703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4287 a_3480_17143# a_3305_15823# a_3622_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X4288 a_44741_36201# a_35244_32411# a_44647_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X4289 a_31214_58138# a_18546_58180# a_31122_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X429 VSS a_20164_27791# a_20616_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4290 a_47035_36495# a_45019_38645# a_46636_36469# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.195e+12p pd=1.039e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4291 VSS a_3175_72641# a_3136_72515# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4292 a_1769_47919# a_1769_13103# a_1937_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u w=1e+06u l=150000u M=2
X4293 a_7865_59861# a_4075_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4294 VSS a_19176_35279# a_19282_35279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4295 a_20570_9460# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4296 a_2325_23413# a_2107_23817# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X4297 a_4984_41935# a_3983_41941# a_4912_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4298 VSS a_1923_53055# a_1881_55357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4299 a_36234_21540# a_18546_21538# a_36142_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X43 a_24773_49257# a_22499_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X430 a_40158_56130# pmat.row_n[0] a_40650_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4300 a_45670_10464# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4301 a_28110_71190# pmat.row_n[15] a_28602_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4302 a_11737_53359# a_4128_64391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X4303 VDD nmat.rowon_n[14] a_30118_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4304 a_28602_20504# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4305 VSS pmat.row_n[12] a_43566_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4306 a_40554_65206# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4307 a_2757_58621# a_2727_58470# a_2685_58621# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4308 a_28202_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4309 a_49286_20536# a_18546_20534# a_49194_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X431 a_27890_32143# a_24374_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4310 a_30863_46831# a_31105_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=0p ps=0u w=650000u l=150000u M=2
X4311 VDD a_33467_46261# a_37791_46811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4312 VSS a_4031_32852# a_3091_33402# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4313 a_33775_29111# a_31263_28309# a_33925_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4314 a_44888_33205# a_30663_50087# a_45545_33551# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X4315 a_27619_36649# a_27605_37127# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4316 a_20315_29098# a_13643_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4317 VDD nmat.rowon_n[13] a_22086_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4318 VSS a_10515_15055# a_14471_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4319 a_36142_63158# pmat.row_n[7] a_36634_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X432 a_24602_48169# a_19541_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X4320 a_20474_68218# pmat.rowon_n[12] a_20078_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4321 a_40650_61512# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4322 VSS pmat.row_n[3] a_46578_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4323 a_43566_56170# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4324 a_29114_12910# a_18162_12504# a_29206_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4325 VDD a_2879_57487# a_3431_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4326 a_10299_51433# a_10245_51335# a_10205_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X4327 a_30210_19532# a_18546_19530# a_30118_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4328 a_5156_28335# a_4075_28335# a_4809_28577# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4329 VDD a_3776_77129# a_3951_77055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X433 a_26194_65166# a_18546_65208# a_26102_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4330 a_50594_57174# pmat.rowon_n[1] a_50198_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4331 a_6634_26133# a_4516_21531# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4332 a_44666_16488# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4333 a_18546_70228# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4334 VSS a_19689_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X4335 VSS pmat.row_n[13] a_29510_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4336 VDD a_36380_34191# a_36486_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4337 VDD a_14589_35286# a_13653_35516# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X4338 a_33526_67214# pmat.rowon_n[11] a_33130_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4339 a_18162_24552# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X434 vcm a_18162_62194# a_23182_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4340 a_34797_51727# a_34942_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X4341 VSS a_11133_34427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X4342 a_6173_42479# a_6007_42479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4343 a_4951_76983# a_4429_76751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4344 a_11163_22057# a_7693_22365# a_11067_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4345 a_23486_59182# pmat.rowon_n[3] a_23090_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4346 a_47582_55166# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4347 VDD nmat.rowon_n[7] a_21082_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4348 a_38242_68178# a_18546_68220# a_38150_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4349 a_35161_49007# a_24867_53135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X435 a_12447_16143# a_20879_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X4350 VSS nmat.sample_n a_18162_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X4351 a_28110_18934# a_18162_18528# a_28202_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4352 a_1643_69653# a_1846_69931# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4353 vcm a_18162_64202# a_48282_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4354 VDD cgen.dlycontrol2_in[3] a_29159_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4355 a_48190_68178# pmat.row_n[12] a_48682_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4356 VSS a_2867_43541# a_2411_43301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4357 a_22086_67174# a_18162_67214# a_22178_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4358 a_27502_58178# pmat.rowon_n[2] a_27106_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4359 a_17141_51843# a_16800_47213# a_17046_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X436 a_26594_69544# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4360 VSS VDD a_24490_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4361 VDD ANTENNA__1197__A.DIODE a_22097_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4362 a_2927_22134# a_1781_9308# a_2468_21959# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4363 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top vcm.sky130_fd_sc_hd__buf_4_3.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=3.16e+06u as=4.35e+11p ps=4.74e+06u w=500000u l=500000u M=2
X4364 a_8723_67191# a_8819_67197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X4365 a_22977_32509# a_22933_32117# a_22811_32521# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X4366 a_44174_8894# a_18162_8488# a_44266_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4367 a_36234_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4368 a_35138_66170# a_18162_66210# a_35230_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4369 a_2215_15823# a_1591_15829# a_2107_16201# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X437 a_23090_66170# pmat.row_n[10] a_23582_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4370 a_2012_28157# a_1895_27962# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4371 cgen.dlycontrol2_in[3] a_1591_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4372 a_46225_47695# a_45112_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X4373 a_10045_59887# a_10195_59861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4374 a_39550_23914# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4375 a_19689_44581# a_17996_44007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X4376 a_17397_48463# a_17049_48579# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X4377 a_8031_61839# a_2215_47375# a_7937_61839# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X4378 VSS pmat.row_n[13] a_43566_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4379 a_25590_7452# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X438 VSS pmat.sample_n a_18162_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X4380 a_21478_7850# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4381 vcm a_18162_70226# a_30210_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4382 a_46674_57496# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4383 a_46968_45743# a_47290_45717# a_47236_45743# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X4384 a_29206_63158# a_18546_63200# a_29114_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4385 VSS a_9395_27791# a_10609_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4386 a_41558_72234# VDD a_41162_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4387 VDD a_22343_50613# pmat.row_n[14] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4388 a_30610_23516# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4389 a_29606_67536# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X439 a_37739_43177# a_36345_42567# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X4390 a_30210_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4391 a_51294_23548# a_18546_23546# a_51202_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4392 a_45489_30511# a_30663_50087# a_45405_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X4393 VSS VDD a_31518_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4394 VDD pmat.rowon_n[9] a_33130_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4395 a_9166_51843# a_8385_51727# a_9084_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4396 a_47278_13508# a_18546_13506# a_47186_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4397 a_29114_57134# a_18162_57174# a_29206_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4398 a_33222_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4399 VDD ANTENNA__1187__B1.DIODE pmat.col_n[11] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X44 a_12815_26409# a_10223_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X440 VSS nmat.sample_n a_18162_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X4400 a_20570_15484# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4401 a_49590_15882# pmat.rowoff_n[7] a_49194_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4402 VSS pmat.row_n[4] a_46578_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4403 a_20474_21906# nmat.rowon_n[2] a_20078_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4404 a_50594_10862# nmat.rowon_n[13] a_50198_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4405 VDD pmat.rowon_n[1] a_23090_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4406 VSS pmat.row_n[14] a_29510_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4407 VSS a_45325_38127# a_47357_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4408 a_38546_70226# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4409 a_33622_14480# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X441 VDD pmat.rowon_n[11] a_30118_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4410 a_33526_20902# pmat.rowoff_n[12] a_33130_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4411 a_31122_15922# a_18162_15516# a_31214_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4412 VSS cgen.dlycontrol1_in[2] a_26767_34967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4413 a_7435_32182# a_4128_64391# a_6976_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4414 vcm a_18162_61190# a_51294_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4415 a_7385_51701# a_7167_52105# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X4416 a_25743_49783# a_25839_49783# a_26141_49871# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X4417 VSS a_6823_58951# a_3938_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4418 VSS a_24270_49783# a_23971_50228# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4419 VDD a_46339_31029# _1194_.B1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=8
X442 a_44266_15516# a_18546_15514# a_44174_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4420 a_23486_12870# pmat.rowoff_n[4] a_23090_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4421 a_35534_63198# pmat.rowon_n[7] a_35138_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4422 VSS vcm.sky130_fd_sc_hd__inv_1_4.Y a_79718_39826# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4423 a_21082_11906# pmat.row_n[3] a_21574_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4424 VSS a_6895_48981# a_6829_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4425 vcm a_18162_21540# a_25190_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4426 a_28202_24552# a_18546_24550# a_28110_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4427 a_34828_37253# a_33765_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4428 a_43170_71190# a_18162_71230# a_43262_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4429 a_48586_62194# pmat.rowon_n[6] a_48190_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X443 VSS a_1923_69823# a_9913_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4430 a_34134_10902# pmat.row_n[2] a_34626_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4431 a_33130_7890# a_18162_7484# a_33222_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4432 VSS a_3305_27791# a_5070_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X4433 VDD a_12447_16143# a_16679_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X4434 vcm a_18162_7484# a_46274_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4435 a_5779_71285# a_8283_71829# a_8231_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X4436 a_32522_68218# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4437 a_5633_71631# a_2879_57487# a_5415_71543# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4438 a_8820_6397# a_8703_6202# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4439 VDD pmat.rowon_n[2] a_27106_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X444 a_26102_59142# a_18162_59182# a_26194_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4440 a_11307_14191# a_10957_14191# a_11212_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4441 a_5136_19783# a_5351_19913# a_5278_19958# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X4442 a_39246_9492# a_18546_9490# a_39154_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4443 a_2439_13889# a_3571_13627# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4444 VSS a_11547_48061# a_11508_48187# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4445 vcm a_18162_67214# a_50290_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4446 a_27502_11866# nmat.rowon_n[12] a_27106_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4447 a_14749_48285# a_14486_47919# a_14336_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4448 VDD a_24867_53135# a_43261_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X4449 a_9217_24233# a_8831_24501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X445 ctopn nmat.sw ctopn VDD sky130_fd_pr__pfet_01v8 ad=2.7075e+12p pd=2.185e+07u as=0p ps=0u w=1.9e+06u l=220000u M=2
X4450 a_27753_35073# a_27687_34967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4451 a_31695_43439# a_31518_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4452 a_47186_70186# a_18162_70226# a_47278_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4453 VSS pmat.row_n[15] a_40554_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4454 a_39550_64202# pmat.rowon_n[8] a_39154_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4455 VDD a_6343_32661# a_6330_33053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4456 a_35534_59182# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4457 vcm a_18162_12504# a_46274_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4458 VSS a_31263_32117# a_7939_31591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4459 a_37638_72556# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X446 a_37680_42919# a_36617_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4460 a_12960_10749# a_11987_10089# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X4461 VDD nmat.rowon_n[2] a_37146_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4462 a_3859_22655# a_3684_22729# a_4038_22717# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4463 VDD pmat.rowon_n[14] a_41162_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4464 vcm a_18162_69222# a_23182_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4465 a_33130_16926# pmat.row_n[8] a_33622_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4466 a_50290_10496# a_18546_10494# a_50198_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4467 a_1895_36666# a_1899_35051# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4468 a_37146_62154# a_18162_62194# a_37238_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4469 a_20078_19938# pmat.row_n[11] a_20570_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X447 a_30210_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4470 a_32035_43177# a_30913_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4471 a_45277_32687# a_44923_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4472 a_41254_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4473 a_23849_51727# _1194_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4474 VSS a_46968_45743# a_30111_47911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4475 a_24186_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4476 VSS _1194_.A2 a_83276_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4477 VSS a_12263_50959# a_18521_46837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4478 VDD a_2747_74549# a_1823_76181# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4479 a_23182_12504# a_18546_12502# a_23090_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X448 VDD a_8744_71689# a_8919_71615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4480 vcm a_18162_68218# a_27198_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4481 a_38242_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4482 a_4579_47919# a_4071_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4483 a_9414_12559# a_8695_12801# a_8851_12533# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X4484 VSS a_4865_8181# a_2972_9991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4485 a_38770_50755# a_25879_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4486 VSS a_1781_9308# a_1725_9334# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4487 vcm a_18162_18528# a_45270_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4488 a_2012_39037# a_1895_38842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4489 a_27198_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X449 a_2407_49289# a_4627_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4490 a_79085_39738# a_79181_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4491 a_44570_17890# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4492 a_2672_26159# a_1591_26159# a_2325_26401# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4493 a_35230_71190# a_18546_71232# a_35138_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4494 VDD a_27603_34191# a_30771_39425# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4495 VDD a_4259_31375# a_7033_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4496 VSS a_13561_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X4497 VDD a_11883_62063# a_11895_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X4498 a_28202_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4499 a_25098_21946# a_18162_21540# a_25190_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X45 VDD a_39505_38780# a_39111_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X450 VSS a_33281_49551# a_10883_3303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X4500 VDD pmat.rowon_n[7] a_35138_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4501 a_22178_18528# a_18546_18526# a_22086_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4502 VDD a_11057_35836# a_11001_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X4503 a_4921_32441# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4504 a_18235_41271# a_17113_41317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4505 a_39246_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4506 a_25224_27247# a_9411_2215# a_24921_27221# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4507 a_14528_68841# a_13327_70741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4508 a_24490_61190# pmat.rowon_n[5] a_24094_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4509 VSS pmat.row_n[9] a_21478_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 VSS a_1644_58229# result_out[3] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4510 a_21891_47081# pmat.rowon_n[7] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4511 VSS a_13605_71017# a_13633_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4512 a_2107_23817# a_1757_23445# a_2012_23805# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4513 a_46182_10902# a_18162_10496# a_46274_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4514 a_36142_71190# pmat.row_n[15] a_36634_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4515 VDD a_6283_31591# a_37471_32149# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4516 a_9133_6005# a_8915_6409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X4517 a_32522_21906# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4518 a_29114_20942# a_18162_20536# a_29206_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4519 VDD pmat.rowon_n[6] a_39154_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X452 a_4071_47919# a_3978_48071# a_3983_47919# VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=6.565e+11p ps=5.92e+06u w=650000u l=150000u
X4520 a_11505_25321# a_9075_28023# a_11251_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u M=2
X4521 a_11541_69929# a_11487_69653# a_8439_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4522 a_35138_57134# pmat.row_n[1] a_35630_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4523 vcm a_18162_14512# a_23182_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4524 a_44266_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4525 VDD a_2407_49289# a_7345_64822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4526 a_46578_55166# VSS a_46182_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4527 a_25190_59142# a_18546_59184# a_25098_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4528 vcm a_18162_56170# a_22178_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4529 VDD nmat.rowon_n[7] pmat.rowon_n[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u M=4
X453 a_35630_8456# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4530 VSS a_41427_31599# a_41427_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X4531 VDD nmat.rowon_n[7] a_14460_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X4532 a_4135_19391# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4533 a_22482_13874# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4534 VSS pmat.row_n[8] a_25494_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4535 a_22787_34709# a_11041_38772# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4536 a_10995_76207# a_11023_76359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4537 a_12543_37277# a_12289_36950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4538 VDD a_42462_48071# a_42138_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4539 a_23182_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X454 a_11985_20969# a_11711_20725# a_11903_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4540 a_9701_32509# a_9666_32275# a_9231_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4541 a_8360_7485# a_8243_7290# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4542 a_40951_31599# a_40678_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4543 a_35534_12870# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4544 a_47582_63198# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4545 VDD a_35465_32441# a_35495_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4546 VSS a_30857_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X4547 VDD a_9103_73791# a_9090_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4548 vcm a_18162_55166# a_26194_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4549 a_10291_77269# a_10494_77547# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X455 a_17323_27791# a_7026_24527# a_17573_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=7.9e+11p ps=7.58e+06u w=1e+06u l=150000u M=2
X4550 a_26102_59142# pmat.row_n[3] a_26594_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4551 VDD a_23700_38567# a_23604_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4552 a_8655_64783# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X4553 vcm a_18162_72234# a_48282_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4554 a_14829_29423# a_13655_26703# a_14471_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=8.6e+11p ps=7.72e+06u w=1e+06u l=150000u
X4555 a_45178_22950# pmat.row_n[14] a_45670_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4556 a_38242_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4557 a_24959_31055# a_22628_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=9.65e+11p pd=7.93e+06u as=0p ps=0u w=1e+06u l=150000u
X4558 VSS pmat.row_n[7] a_24490_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4559 VSS a_6927_30503# a_12371_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X456 a_44174_55126# VDD a_44666_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4560 vcm a_18162_17524# a_21174_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4561 a_38642_17492# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4562 a_38546_23914# pmat.rowoff_n[15] a_38150_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4563 VSS a_4123_76181# a_2999_76922# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4564 a_37542_9858# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4565 a_10677_35303# a_10985_35516# a_10651_35507# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4566 a_36142_18934# a_18162_18528# a_36234_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4567 a_14499_26703# a_13145_26935# a_14391_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X4568 VDD pmat.rowoff_n[7] a_42166_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4569 a_39359_49172# a_38793_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X457 VSS a_9319_50639# a_9184_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4570 a_45019_38645# a_46523_39733# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=8
X4571 a_20776_51959# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4572 a_14645_28381# a_10589_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4573 VSS a_28613_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X4574 a_22578_22512# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4575 VSS a_3879_42997# a_2263_43719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4576 a_49194_21946# pmat.row_n[13] a_49686_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4577 VSS pmat.row_n[1] a_47582_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4578 a_49194_17930# a_18162_17524# a_49286_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4579 a_4809_28577# a_4591_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X458 a_12250_4175# a_9411_2215# a_12164_4175# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4580 a_50198_12910# a_18162_12504# a_50290_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4581 a_13347_64783# a_3339_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X4582 a_7436_58487# a_4843_54826# a_7578_58294# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X4583 a_16837_40955# a_16171_40157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4584 a_17882_31094# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X4585 VSS a_12292_44869# a_12255_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X4586 VSS a_2319_56860# a_2250_56989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X4587 a_39154_13914# pmat.row_n[5] a_39646_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4588 VDD a_41731_49525# a_43267_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X4589 a_38876_39655# a_37813_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 a_30514_22910# nmat.rowon_n[1] a_30118_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4590 a_45282_32143# a_44571_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4591 a_4885_58255# a_4719_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4592 a_43662_11468# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4593 VSS pmat.row_n[8] a_28506_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4594 nmat.col[30] _1196_.B1 a_83656_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4595 VDD a_24895_37429# a_24719_37429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4596 a_26594_21508# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4597 a_30371_37737# a_30765_37692# a_30431_37683# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X4598 a_10769_77295# a_10291_77269# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4599 a_23090_14918# a_18162_14512# a_23182_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X46 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u M=466
X460 a_27106_65166# pmat.row_n[9] a_27598_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4600 VDD a_2199_13887# a_7176_8751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4601 a_26194_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4602 a_47278_21540# a_18546_21538# a_47186_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4603 a_38379_52047# a_13091_28327# pmat.col_n[18] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4604 a_29114_65166# a_18162_65206# a_29206_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4605 a_22743_41001# a_21621_40955# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X4606 a_21087_43177# a_19965_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4607 VSS a_9135_60967# a_12155_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4608 a_33222_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4609 a_30118_60146# a_18162_60186# a_30210_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X461 a_25129_31751# a_24861_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4610 VDD a_14335_16519# a_14195_7351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4611 a_6837_42255# a_6369_39465# a_6554_43255# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4612 a_20170_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4613 VDD nmat.rowon_n[7] a_19074_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4614 a_29053_31375# a_24374_29941# a_29243_31375# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X4615 VDD nmat.rowon_n[12] a_20078_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4616 a_47731_36103# a_40837_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4617 a_31122_23954# a_18162_23548# a_31214_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4618 a_29606_12472# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4619 VSS a_24565_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X462 VSS a_11927_27399# a_16965_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.49925e+12p ps=2.199e+07u w=650000u l=150000u M=4
X4620 a_18272_39429# a_17113_39141# a_18235_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X4621 VDD a_4432_42313# a_4608_41909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4622 a_27106_13914# a_18162_13508# a_27198_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4623 VDD nmat.rowon_n[13] a_33130_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4624 a_14809_53359# a_11067_64015# a_14737_53359# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4625 a_47186_63158# pmat.row_n[7] a_47678_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4626 a_30913_43131# a_30140_43781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4627 a_33765_40229# a_33084_40743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X4628 a_31518_68218# pmat.rowon_n[12] a_31122_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4629 a_51694_61512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X463 VDD a_45112_47607# a_45113_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X4630 VSS a_18241_31698# a_34243_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4631 a_42658_19500# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4632 VDD a_11389_40443# a_24753_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4633 a_4128_64391# a_6343_32661# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4634 vcm a_18162_71230# a_24186_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4635 VSS a_13653_35516# a_13345_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X4636 a_32522_9858# nmat.rowon_n[14] a_32126_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4637 a_11041_26409# a_4068_25615# a_10969_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4638 VDD pmat.rowon_n[0] a_44174_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4639 VSS a_1586_33927# a_1591_38677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X464 nmat.sample a_20711_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X4640 a_15107_35831# a_13985_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4641 a_9135_22057# a_8507_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X4642 a_22097_48579# a_21215_48071# a_22015_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4643 VSS a_24937_41479# a_25319_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X4644 VSS a_2149_45717# a_5857_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4645 VDD pmat.rowon_n[10] a_27106_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4646 a_24586_63520# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4647 VDD a_11823_74895# a_12225_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4648 a_5399_65479# a_4583_68021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4649 a_2107_50095# a_1757_50095# a_2012_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X465 a_48282_14512# a_18546_14510# a_48190_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4650 a_3622_17277# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4651 a_20848_39429# a_19689_39141# a_20752_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4652 a_43262_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4653 a_18546_67216# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X4654 a_49286_68178# a_18546_68220# a_49194_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4655 VDD config_2_in[9] a_2603_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4656 a_9037_73865# a_7847_73493# a_8928_73865# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X4657 VDD _1154_.A a_82787_54421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4658 a_44420_45895# a_44628_45717# a_44562_45743# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4659 a_4403_51701# a_1957_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X466 VSS pmat.row_n[0] a_41558_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4660 a_20078_68178# a_18162_68218# a_20170_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4661 a_39550_72234# VDD a_39154_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4662 vcm a_18162_20536# a_46274_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4663 a_50198_57134# a_18162_57174# a_50290_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4664 VDD a_22628_30485# a_23352_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X4665 a_28602_62516# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4666 a_27313_51701# ANTENNA__1197__B.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X4667 a_33130_67174# a_18162_67214# a_33222_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4668 a_12693_38543# a_12267_38870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4669 VDD pmat.rowon_n[4] a_32126_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X467 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4670 a_13173_68597# a_10991_68591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4671 a_2493_11477# a_2327_11477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4672 a_2012_20541# a_1895_20346# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4673 VDD a_43315_48437# a_45370_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=2
X4674 a_47278_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4675 VDD ANTENNA__1395__A1.DIODE a_39307_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X4676 VSS a_34816_34191# a_34922_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4677 a_5921_11791# a_5579_12394# a_5602_11791# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=4.7125e+11p ps=4.05e+06u w=650000u l=150000u
X4678 vcm a_18162_22544# a_19166_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4679 a_23090_59142# a_18162_59182# a_23182_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X468 VDD nmat.rowon_n[15] a_45178_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4680 a_11067_49871# a_30833_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4681 a_23182_20536# a_18546_20534# a_23090_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4682 a_37542_24918# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4683 a_43566_17890# nmat.rowon_n[6] a_43170_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4684 a_41162_16926# pmat.row_n[8] a_41654_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4685 a_19166_10496# a_18546_10494# a_19074_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4686 a_11883_66191# a_11797_60431# a_9643_66389# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4687 a_26498_69222# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4688 VSS pmat.row_n[11] a_30514_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4689 a_30571_50959# a_41427_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X469 VSS a_20645_42044# a_20337_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X4690 VDD a_5651_66975# a_12265_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4691 VDD clk_ena a_21891_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4692 a_29493_31375# a_29635_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X4693 a_12245_21807# a_11897_21813# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X4694 a_24847_37455# a_11497_38543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X4695 a_44266_56130# a_18546_56172# a_44174_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4696 a_22201_48169# a_18823_50247# a_22105_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4697 a_5687_71829# a_12131_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4698 a_27106_58138# a_18162_58178# a_27198_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4699 VSS pmat.row_n[3] a_20474_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 VSS a_54790_39936# comp.adc_nor_latch_0.NOR_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.65e+11p ps=1.66e+06u w=500000u l=150000u M=2
X470 a_48586_71230# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4700 a_13593_8573# a_13549_8181# a_13427_8585# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4701 nmat.rowoff_n[2] a_14839_9295# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4702 a_47582_16886# nmat.rowon_n[7] a_47186_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4703 VSS pmat.row_n[5] a_44570_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4704 a_12665_69135# a_12152_66415# a_12581_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4705 VDD pmat.rowon_n[15] a_35138_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4706 a_27106_17930# pmat.row_n[9] a_27598_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4707 VSS pmat.row_n[15] a_27502_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4708 cgen.start_conv_in a_1591_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4709 a_9195_60039# a_9135_60967# a_9369_59915# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X471 vcm a_18162_11500# a_45270_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4710 a_31614_15484# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4711 a_31518_21906# nmat.rowon_n[2] a_31122_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4712 a_30999_48071# a_32827_46805# a_32785_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4713 a_35230_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4714 a_48282_55126# a_18546_55168# a_48190_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4715 a_18162_71230# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4716 a_48682_59504# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4717 VSS a_43533_30761# a_46108_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4718 a_21478_55166# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4719 VDD a_6283_31591# a_38391_48469# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X472 a_82833_27497# ANTENNA__1197__A.DIODE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4720 a_21478_13874# nmat.rowon_n[10] a_21082_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4721 a_11347_37277# a_11093_36950# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4722 vcm a_18162_8488# a_50290_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4723 VDD pmat.rowon_n[14] a_39154_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4724 a_4162_64561# a_4128_64391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.58e+11p pd=2.36e+06u as=0p ps=0u w=420000u l=150000u
X4725 a_46578_63198# pmat.rowon_n[7] a_46182_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4726 a_25190_67174# a_18546_67216# a_25098_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4727 vcm a_18162_64202# a_22178_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4728 a_32126_11906# pmat.row_n[3] a_32618_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4729 VDD ANTENNA__1195__A1.DIODE a_83741_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X473 a_44533_33749# a_45908_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X4730 a_11797_65871# a_10921_64786# a_9643_66389# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X4731 a_22086_68178# pmat.row_n[12] a_22578_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4732 vcm a_18162_8488# a_26194_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4733 a_3746_58487# a_4043_33535# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X4734 a_12196_44869# a_12292_44869# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X4735 a_43262_17524# a_18546_17522# a_43170_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4736 a_4161_64239# a_4128_64391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.323e+11p pd=1.47e+06u as=0p ps=0u w=420000u l=150000u
X4737 VDD pmat.rowon_n[3] a_25098_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4738 a_40677_48437# a_40949_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X4739 a_42769_50069# a_28131_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X474 a_7645_17455# a_4976_16091# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X4740 a_18546_7482# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X4741 vcm.sky130_fd_sc_hd__buf_4_2.X a_77428_38962# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X4742 VDD a_1586_33927# a_6007_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4743 a_31504_46831# a_31105_46805# a_30833_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4744 a_35799_35831# a_36193_35805# a_11297_36091# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X4745 result_out[14] a_1644_74549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4746 VSS a_7644_16341# a_11711_20725# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4747 vcm a_18162_63198# a_26194_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4748 a_6564_24527# a_4523_21276# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4749 a_31976_38567# a_32072_38567# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X475 a_12568_35077# a_11409_34789# a_12531_34743# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X4750 a_26102_67174# pmat.row_n[11] a_26594_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4751 a_37542_65206# pmat.rowon_n[9] a_37146_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4752 VDD a_16926_46261# a_13091_18535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4753 a_30610_65528# pmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4754 vcm a_18162_13508# a_44266_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4755 VDD a_25221_46519# a_25189_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X4756 VSS a_9227_20291# a_7779_22583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4757 VSS pmat.row_n[15] a_51598_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4758 VDD a_11803_49551# a_12174_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4759 VSS a_22393_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X476 a_44570_10862# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4760 VDD nmat.rowon_n[2] a_48190_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4761 VSS a_21365_27247# a_22015_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4762 a_3111_53333# a_1591_52815# a_3054_54223# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X4763 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4764 a_20570_57496# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4765 a_26498_22910# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4766 a_48190_62154# a_18162_62194# a_48282_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4767 VSS pmat.row_n[12] a_30514_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4768 VDD a_13779_43123# a_13805_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4769 a_3297_27275# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X477 a_44647_35520# a_43776_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X4770 a_33622_56492# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4771 a_21174_13508# a_18546_13506# a_21082_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4772 a_5081_52521# a_2315_44124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4773 VDD nmat.rowon_n[10] a_38150_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4774 VSS a_9092_31287# a_7619_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4775 a_34226_12504# a_18546_12502# a_34134_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4776 VSS pmat.row_n[4] a_20474_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4777 a_50198_20942# a_18162_20536# a_50290_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4778 a_31307_49871# _1183_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X4779 vcm a_18162_19532# a_43262_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X478 a_51598_8854# nmat.rowon_n[15] a_51202_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4780 VDD a_11547_48061# a_11508_48187# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4781 a_47947_52047# a_24867_53135# pmat.col[28] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4782 a_49286_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4783 VDD a_3571_13627# a_11711_12565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4784 a_11435_58791# a_15655_50613# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X4785 a_9414_63695# a_8695_63937# a_8851_63669# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X4786 a_44697_48783# a_45370_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4787 VSS pmat.row_n[6] a_45574_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4788 a_42562_18894# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4789 VSS a_19865_46983# a_19678_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X479 a_36178_48169# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X4790 a_1757_23445# a_1591_23445# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4791 a_4441_74281# a_4409_74183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4792 VSS VDD a_28506_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4793 a_32522_70226# pmat.rowon_n[14] a_32126_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4794 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4795 VDD a_78165_39738# a_77978_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4796 VSS a_4461_46805# a_4395_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4797 a_23090_22950# a_18162_22544# a_23182_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4798 a_13655_26703# a_13437_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X4799 a_46274_71190# a_18546_71232# a_46182_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X48 vcm a_18162_55166# a_31214_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X480 a_2007_25597# a_2879_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X4800 a_3795_70223# a_3710_70455# a_3577_70197# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4801 VSS a_20411_51157# a_14653_53458# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X4802 a_27887_41271# a_27947_41245# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X4803 a_50290_58138# a_18546_58180# a_50198_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4804 a_12592_18365# a_11145_17999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X4805 VDD pmat.rowon_n[7] a_46182_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4806 a_22482_62194# pmat.rowon_n[6] a_22086_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4807 a_47011_31029# a_47685_30517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X4808 VDD a_25575_31055# a_40967_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X4809 VDD a_3305_17999# a_5705_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 a_21574_55488# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4810 VDD nmat.rowon_n[14] a_19793_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4811 VDD a_20616_27791# a_26899_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X4812 VDD a_6975_76823# a_8481_75663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4813 VSS pmat.row_n[9] a_32522_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4814 VDD a_24833_34191# a_25647_34343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4815 VSS a_9463_50877# a_10319_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X4816 a_47186_71190# pmat.row_n[15] a_47678_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4817 a_42258_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4818 VSS ANTENNA__1190__B1.DIODE a_45469_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X4819 a_7808_61493# a_1823_66941# a_8031_61839# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X482 VDD a_6559_6031# a_7206_5853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4820 vcm a_18162_57174# a_20170_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4821 a_12155_27791# a_11711_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4822 a_19470_60186# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4823 a_18162_58178# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X4824 a_19470_19898# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4825 a_36175_50345# a_30663_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.95e+11p pd=5.19e+06u as=0p ps=0u w=1e+06u l=150000u
X4826 a_21082_70186# a_18162_70226# a_21174_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4827 a_19488_52423# a_16800_47213# a_19719_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4828 a_20474_14878# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4829 vcm a_18162_56170# a_33222_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X483 a_27502_20902# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4830 a_33526_13874# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4831 a_9480_6409# a_8399_6037# a_9133_6005# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X4832 a_20879_47893# a_21215_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X4833 a_6649_75983# a_6607_75895# a_5497_73719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X4834 a_46130_34639# a_29937_31055# a_46130_34319# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4835 a_12905_17973# a_12687_18377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X4836 a_34226_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4837 a_24586_71552# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4838 VSS a_5341_59317# a_4956_59317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4839 VDD pmat.rowoff_n[12] a_24094_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X484 VSS a_36265_48981# a_22499_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8675e+11p ps=3.79e+06u w=650000u l=150000u M=2
X4840 VSS a_16355_43123# a_16295_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4841 VDD a_13140_50247# a_13091_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4842 VSS a_13227_42333# a_13167_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4843 a_15324_44007# a_14261_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4844 a_24094_61150# a_18162_61190# a_24186_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4845 a_4025_54965# a_6559_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X4846 VDD a_23821_35279# a_28591_36519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4847 VSS pmat.row_n[13] a_48586_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4848 a_45574_66210# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4849 VSS pmat.row_n[0] a_36538_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X485 VDD a_9839_47679# a_9826_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4850 a_14289_5737# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X4851 a_11497_38543# a_11071_38870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4852 VSS a_1644_71285# result_out[12] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4853 a_43170_23954# pmat.row_n[15] a_43662_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4854 a_43170_19938# a_18162_19532# a_43262_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4855 a_39469_38053# a_37776_37479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4856 a_4675_54599# a_4025_54965# a_4909_54447# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4857 a_4351_55527# a_4927_50613# a_4535_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4858 a_46578_8854# nmat.rowon_n[15] a_46182_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4859 a_50198_65166# a_18162_65206# a_50290_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X486 vcm a_18162_23548# a_22178_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4860 VDD a_5012_10927# a_3576_17143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X4861 a_28602_70548# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4862 a_49286_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4863 VDD ANTENNA__1197__A.DIODE a_42987_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X4864 a_42562_59182# pmat.rowon_n[3] a_42166_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4865 a_36634_18496# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4866 a_36538_24918# nmat.en_bit_n[0] a_36142_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4867 a_18546_24550# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4868 a_25190_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4869 a_1923_69823# a_2387_70483# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X487 vcm.sky130_fd_sc_hd__buf_4_0.A vcm.sky130_fd_sc_hd__dlymetal6s6s_1_3.X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4870 a_17740_31287# a_12851_28853# a_17882_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X4871 VDD nmat.rowon_n[7] a_40158_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4872 a_25494_69222# pmat.rowon_n[13] a_25098_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4873 VSS pmat.row_n[10] a_22482_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4874 a_49590_65206# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4875 a_34530_8854# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4876 vcm a_18162_17524# a_32218_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4877 a_19873_44219# a_19417_43990# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X4878 a_49686_17492# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4879 VSS a_5043_37191# a_4127_37013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X488 VSS pmat.row_n[5] a_42562_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4880 a_3824_57487# a_3770_57399# a_3704_57487# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X4881 a_47186_18934# a_18162_18528# a_47278_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4882 VDD ANTENNA__1190__A1.DIODE a_27623_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X4883 a_10423_16055# a_10167_16950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4884 VSS a_47223_38671# _1192_.B1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4885 a_39550_57174# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4886 VSS a_18660_47607# a_18083_47593# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4887 a_41162_67174# a_18162_67214# a_41254_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4888 VSS VDD a_43566_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4889 a_33109_52245# a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X489 a_31122_12910# pmat.row_n[4] a_31614_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4890 a_38150_8894# a_18162_8488# a_38242_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4891 a_12813_31029# a_12595_31433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X4892 VDD a_39647_47679# a_39634_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4893 a_29510_68218# pmat.rowon_n[12] a_29114_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4894 VSS pmat.row_n[9] a_26498_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4895 VSS a_24407_31375# a_39392_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4896 VDD a_30699_29397# a_31154_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4897 VDD nmat.rowon_n[6] a_26102_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4898 a_37463_39095# a_36341_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4899 a_24186_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X49 a_44266_9492# a_18546_9490# a_44174_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X490 a_39246_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4900 VDD a_4383_7093# a_6641_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4901 a_13335_31359# a_13160_31433# a_13514_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4902 a_44266_64162# a_18546_64204# a_44174_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4903 nmat.col[17] a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X4904 a_44666_68540# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4905 a_26479_32117# a_27443_32143# a_27976_32463# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X4906 a_2203_28169# a_1757_27797# a_2107_28169# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X4907 a_20474_55166# pmat.en_C0_n a_20078_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4908 a_3521_33205# a_3303_33609# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X4909 a_14340_19783# a_9963_13967# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=0p ps=0u w=650000u l=150000u
X491 VDD a_11435_58791# a_13645_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X4910 a_35885_36165# a_11297_36091# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4911 a_19566_7452# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4912 VDD a_22063_46519# a_21837_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4913 VSS pmat.row_n[0] a_29510_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4914 a_7263_52105# a_6817_51733# a_7167_52105# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X4915 a_31214_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4916 a_18162_11500# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X4917 a_4897_58575# a_1823_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X4918 a_27598_13476# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4919 a_41475_31751# a_39939_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X492 a_27502_8854# nmat.rowon_n[15] a_27106_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4920 a_33084_40743# a_31925_40955# a_32988_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4921 VDD nmat.rowon_n[12] a_31122_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4922 a_48282_63158# a_18546_63200# a_48190_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4923 vcm a_18162_60186# a_45270_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4924 VDD a_23883_34165# a_23707_34165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4925 VDD pmat.rowon_n[12] a_21082_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4926 VSS a_4491_53511# a_4123_52789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4927 VDD a_2672_41225# a_2847_41151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4928 a_48682_67536# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4929 a_45178_64162# pmat.row_n[8] a_45670_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X493 a_36161_37462# a_36341_38053# a_37463_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4930 a_21478_63198# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4931 a_34883_28111# ANTENNA__1195__A1.DIODE nmat.col[14] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4932 a_20911_51843# a_18823_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4933 a_31393_49551# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.55e+11p pd=2.51e+06u as=0p ps=0u w=1e+06u l=150000u
X4934 a_25794_49007# a_25839_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4935 VSS pmat.row_n[15] a_35534_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4936 a_34530_62194# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4937 VDD a_54790_39936# comp.adc_nor_latch_0.NOR_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u M=2
X4938 vcm a_18162_72234# a_22178_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4939 VDD pmat.rowon_n[1] a_42166_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X494 a_22178_11500# a_18546_11498# a_22086_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4940 VSS pmat.row_n[14] a_48586_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4941 a_4752_42301# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4942 vcm a_18162_22544# a_40250_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4943 VDD a_26552_36165# a_26456_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4944 a_22178_60146# a_18546_60188# a_22086_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4945 vcm a_18162_71230# a_35230_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4946 VDD pmat.rowon_n[11] a_25098_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4947 a_39246_15516# a_18546_15514# a_39154_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4948 a_22578_64524# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4949 VSS a_3305_17999# a_5825_22901# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X495 a_6641_25731# a_4068_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4950 a_14562_46403# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X4951 a_9020_7497# a_7939_7125# a_8673_7093# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4952 a_25190_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4953 a_23182_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4954 a_13909_66959# a_13432_62581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=0p ps=0u w=1e+06u l=150000u
X4955 VDD a_5731_58951# a_5731_58799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4956 VDD a_1923_69823# a_1643_74005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4957 a_1643_52789# a_1846_52947# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4958 a_28848_42919# a_27785_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4959 a_42562_12870# pmat.rowoff_n[4] a_42166_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X496 vcm a_18162_22544# a_35230_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4960 VDD a_25802_48169# a_26242_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X4961 a_2847_36799# a_2672_36873# a_3026_36861# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4962 VSS ANTENNA__1197__B.DIODE a_46934_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4963 a_39154_55126# VDD a_39646_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4964 VDD a_2325_26401# a_2215_26525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4965 a_25494_22910# nmat.rowon_n[1] a_25098_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4966 VDD a_4579_47919# a_6829_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4967 VDD a_12693_38543# a_17525_36911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4968 vcm a_18162_21540# a_44266_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4969 a_11058_62063# a_10286_60405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X497 a_11023_76359# a_10699_75119# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4970 a_23090_60146# pmat.row_n[4] a_23582_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4971 a_51598_68218# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4972 a_30860_48783# a_28901_48437# a_30189_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4973 a_35353_50959# a_30571_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4974 a_39550_10862# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4975 VSS a_2563_34837# a_2509_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4976 VDD a_7407_17455# a_7809_17705# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4977 a_24861_29673# a_8583_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4978 a_5253_11177# a_5223_11079# a_4998_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.05e+11p ps=7.61e+06u w=1e+06u l=150000u M=2
X4979 a_27001_30511# a_23933_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X498 VSS a_1957_43567# a_14209_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4980 VDD a_5351_19913# a_6836_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4981 a_29510_21906# nmat.rowon_n[2] a_29114_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4982 VSS pmat.row_n[5] a_37542_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4983 a_26102_12910# pmat.row_n[4] a_26594_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4984 VDD a_5687_71829# a_11990_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4985 a_21174_21540# a_18546_21538# a_21082_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4986 VDD a_16911_52423# a_14287_70543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X4987 a_30610_10464# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4988 a_41558_18894# nmat.rowon_n[5] a_41162_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4989 VDD a_23541_52245# pmat.col[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X499 a_1846_31851# a_2163_31741# a_2121_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X4990 VSS _1187_.A2 a_29825_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4991 a_32740_50095# a_28915_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.8675e+11p pd=3.79e+06u as=0p ps=0u w=650000u l=150000u
X4992 a_34226_20536# a_18546_20534# a_34134_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4993 a_22015_48579# a_18823_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4994 a_48586_24918# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4995 a_5749_57685# a_4351_55527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4996 VSS a_2199_13887# a_4853_14013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4997 VSS a_3305_15823# a_6469_21813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4998 a_12479_41046# a_12228_40693# a_12020_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4999 a_19470_13874# nmat.rowon_n[10] a_19074_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5 VSS a_4421_67477# a_4036_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X50 a_25209_44581# a_23700_44869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X500 VDD comp.adc_inverter_1.out comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=3.32e+06u w=500000u l=150000u M=4
X5000 vcm a_18162_69222# a_42258_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5001 VSS a_13459_28111# a_47947_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X5002 vcm a_18162_59182# a_38242_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5003 a_37146_9898# pmat.row_n[1] a_37638_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5004 a_4697_74005# a_4225_71311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X5005 a_42258_57134# a_18546_57176# a_42166_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5006 VSS a_24407_31375# a_30100_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5007 VSS a_5779_71285# a_6772_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X5008 a_39154_72194# a_18162_72234# a_39246_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5009 a_5545_17027# a_5271_17271# a_5463_17027# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X501 a_26411_42717# a_11041_40948# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X5010 a_20848_38341# a_19689_38053# a_20752_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5011 a_38546_16886# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5012 a_9460_10615# a_9668_10651# a_9602_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5013 a_43262_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5014 a_35099_34191# a_34922_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5015 VSS pmat.row_n[6] a_42562_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5016 a_47678_9460# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5017 a_21082_63158# pmat.row_n[7] a_21574_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5018 a_3208_33597# a_3091_33402# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5019 a_12217_46831# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X502 a_24490_13874# nmat.rowon_n[10] a_24094_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5020 VSS pmat.row_n[3] a_31518_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5021 a_25098_18934# pmat.row_n[10] a_25590_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5022 result_out[6] a_1644_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X5023 VDD a_4921_32441# a_4951_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5024 vcm a_18162_68218# a_46274_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5025 VDD pmat.rowon_n[15] a_46182_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5026 a_23479_35831# a_22357_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5027 a_7536_48579# a_6787_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5028 VSS a_2387_70483# a_1923_69823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X5029 a_25190_7484# a_18546_7482# a_25098_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X503 VSS pmat.row_n[2] a_21478_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5030 a_19948_51959# a_12263_50959# a_20179_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5031 a_46274_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5032 VSS a_4075_50087# a_4627_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X5033 VSS a_12851_28853# a_17702_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X5034 vcm a_18162_9492# a_30210_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5035 a_29206_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5036 a_11781_46831# a_11071_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5037 a_9681_8527# a_2648_29397# a_9463_8439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5038 VSS a_1591_31599# a_1683_46295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5039 a_32522_55166# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X504 VDD a_13091_7655# a_13551_8751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5040 a_23182_68178# a_18546_68220# a_23090_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5041 vcm a_18162_65206# a_20170_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5042 a_44174_21946# a_18162_21540# a_44266_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5043 a_28079_39913# a_28116_39655# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X5044 a_20078_69182# pmat.row_n[13] a_20570_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5045 a_19166_58138# a_18546_58180# a_19074_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5046 a_41254_18528# a_18546_18526# a_41162_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5047 VDD a_8491_47911# a_12613_57141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5048 vcm a_18162_64202# a_33222_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5049 a_29114_19938# pmat.row_n[11] a_29606_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X505 vcm a_18162_59182# a_43262_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5050 a_33130_68178# pmat.row_n[12] a_33622_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5051 a_6574_5853# a_6448_5755# a_6170_5739# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5052 VSS pmat.row_n[9] a_40554_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5053 a_1757_38677# a_1591_38677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5054 a_82789_26677# ANTENNA__1395__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X5055 a_79368_39738# vcm.sky130_fd_sc_hd__nand2_1_1.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5056 a_6311_42692# a_6554_43255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5057 a_2464_59165# a_2250_59165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5058 a_51598_21906# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5059 a_21174_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X506 a_5865_18543# a_5821_18785# a_5699_18543# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5060 a_17808_34215# a_16745_34427# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5061 vcm a_18162_14512# a_42258_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5062 VSS a_25287_32117# a_6007_33767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5063 vcm a_18162_56170# a_41254_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5064 VDD a_9323_28879# a_9785_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X5065 ANTENNA__1395__A2.DIODE a_37820_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5066 VDD nmat.rowon_n[14] a_32126_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5067 a_30913_38053# a_29220_37253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X5068 a_48586_65206# pmat.rowon_n[9] a_48190_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5069 VSS a_2319_31836# a_2250_31965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X507 a_14696_26409# a_8861_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5070 a_41558_13874# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5071 a_4843_54826# a_8749_57141# a_8697_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5072 a_24490_23914# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5073 a_4492_32375# a_3746_58487# a_4634_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5074 a_9103_56383# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5075 a_2847_26133# a_2672_26159# a_3026_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5076 a_14553_29423# a_14465_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5077 a_25190_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5078 a_36234_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5079 VDD a_6283_31591# a_38391_47381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X508 VSS a_30913_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5080 a_38546_57174# pmat.rowon_n[1] a_38150_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5081 a_31614_57496# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5082 VSS a_2648_29397# a_2592_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5083 VDD a_45805_32661# a_45119_32661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5084 a_6522_32687# a_2411_33749# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5085 vcm a_18162_15516# a_28202_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5086 VSS a_2244_20871# cgen.dlycontrol4_in[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5087 a_18769_36965# a_18180_38341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X5088 VSS a_12429_62607# a_13015_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5089 a_32218_13508# a_18546_13506# a_32126_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X509 a_44174_72194# a_18162_72234# a_44266_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5090 a_10569_64489# a_5363_70543# a_10497_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5091 a_14163_55295# a_13988_55369# a_14342_55357# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5092 nmat.rowon_n[10] a_14458_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5093 a_2629_55357# a_2250_54991# a_2557_55357# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5094 VSS pmat.row_n[4] a_31518_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5095 a_32988_40743# a_31925_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5096 VSS pmat.row_n[7] a_43566_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5097 a_40554_60186# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5098 VSS a_6821_18543# a_10239_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5099 a_40554_19898# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X51 a_1674_68047# a_1644_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X510 a_49590_63198# pmat.rowon_n[7] a_49194_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5100 a_23486_70226# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5101 a_30118_9898# a_18162_9492# a_30210_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5102 a_4227_34293# a_4514_34451# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5103 a_48586_7850# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5104 a_17424_27497# a_7026_24527# a_17047_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.175e+12p ps=1.035e+07u w=1e+06u l=150000u M=4
X5105 a_44266_72194# a_18546_72236# a_44174_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5106 a_37146_24958# VDD a_37638_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5107 a_2334_49334# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X5108 VSS a_35036_32375# a_31263_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5109 VDD a_32072_42919# a_31976_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X511 VSS pmat.row_n[4] a_46578_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5110 a_41654_22512# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5111 a_31393_31055# a_31263_28309# a_30527_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X5112 a_20474_63198# pmat.rowon_n[7] a_20078_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5113 a_6061_38377# a_5687_38279# a_5989_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5114 VSS a_4535_56623# a_2879_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5115 a_19439_28585# a_7840_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X5116 VDD nmat.rowon_n[6] a_34134_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5117 a_33526_62194# pmat.rowon_n[6] a_33130_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5118 VSS a_5065_63669# a_4680_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X5119 VDD a_44449_31029# a_37291_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u M=2
X512 VSS pmat.row_n[11] a_46578_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5120 a_9741_28585# a_4339_27804# a_9669_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5121 a_45178_72194# VDD a_45670_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5122 a_46182_8894# a_18162_8488# a_46274_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5123 a_45670_21508# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5124 a_45270_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5125 a_42166_14918# a_18162_14512# a_42258_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5126 a_41162_7890# VDD a_41654_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5127 ANTENNA__1197__B.DIODE a_40837_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=8
X5128 a_35534_7850# VDD a_35138_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5129 a_51694_7452# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X513 a_43566_16886# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5130 a_14471_20175# a_9963_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5131 a_32126_70186# a_18162_70226# a_32218_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5132 a_35630_13476# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5133 a_78165_40202# a_78261_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5134 a_24490_64202# pmat.rowon_n[8] a_24094_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5135 VDD VSS a_38150_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5136 a_4445_64239# a_4162_64561# a_4032_64391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5137 vcm a_18162_12504# a_31214_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5138 a_18162_19532# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X5139 a_39246_23548# a_18546_23546# a_39154_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X514 a_43170_8894# a_18162_8488# a_43262_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5140 VDD a_45345_31029# a_34204_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5141 a_22578_72556# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5142 a_48682_12472# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5143 VDD nmat.rowon_n[2] a_22086_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5144 a_2953_33237# a_2787_33237# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5145 a_36723_27247# _1154_.X nmat.col[17] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X5146 a_46182_13914# a_18162_13508# a_46274_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5147 a_14734_4175# a_9411_2215# a_14648_4175# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X5148 a_25190_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5149 a_22086_62154# a_18162_62194# a_22178_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X515 a_41443_28879# a_41192_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5150 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5151 a_11793_67503# a_10975_67503# a_11019_71543# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5152 a_43566_67214# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5153 VSS _1224_.X a_83238_4175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2675e+12p ps=1.3e+07u w=650000u l=150000u M=4
X5154 VSS a_11057_35836# a_11001_35862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5155 a_50594_68218# pmat.rowon_n[12] a_50198_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5156 VSS a_1717_13647# a_8257_10422# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5157 VSS a_27579_34967# a_14600_37607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5158 VSS VDD a_33526_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5159 a_35138_61150# a_18162_61190# a_35230_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X516 a_45747_51433# a_17139_30503# a_45529_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5160 a_38546_10862# nmat.rowon_n[13] a_38150_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5161 a_26498_9858# nmat.rowon_n[14] a_26102_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5162 VDD a_19817_37692# a_19423_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5163 a_7177_27907# a_7140_27805# a_7105_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5164 a_3063_55535# a_2727_58470# a_2969_55535# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X5165 a_19074_15922# a_18162_15516# a_19166_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5166 VDD pmat.rowoff_n[4] a_25098_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5167 VDD a_14839_54599# a_14839_54447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5168 a_14427_46519# a_14699_46377# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5169 a_8287_71311# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X517 a_27339_30511# a_24861_29673# a_27001_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X5170 vcm a_18162_61190# a_39246_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5171 a_23182_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5172 a_14899_31599# a_14453_31599# a_14803_31599# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X5173 a_43662_63520# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5174 a_42617_47081# a_35186_47375# a_42191_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X5175 a_2897_21781# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5176 a_12175_27221# a_12075_24847# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5177 a_37238_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5178 vcm a_18162_18528# a_30210_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5179 a_47678_18496# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X518 VSS pmat.row_n[14] a_29510_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5180 VSS a_2407_49289# a_7352_65149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5181 a_2407_49289# a_4627_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X5182 VSS a_17625_42902# a_16689_43132# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X5183 VDD a_6787_47607# a_11793_75663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5184 a_12700_16367# a_11785_16367# a_12353_16609# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5185 VDD nmat.rowon_n[7] a_51202_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5186 VSS nmat.sample_n a_18162_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X5187 VDD a_5715_16911# a_5731_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5188 a_5893_46831# a_4985_51433# a_5455_46831# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=5.07e+11p ps=5.46e+06u w=650000u l=150000u
X5189 a_10921_64786# a_14289_66421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X519 a_11977_66415# a_11883_62063# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X5190 a_20170_71190# a_18546_71232# a_20078_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5191 a_37542_58178# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5192 VDD nmat.rowon_n[12] a_29114_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5193 VSS a_18243_28327# a_41784_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5194 VDD pmat.rowon_n[12] a_19074_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5195 a_4613_19087# a_4135_19391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5196 a_2334_49007# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5197 a_10190_60663# a_11007_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5198 a_5797_24233# a_4337_22351# a_5725_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5199 VDD pmat.rowon_n[7] a_20078_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X52 a_31122_59142# pmat.row_n[3] a_31614_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X520 a_2833_14013# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5200 VSS a_1957_43567# a_11541_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5201 a_45832_51183# ANTENNA__1197__A.DIODE a_45529_51157# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X5202 a_35138_7890# a_18162_7484# a_35230_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5203 vcm a_18162_67214# a_38242_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5204 a_20874_32509# a_1858_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5205 VSS a_7079_40277# a_7013_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X5206 a_42258_65166# a_18546_65208# a_42166_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5207 a_42658_69544# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5208 nmat.col[26] _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X5209 pmat.rowon_n[1] a_14839_54447# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X521 VSS a_11435_58791# a_14257_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5210 a_28020_38567# a_26957_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X5211 a_38012_52271# a_11067_27239# a_37709_52245# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X5212 pmat.rowon_n[7] a_21647_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5213 a_12902_26159# a_10223_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5214 VSS a_1644_76181# result_out[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5215 VDD a_17902_43439# a_21815_42351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5216 a_31122_10902# a_18162_10496# a_31214_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5217 a_21082_71190# pmat.row_n[15] a_21574_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5218 a_42166_59142# a_18162_59182# a_42258_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5219 a_25098_69182# a_18162_69222# a_25190_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X522 VDD pmat.rowoff_n[15] a_34134_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5220 VSS pmat.row_n[1] a_27502_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5221 VDD pmat.rowon_n[6] a_24094_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5222 a_38242_10496# a_18546_10494# a_38150_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5223 a_31518_55166# VSS a_31122_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5224 a_18162_9492# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X5225 a_13268_2223# ANTENNA__1196__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5226 VSS a_77245_39738# a_77058_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5227 VSS a_2411_33749# a_6601_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5228 a_6263_49373# a_5639_49007# a_6155_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5229 nmat.col_n[13] a_14734_4175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X523 a_30118_18934# pmat.row_n[10] a_30610_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5230 a_32371_47349# a_11067_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X5231 a_43170_65166# pmat.row_n[9] a_43662_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5232 a_12513_39100# a_13555_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5233 a_13549_21263# a_4523_21276# a_13467_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5234 a_26456_41605# a_26317_40726# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X5235 VSS a_11389_40443# a_24667_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X5236 VDD nmat.rowon_n[4] a_28110_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5237 a_13146_58621# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5238 a_10791_26409# a_4068_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5239 a_46182_58138# a_18162_58178# a_46274_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X524 a_19074_8894# a_18162_8488# a_19166_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5240 a_32522_63198# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5241 a_29114_68178# a_18162_68218# a_29206_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5242 a_9183_72007# a_9375_72007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5243 VSS a_5081_53135# a_6978_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5244 a_7066_40669# a_5989_40303# a_6904_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5245 a_46182_17930# pmat.row_n[9] a_46674_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5246 VSS pmat.row_n[15] a_46578_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5247 a_6037_59887# a_6175_60039# a_6128_59887# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=0p ps=0u w=650000u l=150000u
X5248 a_43566_20902# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5249 a_50690_15484# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X525 a_27198_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5250 a_50594_21906# nmat.rowon_n[2] a_50198_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5251 VDD a_2467_46506# a_1987_45370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5252 a_40250_9492# a_18546_9490# a_40158_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5253 vcm a_18162_72234# a_33222_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5254 a_37238_16520# a_18546_16518# a_37146_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5255 a_30118_22950# pmat.row_n[14] a_30610_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5256 VSS a_6343_32661# a_6277_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5257 VSS a_14917_23983# a_18397_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5258 a_23182_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5259 a_20078_55126# a_18162_55166# a_20170_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X526 a_37927_52521# a_24591_28327# a_37709_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5260 a_7275_51727# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X5261 VSS pmat.row_n[7] a_36538_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5262 a_39550_18894# nmat.rowon_n[5] a_39154_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5263 a_10045_59887# a_8491_47911# a_8841_60405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5264 a_40554_13874# nmat.rowon_n[10] a_40158_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5265 VDD a_4337_22351# a_5271_23447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5266 a_40317_52271# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X5267 a_23582_17492# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5268 a_23486_23914# pmat.rowoff_n[15] a_23090_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5269 a_20078_14918# pmat.row_n[6] a_20570_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X527 vcm a_18162_68218# a_51294_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5270 a_21082_18934# a_18162_18528# a_21174_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5271 a_51202_11906# pmat.row_n[3] a_51694_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5272 VSS a_1899_35051# a_6127_40516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5273 vcm a_18162_64202# a_41254_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5274 a_25393_35877# a_24937_36039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X5275 a_41162_68178# pmat.row_n[12] a_41654_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5276 VSS a_41443_28879# a_41964_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5277 VSS a_9135_60967# a_9976_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X5278 a_37146_58138# pmat.row_n[2] a_37638_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5279 a_41481_52245# _1187_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X528 VDD nmat.rowon_n[1] a_47186_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5280 a_34134_21946# pmat.row_n[13] a_34626_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5281 VDD a_39045_37692# a_38651_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5282 a_34134_17930# a_18162_17524# a_34226_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5283 a_29079_47375# a_28455_47381# a_28971_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5284 VDD pmat.rowon_n[3] a_44174_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5285 a_7281_51183# a_4259_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X5286 VDD a_2099_25236# a_1895_26372# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5287 a_37542_11866# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5288 a_12040_16367# a_11881_16911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5289 VDD a_14427_46519# a_14379_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X529 vcm a_18162_58178# a_47278_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5290 a_8215_69929# a_8439_69653# a_7730_69109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5291 a_26498_56170# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5292 a_46921_30511# a_30571_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5293 a_33331_31599# a_29163_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.646e+11p pd=2.94e+06u as=0p ps=0u w=420000u l=150000u
X5294 a_25671_40719# cgen.dlycontrol3_in[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5295 a_2467_46506# a_2559_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5296 a_24094_13914# pmat.row_n[5] a_24586_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5297 VDD a_2651_8916# a_1949_9308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5298 a_11041_39860# a_11347_40214# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5299 a_27598_55488# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X53 vcm.sky130_fd_sc_hd__buf_4_0.X a_77428_40594# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X530 a_5038_28853# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X5300 vcm a_18162_23548# a_28202_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5301 a_32218_21540# a_18546_21538# a_32126_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5302 a_2163_74173# a_1674_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5303 a_10781_42364# a_30955_42689# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5304 VDD nmat.en_bit_n[0] a_36142_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5305 a_17285_32117# pmat.rowon_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5306 a_4680_63669# a_2407_49289# a_4903_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X5307 VSS a_4991_69831# a_8538_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5308 VSS pmat.row_n[2] a_27502_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5309 a_50198_19938# pmat.row_n[11] a_50690_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X531 a_82736_4943# _1154_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.955e+12p pd=1.791e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X5310 a_9050_14774# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X5311 VSS a_17021_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5312 a_45279_50959# a_24867_53135# pmat.col[26] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5313 vcm a_18162_15516# a_36234_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5314 VSS a_14457_15823# a_14747_7663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5315 VDD ANTENNA__1195__A1.DIODE a_33141_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X5316 a_40250_13508# a_18546_13506# a_40158_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5317 a_16381_35286# a_16745_34427# a_17867_34473# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5318 a_8831_24501# a_8399_18115# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5319 a_32126_63158# pmat.row_n[7] a_32618_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X532 VDD pmat.rowon_n[15] a_51202_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5320 a_40250_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5321 a_37638_20504# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5322 VSS a_7717_14735# a_13275_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X5323 a_27789_36039# a_27049_35515# a_28112_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5324 a_37238_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5325 a_19522_27247# a_7840_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X5326 a_44266_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5327 VSS a_19405_28853# a_31165_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5328 VDD a_29685_34954# a_20534_35431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5329 VDD a_5558_9527# a_5935_6575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X533 VSS pmat.row_n[6] a_19470_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5330 a_28245_35877# a_27789_36039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X5331 VDD a_11965_42583# a_11910_43047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5332 a_27198_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5333 a_10932_21959# a_5899_21807# a_11163_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5334 a_33719_34191# a_33542_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5335 a_1937_48169# a_1769_14735# a_1683_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5336 a_25667_35253# a_11317_36924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5337 a_5320_30199# a_4719_30287# a_5462_30333# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5338 a_1881_74031# a_1846_74283# a_1643_74005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5339 VSS a_6970_67191# a_6612_66933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X534 a_21174_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5340 a_39550_9858# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5341 a_42166_22950# a_18162_22544# a_42258_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5342 a_38150_12910# a_18162_12504# a_38242_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5343 a_13427_18303# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5344 a_34226_68178# a_18546_68220# a_34134_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5345 VSS a_30111_47911# a_45201_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.085e+11p ps=7.38e+06u w=650000u l=150000u M=2
X5346 VSS pmat.row_n[1] a_49590_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5347 a_30473_49871# ANTENNA__1187__B1.DIODE a_30255_49783# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5348 VDD a_14887_46377# a_14699_46377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5349 a_24490_72234# VDD a_24094_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X535 a_23486_60186# pmat.rowon_n[4] a_23090_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5350 a_11455_50237# a_5363_33551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5351 VDD a_2897_21781# a_2927_22134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5352 VDD a_7658_71543# a_7847_73493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5353 vcm a_18162_20536# a_31214_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5354 VSS pmat.row_n[9] a_51598_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5355 VSS a_11261_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5356 vcm a_18162_10496# a_27198_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5357 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5358 a_8443_20719# a_7935_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5359 a_12764_37277# a_12513_36924# a_12543_36950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X536 a_29206_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5360 VSS a_1781_9308# a_1725_11254# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5361 VDD pmat.sample_n a_18162_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X5362 a_32218_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5363 VSS a_9459_5461# a_8703_6202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5364 VSS a_13779_43123# a_13719_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X5365 a_3938_76751# a_2861_76757# a_3776_77129# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5366 VSS a_11067_30287# a_16945_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5367 a_14655_59343# a_10515_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5368 a_45450_48695# a_33423_47695# a_46225_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5369 a_22482_24918# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X537 a_23486_19898# nmat.rowon_n[4] a_23090_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5370 a_16311_28327# a_45915_29941# a_45861_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=2.44e+12p ps=2.288e+07u w=1e+06u l=150000u M=8
X5371 a_19074_23954# a_18162_23548# a_19166_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5372 VDD a_2099_24746# a_1895_23610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5373 a_6082_46831# a_5455_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5374 a_39125_47349# a_38907_47753# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X5375 a_36538_58178# pmat.rowon_n[2] a_36142_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5376 VSS comp.adc_comp_circuit_0.adc_comp_buffer_1.in a_54790_39198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.55e+11p ps=1.62e+06u w=500000u l=150000u
X5377 a_43662_71552# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5378 a_35534_23914# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5379 VDD a_29076_48695# a_28573_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X538 a_4031_40455# a_2935_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X5380 a_39646_61512# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5381 a_6749_66959# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X5382 a_29206_19532# a_18546_19530# a_29114_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5383 VDD a_2007_25597# a_35860_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5384 a_12542_47197# a_11784_47099# a_11979_47068# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5385 a_47278_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5386 a_34611_44265# a_33489_44219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X5387 VDD a_4259_31375# a_9166_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5388 a_9976_58575# a_9577_58229# a_9305_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5389 a_6917_15055# a_6853_14967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X539 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5390 a_5989_34863# a_5823_34863# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5391 a_26102_71190# a_18162_71230# a_26194_71190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5392 VSS a_6639_23413# nmat.sw VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5393 a_25494_15882# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5394 VSS pmat.row_n[10] a_28506_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5395 a_2192_49159# a_2407_49289# a_2334_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5396 a_32522_16886# nmat.rowon_n[7] a_32126_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5397 a_43548_30287# a_41227_29423# a_43442_30287# VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=0p ps=0u w=650000u l=150000u
X5398 VSS ANTENNA__1395__B1.DIODE a_24673_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5399 VDD pmat.rowon_n[15] a_20078_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X54 nmat.col[12] ANTENNA__1184__B1.DIODE a_14471_3561# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X540 a_24586_7452# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5400 VSS a_1643_61493# a_1591_61519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5401 a_28506_8854# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5402 a_20170_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5403 a_44570_69222# pmat.rowon_n[13] a_44174_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5404 vcm a_18162_57174# a_29206_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5405 a_25575_31055# a_25042_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5406 VSS pmat.row_n[10] a_41558_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5407 vcm a_18162_17524# a_51294_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5408 a_33222_55126# a_18546_55168# a_33130_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5409 a_33622_59504# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X541 a_20474_7850# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5410 VDD a_20475_49783# a_20425_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5411 a_29510_14878# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5412 a_34887_39095# a_33765_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5413 a_45270_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5414 a_48190_24958# VDD a_48682_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5415 VDD a_3891_60431# a_3339_59879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X5416 a_38150_57134# a_18162_57174# a_38242_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5417 a_20349_50345# a_18547_51565# a_20267_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5418 VSS a_16505_40157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5419 VDD pmat.rowon_n[14] a_24094_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X542 a_51294_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5420 a_24270_49783# a_22499_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X5421 a_42258_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5422 a_31518_63198# pmat.rowon_n[7] a_31122_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5423 VSS a_11007_58229# a_12155_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5424 VSS a_33765_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5425 a_6777_61519# a_5731_58951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5426 VSS pmat.row_n[9] a_45574_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5427 a_17882_31421# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5428 VDD nmat.rowon_n[6] a_45178_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5429 a_42658_14480# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X543 VSS a_1923_31743# a_4945_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5430 VDD a_12437_28585# a_15393_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5431 VDD a_20572_40517# a_20476_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5432 a_40158_15922# a_18162_15516# a_40250_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5433 a_43262_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5434 a_21082_8894# pmat.row_n[0] a_21574_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5435 a_10907_42390# a_10725_42390# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5436 a_34030_47893# ANTENNA__1197__B.DIODE a_34245_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5437 a_5968_77295# a_5725_76207# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5438 VDD a_2879_26703# a_2007_25597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X5439 a_26456_36165# a_25393_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X544 a_13102_71631# a_13158_71285# a_13102_71311# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5440 VSS pmat.row_n[1] a_35534_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5441 a_31614_8456# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5442 VDD a_28336_29967# a_43359_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5443 a_10016_30511# a_9899_30724# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5444 a_18546_62196# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X5445 a_22482_65206# pmat.rowon_n[9] a_22086_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5446 VSS pmat.row_n[0] a_48586_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5447 a_5266_17143# a_6621_16885# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X5448 a_37238_24552# a_18546_24550# a_37146_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5449 a_50290_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X545 a_2950_74707# a_3267_74817# a_3225_74941# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X5450 VDD nmat.rowon_n[7] a_49194_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5451 a_36234_66170# a_18546_66212# a_36142_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5452 a_46674_13476# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5453 a_43170_10902# pmat.row_n[2] a_43662_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5454 VDD nmat.rowon_n[12] a_50198_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5455 a_20078_63158# a_18162_63198# a_20170_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5456 a_29606_23516# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5457 VDD pmat.rowon_n[12] a_40158_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5458 a_29206_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5459 VSS a_77245_40202# a_77058_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X546 VDD nmat.rowon_n[9] a_37146_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5460 VSS a_2935_38279# a_6800_44629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5461 VDD pmat.rowon_n[2] a_36142_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5462 VDD nmat.rowon_n[2] a_33130_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5463 VDD a_29076_48695# a_29300_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5464 a_33130_62154# a_18162_62194# a_33222_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5465 a_36538_11866# nmat.rowon_n[12] a_36142_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5466 VDD a_29217_41570# a_31976_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5467 a_43971_28487# a_38851_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5468 VDD a_31085_27221# nmat.col[11] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5469 a_1644_62581# a_1591_61519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X547 a_34226_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5470 a_20251_42089# a_20645_42044# a_14149_39747# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X5471 a_11257_60137# a_10878_58487# a_10286_60405# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5472 a_25494_56170# pmat.rowon_n[0] a_25098_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5473 a_19566_15484# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5474 a_39193_43131# a_37960_42693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X5475 vcm a_18162_72234# a_41254_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5476 VDD a_11067_27239# a_22830_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X5477 VDD a_14943_26703# a_16285_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X5478 VSS a_27411_46805# a_14887_46377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5479 VDD nmat.rowon_n[10] a_23090_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X548 a_35230_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5480 VDD a_30663_50087# a_41335_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X5481 vcm a_18162_62194# a_37238_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5482 a_37146_66170# pmat.row_n[10] a_37638_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5483 a_41254_60146# a_18546_60188# a_41162_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5484 a_14633_50095# a_13432_62581# a_14287_50345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X5485 VDD a_47011_31029# a_46339_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u M=3
X5486 VDD pmat.rowon_n[11] a_44174_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5487 a_14369_60137# a_10515_15055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=0p ps=0u w=1e+06u l=150000u
X5488 a_41654_64524# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5489 a_6796_15279# a_6679_15492# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X549 nmat.col_n[3] a_12250_4175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5490 a_34226_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5491 VSS a_44849_45717# a_44783_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5492 VDD a_10139_32117# a_10070_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X5493 a_5747_44905# a_4257_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5494 VSS pmat.row_n[6] a_30514_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5495 VSS a_8197_20871# a_10441_21263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X5496 VSS config_2_in[6] a_1591_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5497 a_5597_69473# a_2419_53351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5498 a_29510_55166# VSS a_29114_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5499 a_11200_42895# a_10949_43124# a_10979_43222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X55 a_1644_65845# a_1591_65327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X550 VDD a_7732_52105# a_7907_52031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5500 a_3609_9295# a_3663_9269# a_3609_9615# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5501 a_44570_22910# nmat.rowon_n[1] a_44174_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5502 a_8643_77129# a_8197_76757# a_8547_77129# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X5503 a_31214_71190# a_18546_71232# a_31122_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5504 a_48586_58178# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5505 a_42166_60146# pmat.row_n[4] a_42658_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5506 a_27198_61150# a_18546_61192# a_27106_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5507 a_50198_68178# a_18162_68218# a_50290_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5508 a_33986_47375# a_32687_46607# a_33986_47695# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X5509 VDD pmat.rowon_n[7] a_31122_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X551 a_3986_74575# a_3228_74691# a_3423_74549# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5510 VSS a_21365_27247# a_31217_29429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5511 VDD a_5257_62215# a_4413_62037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X5512 VSS a_5715_16911# a_5731_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5513 a_35630_55488# pmat.en_bit_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5514 vcm a_18162_23548# a_36234_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5515 a_6817_51733# a_6651_51733# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5516 a_40250_21540# a_18546_21538# a_40158_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5517 a_33870_29967# a_20439_27247# a_33567_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X5518 VDD a_16657_42567# a_17808_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5519 a_2250_59165# a_2163_58941# a_1846_59051# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X552 nmat.rowoff_n[13] a_12447_16143# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X5520 VSS pmat.row_n[15] a_39550_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5521 a_6750_60797# a_4351_55527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5522 a_36234_11500# a_18546_11498# a_36142_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5523 VDD a_12500_68021# a_9545_66567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X5524 a_32126_71190# pmat.row_n[15] a_32618_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5525 vcm a_18162_22544# a_49286_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5526 a_12687_18377# a_12171_18005# a_12592_18365# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X5527 a_28110_61150# pmat.row_n[5] a_28602_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5528 a_37238_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5529 a_49286_10496# a_18546_10494# a_49194_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X553 a_2369_33775# a_2325_34017# a_2203_33775# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5530 VSS pmat.row_n[2] a_35534_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5531 VSS a_38851_28327# a_44023_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5532 a_26576_46831# a_25681_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5533 VSS a_25129_31751# a_25084_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5534 a_26194_22544# a_18546_22542# a_26102_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5535 VSS pmat.row_n[3] a_50594_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5536 a_44174_18934# pmat.row_n[10] a_44666_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5537 VSS VDD a_44570_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5538 a_10239_14183# a_14287_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5539 VSS a_27329_42902# a_27519_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X554 a_24186_58138# a_18546_58180# a_24094_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5540 a_38150_20942# a_18162_20536# a_38242_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5541 VSS pmat.row_n[13] a_33526_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5542 a_30514_66210# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5543 a_35621_27247# a_13091_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5544 VSS a_4075_50087# a_7431_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5545 a_19166_7484# a_18546_7482# a_19074_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5546 a_11568_37277# a_11317_36924# a_11347_36950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X5547 VSS a_22393_37692# a_22085_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X5548 VSS a_33467_46261# a_37791_46811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5549 a_35230_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X555 a_2419_53351# a_3707_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X5550 a_37542_60186# pmat.rowon_n[4] a_37146_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5551 a_37542_19898# nmat.rowon_n[4] a_37146_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5552 a_7415_29397# a_10097_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X5553 a_34226_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5554 a_48282_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5555 VSS pmat.row_n[7] a_47582_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5556 a_21574_18496# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5557 VDD a_6800_22869# a_6830_22895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5558 a_21478_24918# VSS a_21082_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5559 a_3784_62607# a_3305_62607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X556 VSS a_41731_49525# a_21739_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X5560 VDD a_1957_43567# a_12860_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5561 a_51598_13874# nmat.rowon_n[10] a_51202_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5562 a_4193_40303# a_2839_38101# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5563 VSS a_22817_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5564 a_34530_65206# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5565 a_38242_58138# a_18546_58180# a_38150_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5566 a_34626_17492# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5567 VSS a_23815_48981# pmat.row_n[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X5568 a_8175_63669# a_8378_63827# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5569 a_30044_43781# a_28981_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X557 a_48282_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5570 a_32126_18934# a_18162_18528# a_32218_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5571 a_7456_15279# a_6375_15279# a_7109_15521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X5572 VDD a_41665_46805# a_40949_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5573 a_13656_62927# a_13432_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5574 a_48190_58138# pmat.row_n[2] a_48682_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5575 a_3305_17999# a_2847_18303# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X5576 VSS a_4492_32375# a_4123_32661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5577 a_24490_57174# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5578 a_48586_11866# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5579 a_40250_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X558 a_45178_11906# a_18162_11500# a_45270_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5580 VDD a_3305_17999# a_6467_29415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5581 a_7367_31055# a_6743_31061# a_7259_31433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5582 VDD a_28591_36519# a_11149_36924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X5583 a_28202_69182# a_18546_69224# a_28110_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5584 vcm a_18162_66210# a_25190_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5585 a_35138_13914# pmat.row_n[5] a_35630_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5586 a_36234_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5587 a_32405_32463# a_18241_31698# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X5588 VDD nmat.rowon_n[14] a_26102_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5589 a_8908_14967# a_7644_16341# a_9050_14774# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X559 a_34134_19938# pmat.row_n[11] a_34626_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5590 VSS a_2847_8511# a_2781_8585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5591 a_20520_32521# a_19605_32149# a_20173_32117# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5592 a_25590_19500# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5593 a_3320_30333# a_3202_29941# a_3248_30333# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5594 a_6323_26409# a_5320_27023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5595 VDD a_12069_38517# a_12013_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5596 VSS a_33386_30485# a_31675_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5597 a_28506_14878# nmat.rowon_n[9] a_28110_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5598 a_2325_15797# a_2107_16201# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X5599 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X56 VSS a_15299_28879# a_15753_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X560 a_45405_30511# a_41731_49525# a_45212_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=1.195e+12p ps=1.039e+07u w=1e+06u l=150000u M=2
X5600 VSS a_29864_39429# a_29827_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X5601 VSS a_4866_52245# a_4259_73807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5602 vcm a_18162_65206# a_29206_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5603 a_50690_57496# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5604 a_29114_69182# pmat.row_n[13] a_29606_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5605 a_19509_39638# a_19505_38779# a_20627_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5606 a_33222_63158# a_18546_63200# a_33130_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5607 vcm a_18162_60186# a_30210_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5608 VSS pmat.row_n[8] a_37542_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5609 a_33622_67536# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X561 a_5589_14967# a_5451_14557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5610 vcm a_18162_15516# a_47278_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5611 a_30118_64162# pmat.row_n[8] a_30610_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5612 a_4231_60975# a_1591_61519# a_4041_61225# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5613 a_38661_32521# a_37471_32149# a_38552_32521# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5614 a_10497_54697# a_10117_54697# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5615 a_51294_13508# a_18546_13506# a_51202_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5616 VSS a_22186_30485# pmat.en_bit_n[2] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X5617 VSS pmat.row_n[0] a_38546_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5618 a_38150_65166# a_18162_65206# a_38242_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5619 a_5069_40303# a_4955_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X562 VDD a_7644_16341# a_12077_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5620 a_2319_72092# a_2124_72123# a_2629_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X5621 VSS pmat.row_n[15] a_20474_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5622 a_13641_54965# a_13423_55369# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X5623 a_42258_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5624 VSS a_3339_70759# a_6637_69367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5625 VDD a_4351_55527# a_5760_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.5e+11p ps=5.7e+06u w=1e+06u l=150000u
X5626 VSS pmat.row_n[4] a_50594_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5627 a_15667_27239# a_41731_49525# a_44463_29199# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X5628 a_20078_56130# pmat.row_n[0] a_20570_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5629 a_46523_39733# a_44444_32233# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u M=3
X563 VDD a_5423_67191# a_4421_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X5630 a_48586_8854# nmat.rowon_n[15] a_48190_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5631 a_11409_34789# a_10953_34951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X5632 VSS pmat.row_n[14] a_33526_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5633 a_42562_70226# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5634 a_32219_44535# a_31097_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5635 a_24186_15516# a_18546_15514# a_24094_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5636 a_40158_23954# a_18162_23548# a_40250_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5637 a_4319_71311# a_4265_71543# a_4225_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X5638 a_44745_44111# a_31675_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5639 VDD a_7717_14735# a_21279_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X564 a_26329_28111# a_13091_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X5640 ANTENNA__1190__A2.DIODE a_46863_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5641 a_24094_55126# VDD a_24586_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5642 a_25997_42902# a_25209_42043# a_26272_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5643 a_33925_28879# a_13641_23439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5644 a_45574_61190# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5645 a_2107_33775# a_1757_33775# a_2012_33775# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5646 VDD a_5809_51335# a_5731_58951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X5647 VSS a_1586_33927# a_6007_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5648 a_2369_8573# a_2325_8181# a_2203_8585# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5649 a_9651_69679# a_9135_69679# a_9556_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X565 a_24965_50639# a_17139_30503# pmat.col[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X5650 a_9184_51335# a_9457_51163# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5651 a_28202_14512# a_18546_14510# a_28110_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5652 a_28506_71230# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5653 vcm a_18162_11500# a_25190_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5654 VSS a_20616_27791# a_25129_31751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5655 VDD config_1_in[7] a_1591_4399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5656 VDD pmat.rowon_n[10] a_36142_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5657 a_1761_11471# a_1591_11471# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5658 VDD a_4337_22351# a_4509_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5659 a_24490_10862# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X566 vcm a_18162_10496# a_21174_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5660 a_35730_47919# a_35786_47893# a_33957_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5661 pmat.row_n[7] a_17007_50613# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X5662 VDD a_5731_58799# a_3866_57399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5663 a_36234_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5664 vcm a_18162_57174# a_50290_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5665 a_5417_11445# a_5768_9527# a_5921_11791# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5666 VSS pmat.row_n[5] a_22482_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5667 a_49590_60186# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5668 VSS a_47449_52271# ANTENNA__1190__A1.DIODE VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X5669 a_19166_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X567 VSS a_5363_70543# a_7845_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X5670 a_49590_19898# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5671 VSS a_6608_70455# a_6559_70223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5672 a_51202_70186# a_18162_70226# a_51294_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5673 VDD a_13597_37571# a_19509_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5674 vcm a_18162_70226# a_37238_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5675 a_50594_14878# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5676 a_41654_72556# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5677 a_33526_24918# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5678 VSS a_12069_38517# a_12013_38870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5679 pmat.col[24] a_16311_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X568 a_38642_10464# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5680 VSS a_25393_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5681 a_37638_62516# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5682 VSS a_12967_58559# a_11007_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5683 a_28352_50959# a_11067_27239# a_28049_50613# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X5684 a_16025_29469# a_14691_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5685 VDD a_15435_29111# a_12851_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X5686 a_41162_62154# a_18162_62194# a_41254_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5687 VDD pmat.rowon_n[4] a_41162_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5688 vcm a_18162_59182# a_23182_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5689 VSS a_5595_65301# a_6612_65845# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X569 VDD a_2319_69916# a_2250_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X5690 VSS VDD a_27502_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5691 a_20520_32521# a_19439_32149# a_20173_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5692 a_27973_41605# a_28281_41245# a_27947_41245# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5693 VSS pmat.sample_n a_18162_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X5694 a_22273_48169# a_21279_48999# a_22201_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5695 a_24094_72194# a_18162_72234# a_24186_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5696 a_29510_63198# pmat.rowon_n[7] a_29114_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5697 VSS pmat.row_n[4] a_26498_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5698 VSS pmat.row_n[11] a_26498_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5699 a_27789_44743# a_27509_44219# a_28572_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X57 a_5357_30511# a_4167_30511# a_5248_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X570 a_14887_46377# a_27411_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5700 a_23486_16886# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5701 a_13686_13967# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5702 a_6981_21263# a_3351_27249# a_6909_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5703 a_2121_69679# a_1643_69653# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5704 a_28267_50639# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X5705 a_46135_38127# a_45884_38377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X5706 a_78802_39738# a_78898_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5707 VDD pmat.rowoff_n[4] a_44174_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5708 a_15435_29111# a_15543_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5709 a_9201_27907# a_4516_21531# a_9129_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X571 VDD a_10795_47893# a_5363_70543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X5710 vcm a_18162_68218# a_31214_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5711 VDD nmat.rowon_n[1] a_27106_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5712 vcm a_18162_58178# a_27198_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5713 a_20253_46287# a_20076_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5714 VDD pmat.rowon_n[15] a_31122_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5715 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5716 a_10954_73195# a_11271_73085# a_11229_72943# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X5717 a_31214_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5718 a_25190_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5719 a_20570_7452# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X572 VSS a_8175_12533# a_5579_12394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5720 a_2099_8725# a_1979_9334# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5721 a_35230_61150# a_18546_61192# a_35138_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5722 a_39550_68218# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5723 VDD a_82783_53524# pmat.col[31] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5724 VDD VDD a_30118_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5725 a_28202_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5726 a_25098_11906# a_18162_11500# a_25190_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5727 a_19049_41959# a_19145_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5728 VDD nmat.rowon_n[5] a_43170_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5729 a_2882_70045# a_2163_69821# a_2319_69916# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X573 VDD VDD a_28110_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5730 VDD a_2847_28095# a_2834_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5731 a_9581_56079# a_9103_56383# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5732 a_4683_30511# a_4167_30511# a_4588_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X5733 VSS a_15435_29111# a_12851_28853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X5734 a_6749_65871# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X5735 VDD a_10195_59861# a_10153_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5736 VSS a_2219_4943# a_2695_4943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5737 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5738 a_11307_14191# a_10791_14191# a_11212_14191# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X5739 a_79718_39826# vcm.sky130_fd_sc_hd__nand2_1_1.A vcm.sky130_fd_sc_hd__nand2_1_1.Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X574 VSS pmat.row_n[12] a_36538_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5740 a_36142_61150# pmat.row_n[5] a_36634_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5741 a_6981_21263# a_6579_21583# a_6817_21583# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X5742 VSS a_13561_42333# a_13253_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X5743 vcm a_18162_19532# a_26194_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5744 a_6168_18543# a_5087_18543# a_5821_18785# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X5745 a_44174_69182# a_18162_69222# a_44266_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5746 VSS pmat.row_n[1] a_46578_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5747 a_4490_6031# a_3413_6037# a_4328_6409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5748 a_13277_14441# a_10515_13967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X5749 VSS pmat.row_n[11] a_29510_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X575 VDD a_15899_47939# a_24602_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5750 a_33526_65206# pmat.rowon_n[9] a_33130_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5751 a_8547_65161# a_8197_64789# a_8452_65149# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5752 result_out[3] a_1644_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5753 a_47278_66170# a_18546_66212# a_47186_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5754 VDD a_1717_13647# a_8257_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5755 a_30999_48071# a_31675_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5756 a_31339_31787# a_18563_27791# a_38299_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5757 a_39154_9898# pmat.row_n[1] a_39646_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5758 VDD nmat.rowon_n[4] a_47186_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5759 VDD pmat.rowon_n[12] a_51202_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X576 vcm a_18162_19532# a_46274_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5760 a_2121_61885# a_1643_61493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5761 VSS pmat.row_n[3] a_19470_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5762 VSS a_2439_13889# a_2400_13763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5763 VDD a_43776_30287# a_45719_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5764 a_51598_63198# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5765 a_21174_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5766 vcm a_18162_7484# a_41254_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5767 a_23486_57174# pmat.rowon_n[1] a_23090_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5768 a_13331_8585# a_12981_8213# a_13236_8573# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5769 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X577 VDD a_2511_25615# a_1923_31743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X5770 a_12199_62621# a_11797_60431# a_12162_64015# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X5771 a_4866_52245# a_5123_52423# a_5081_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5772 a_49686_9460# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5773 a_13685_55357# a_13641_54965# a_13519_55369# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5774 VDD pmat.rowon_n[7] a_29114_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5775 VSS nmat.sample_n a_18162_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X5776 VDD a_8569_60405# a_6175_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X5777 a_51294_7484# a_18546_7482# a_51202_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5778 a_12053_27497# a_12175_27221# a_11885_27247# VSS sky130_fd_pr__nfet_01v8 ad=2.21e+11p pd=1.98e+06u as=0p ps=0u w=650000u l=150000u
X5779 a_7939_31591# a_1781_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X578 a_22178_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5780 a_6790_77661# a_5713_77295# a_6628_77295# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5781 vcm a_18162_62194# a_48282_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5782 a_48190_66170# pmat.row_n[10] a_48682_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5783 a_7377_14441# a_5266_17143# a_7295_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5784 a_25190_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5785 a_47035_27497# a_17139_30503# a_46817_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5786 a_13239_65161# a_12889_64789# a_13144_65149# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5787 VDD a_2847_8511# a_2021_9563# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5788 vcm a_18162_9492# a_32218_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5789 a_42562_23914# pmat.rowoff_n[15] a_42166_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X579 VSS a_6664_26159# a_33386_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5790 a_24833_40719# a_24667_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5791 VDD a_6283_31591# a_22199_32149# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5792 VDD a_40467_46261# a_11948_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5793 a_42658_56492# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5794 a_35290_44527# a_35113_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5795 a_22086_24958# VDD a_22578_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5796 VDD pmat.rowon_n[13] a_28110_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5797 a_4085_7663# a_3663_9269# a_4003_7663# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5798 VDD a_10589_22351# a_14287_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5799 a_19860_32509# a_7939_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X58 a_50198_22950# pmat.row_n[14] a_50690_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X580 a_28202_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5800 a_13641_23439# a_9528_20407# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5801 a_4036_70741# a_1591_71855# a_4259_70767# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5802 a_28202_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5803 a_25098_56130# a_18162_56170# a_25190_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5804 a_39550_21906# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5805 a_16745_44581# a_13779_43123# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X5806 VSS _1192_.B1 a_26511_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X5807 a_8782_63695# a_8695_63937# a_8378_63827# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5808 a_28810_52521# _1187_.A2 a_28507_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X5809 a_46674_55488# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X581 VSS pmat.row_n[11] a_49590_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5810 VSS VDD a_37542_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5811 a_26102_23954# pmat.row_n[15] a_26594_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5812 a_30771_39425# a_23821_35279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5813 a_39581_48841# a_38391_48469# a_39472_48841# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5814 a_26102_19938# a_18162_19532# a_26194_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5815 a_30118_72194# VDD a_30610_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5816 vcm a_18162_23548# a_47278_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5817 a_41558_70226# pmat.rowon_n[14] a_41162_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5818 a_30610_21508# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5819 VSS a_7355_37013# a_7289_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X582 VSS a_4068_25615# a_6634_26133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5820 a_29606_65528# pmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5821 a_30210_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5822 a_51294_21540# a_18546_21538# a_51202_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5823 a_47278_11500# a_18546_11498# a_47186_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5824 VSS a_9889_10681# a_9823_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5825 a_37739_43177# a_36617_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5826 a_29114_55126# a_18162_55166# a_29206_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5827 a_19470_24918# VSS a_19074_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5828 VDD a_11339_39319# a_11327_39087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5829 cgen.dlycontrol2_in[2] a_1591_40303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X583 a_40105_47375# a_39647_47679# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X5830 a_49590_13874# nmat.rowon_n[10] a_49194_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5831 a_7109_15521# a_6891_15279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X5832 a_20570_13476# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5833 VSS pmat.row_n[2] a_46578_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5834 a_19566_57496# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5835 VDD VSS a_23090_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5836 a_29114_14918# pmat.row_n[6] a_29606_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5837 VSS pmat.row_n[12] a_29510_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5838 a_24186_23548# a_18546_23546# a_24094_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5839 a_9783_67075# a_9643_66389# a_9687_67075# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X584 a_29124_37253# a_29220_37253# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X5840 a_33622_12472# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5841 nmat.col[1] _1196_.B1 VSS VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=0p ps=0u w=650000u l=150000u M=2
X5842 a_2557_53181# a_1923_53055# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5843 a_31122_13914# a_18162_13508# a_31214_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5844 VDD a_11067_16359# a_14103_15936# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X5845 a_51202_63158# pmat.row_n[7] a_51694_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5846 a_29220_37253# a_28061_36965# a_29183_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X5847 VSS pmat.row_n[4] a_19470_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5848 a_23486_10862# nmat.rowon_n[13] a_23090_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5849 VDD a_4991_69831# a_13553_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X585 a_17131_48579# a_12263_50959# a_17049_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5850 a_13549_74549# a_13331_74953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X5851 VSS a_10423_16055# a_10423_15823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5852 a_3056_9839# a_2972_9991# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5853 VSS a_15049_36374# a_14113_36604# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X5854 a_46274_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5855 a_48586_60186# pmat.rowon_n[4] a_48190_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5856 vcm a_18162_61190# a_24186_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5857 a_48586_19898# nmat.rowon_n[4] a_48190_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5858 a_32740_50095# a_32514_50141# a_32371_50247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5859 VDD a_3688_17179# a_8649_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X586 VDD a_4383_7093# a_11209_17782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X5860 VSS a_7779_22583# a_8356_23671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5861 a_32126_9898# a_18162_9492# a_32218_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5862 a_46947_39215# a_46705_38671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X5863 a_23604_39655# a_22541_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X5864 a_16926_46261# a_12447_16143# a_17234_46403# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5865 a_32618_18496# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5866 a_36234_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5867 VDD a_33281_49551# a_10883_3303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=6
X5868 vcm a_18162_65206# a_50290_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5869 a_50198_69182# pmat.row_n[13] a_50690_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X587 a_4801_69679# a_1823_74557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X5870 a_14471_29673# a_14466_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5871 a_49286_58138# a_18546_58180# a_49194_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5872 a_29051_39783# a_23821_35279# a_29225_39659# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5873 a_22482_58178# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5874 a_14065_22671# a_14005_22589# a_13962_22671# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X5875 a_36538_71230# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5876 a_3413_6037# a_3247_6037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5877 VDD a_19405_28853# a_19351_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5878 VSS a_5411_12167# a_5363_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5879 a_35534_57174# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 a_83005_26159# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X5880 vcm a_18162_10496# a_46274_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5881 a_37638_70548# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5882 a_4871_17429# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X5883 VDD a_1643_31573# a_1591_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5884 a_18660_47607# a_16083_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X5885 vcm a_18162_67214# a_23182_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5886 a_2999_76922# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5887 a_3410_66003# a_3688_65987# a_3644_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5888 a_26889_47073# a_26671_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X5889 a_37146_60146# a_18162_60186# a_37238_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X589 vcm a_18162_7484# a_45270_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5890 a_26583_34343# cgen.dlycontrol1_in[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X5891 a_18235_35831# a_17113_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5892 VSS a_2791_57703# a_5329_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5893 a_51294_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5894 VSS a_4921_32441# a_4855_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5895 a_47278_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5896 a_17959_44265# a_17996_44007# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X5897 VDD a_40628_39429# a_39781_40157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X5898 vcm a_18162_12504# a_19166_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5899 a_41558_24918# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X59 a_31923_42367# cgen.dlycontrol4_in[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X590 a_26102_22950# a_18162_22544# a_26194_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5900 a_23021_29199# a_20616_27791# a_23033_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5901 a_16761_51183# a_11067_16359# a_16679_51183# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5902 a_1775_5059# a_1761_2767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5903 a_37542_7850# VDD a_37146_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5904 a_11021_42619# a_13985_41317# a_15107_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5905 a_3092_72399# a_2655_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5906 a_23182_10496# a_18546_10494# a_23090_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5907 VDD a_3123_27399# a_2743_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X5908 a_14565_16911# a_11067_16359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5909 a_4719_58255# a_2419_69455# a_4897_58575# VSS sky130_fd_pr__nfet_01v8 ad=5.07e+11p pd=5.46e+06u as=0p ps=0u w=650000u l=150000u
X591 VSS pmat.row_n[3] a_39550_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5910 a_26276_39429# a_25117_39141# a_26239_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5911 VSS pmat.row_n[1] a_42562_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5912 VDD a_22043_35041# a_21867_34709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5913 a_38546_68218# pmat.rowon_n[12] a_38150_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5914 vcm a_18162_16520# a_45270_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5915 a_48282_19532# a_18546_19530# a_48190_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5916 a_33436_34191# a_33259_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5917 a_11980_3087# _1184_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5918 a_31122_58138# a_18162_58178# a_31214_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5919 a_44570_15882# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X592 a_3325_23439# a_2847_23743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5920 VSS a_3923_68021# a_3069_69367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5921 ANTENNA__1395__B1.DIODE a_45019_38645# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=8
X5922 a_11927_27399# a_13151_23957# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X5923 a_21147_49525# a_20619_49551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X5924 a_20476_40517# a_19413_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5925 VDD a_4167_9615# a_4169_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5926 a_28506_9858# nmat.rowon_n[14] a_28110_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5927 a_31122_17930# pmat.row_n[9] a_31614_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5928 VSS pmat.row_n[15] a_31518_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5929 VDD a_20520_32521# a_20695_32447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X593 VDD a_21063_48723# a_10515_13967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X5930 a_31097_44581# a_30641_44743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X5931 VSS a_5245_56053# a_3967_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X5932 a_28202_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5933 VDD a_1591_69679# a_3123_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X5934 VDD pmat.rowon_n[5] a_35138_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5935 a_24643_51959# a_13459_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X5936 a_22178_16520# a_18546_16518# a_22086_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5937 a_12557_32441# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5938 a_15163_32375# pmat.rowon_n[7] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5939 VDD a_36663_34191# a_36769_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X594 vcm a_18162_16520# a_20170_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5940 a_5161_40553# a_4955_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5941 VSS a_1923_53055# a_2433_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5942 VSS a_28981_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5943 a_39246_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5944 VSS pmat.row_n[7] a_21478_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5945 a_24490_18894# nmat.rowon_n[5] a_24094_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5946 VDD a_1586_50247# a_7479_53909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5947 VDD a_6639_63927# a_4266_63303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X5948 a_11883_62063# a_5651_66975# a_11798_62063# VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X5949 a_43566_62194# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X595 a_23182_19532# a_18546_19530# a_23090_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5950 a_11207_11079# comp_latch VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5951 a_50594_63198# pmat.rowon_n[7] a_50198_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5952 VDD pmat.rowon_n[4] a_39154_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5953 VDD a_10515_61839# a_14125_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u M=4
X5954 a_35138_55126# pmat.en_bit_n[2] a_35630_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5955 VSS a_33869_31599# a_35084_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5956 a_13697_47349# a_13830_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X5957 a_25190_57134# a_18546_57176# a_25098_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5958 a_25409_29245# a_25325_29125# a_25327_28992# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5959 a_22086_58138# pmat.row_n[2] a_22578_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X596 a_30210_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5960 VSS pmat.row_n[6] a_25494_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5961 a_22482_11866# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5962 a_19074_10902# a_18162_10496# a_19166_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5963 VSS a_6651_33239# a_2046_30184# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5964 a_44666_24520# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5965 a_36485_49007# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5966 a_17845_27791# a_7415_29397# a_18035_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5967 VSS a_7026_24527# a_17323_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5968 a_35534_10862# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5969 a_2886_25398# a_2648_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X597 a_41254_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5970 a_2834_40847# a_1757_40853# a_2672_41225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5971 VDD a_45450_48695# a_45502_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u M=4
X5972 VDD pmat.rowon_n[15] a_29114_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5973 a_47278_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5974 a_28078_29967# a_27001_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5975 a_44917_43023# a_44733_44431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X5976 a_2893_38377# a_2839_38101# a_2283_39189# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5977 a_34797_27791# a_34204_27765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X5978 vcm a_18162_70226# a_48282_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5979 VDD VSS a_21082_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X598 a_43566_57174# pmat.rowon_n[1] a_43170_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5980 VSS a_10239_14183# a_14718_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X5981 a_48682_23516# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5982 a_45178_20942# pmat.row_n[12] a_45670_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5983 a_25139_27497# _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X5984 a_45178_16926# a_18162_16520# a_45270_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5985 a_48282_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5986 a_12700_16367# a_11619_16367# a_12353_16609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5987 VDD a_1586_8439# a_2327_11477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5988 VSS a_2651_8916# a_1949_9308# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5989 a_22541_38779# a_22085_38550# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X599 a_5972_51433# a_2389_45859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5990 a_4893_63151# a_4583_68021# a_4509_62037# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5991 VSS a_7026_24527# a_13641_23439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5992 VSS a_37709_52245# pmat.col[18] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5993 a_27249_27791# ANTENNA__1197__B.DIODE nmat.col_n[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5994 vcm a_18162_15516# a_21174_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5995 a_44570_56170# pmat.rowon_n[0] a_44174_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5996 a_2012_39037# a_1895_38842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5997 a_38642_15484# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5998 a_38546_21906# nmat.rowon_n[2] a_38150_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5999 a_12289_46831# a_11910_47197# a_12217_46831# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X6 a_37146_61150# pmat.row_n[5] a_37638_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X60 a_43262_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X600 a_37638_16488# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6000 a_35138_72194# a_18162_72234# a_35230_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6001 VDD nmat.rowon_n[10] a_42166_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6002 a_27502_66210# pmat.rowon_n[10] a_27106_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6003 a_40954_29423# a_17842_27497# a_40868_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6004 VSS a_4984_41935# a_5558_41935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6005 VDD pmat.rowoff_n[15] a_25098_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6006 a_24015_36911# cgen.dlycontrol3_in[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6007 a_8264_11703# a_8472_11739# a_8406_11837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6008 a_22578_20504# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6009 a_22178_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X601 a_3026_20541# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X6010 a_49194_15922# a_18162_15516# a_49286_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6011 a_25098_64162# a_18162_64202# a_25190_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6012 result_out[4] a_1644_59861# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6013 VSS a_82787_54421# _1179_.X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X6014 pmat.rowoff_n[12] a_10055_31591# a_16879_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6015 a_10781_42869# a_31783_42689# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6016 a_2555_49007# a_2407_49289# a_2192_49159# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6017 a_4801_58255# a_4720_58487# a_4719_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6018 a_9463_53511# a_10455_53387# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X6019 a_39154_11906# pmat.row_n[3] a_39646_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X602 a_33309_36039# a_33489_36603# a_34552_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6020 a_4259_65103# a_1591_65327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6021 VSS a_10379_8439# a_9731_8439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6022 a_29768_39429# a_29864_39429# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X6023 VDD nmat.rowon_n[9] a_28110_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6024 VSS a_9213_53903# a_10217_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X6025 a_50290_71190# a_18546_71232# a_50198_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6026 a_26194_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6027 a_7026_74358# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6028 a_23090_12910# a_18162_12504# a_23182_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6029 a_46274_61150# a_18546_61192# a_46182_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X603 a_12821_69929# a_12067_67279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X6030 comp.adc_inverter_1.out comp.adc_inverter_1.in VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6031 a_29114_63158# a_18162_63198# a_29206_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6032 a_9369_59915# a_1769_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6033 VSS a_4075_31591# a_13620_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6034 VDD pmat.rowon_n[12] a_49194_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6035 a_10913_55535# a_10497_54697# a_11004_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6036 a_10400_15279# a_9485_15279# a_10053_15521# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X6037 VDD pmat.rowon_n[7] a_50198_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6038 a_9747_62985# a_9301_62613# a_9651_62985# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X6039 a_15259_31029# clk_ena VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X604 VSS a_3399_24787# a_2952_25045# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X6040 a_29606_10464# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6041 VDD _1179_.X a_24946_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X6042 VSS pmat.row_n[2] a_44570_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6043 a_51202_71190# pmat.row_n[15] a_51694_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6044 VSS pmat.row_n[12] a_27502_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6045 a_47186_61150# pmat.row_n[5] a_47678_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6046 VDD a_4031_53034# a_3496_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X6047 VSS a_4339_27804# a_10515_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6048 VDD a_3325_40847# a_3659_39733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6049 a_38150_19938# pmat.row_n[11] a_38642_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X605 VDD a_10697_75218# a_10383_75637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.646e+11p ps=2.94e+06u w=420000u l=150000u
X6050 a_12069_38517# a_29023_38571# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6051 a_4327_60975# a_2727_58470# a_4231_60975# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X6052 a_19860_32509# a_7939_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X6053 VSS a_44774_40821# a_45921_42167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6054 a_21478_58178# pmat.rowon_n[2] a_21082_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6055 vcm a_18162_8488# a_21174_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6056 a_35534_71230# pmat.rowon_n[15] a_35138_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6057 VSS a_9545_66567# a_9493_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6058 a_31469_40726# a_30913_39867# a_31976_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6059 a_45270_22544# a_18546_22542# a_45178_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X606 a_26498_67214# pmat.rowon_n[11] a_26102_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6060 VDD pmat.rowon_n[8] a_27106_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6061 a_24586_61512# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6062 a_32218_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6063 a_5423_30485# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6064 a_31214_8488# a_18546_8486# a_31122_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6065 VSS a_12044_49641# a_13290_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6066 a_18546_65208# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X6067 VSS a_24867_53135# a_30479_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X6068 a_12162_39631# a_12116_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6069 a_42683_32375# a_40837_46261# a_42857_32481# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X607 VDD pmat.rowon_n[7] a_49194_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6070 ndecision_finish comp.adc_nor_latch_0.NOR_1/A a_55770_39250# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6071 a_39550_70226# pmat.rowon_n[14] a_39154_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6072 a_1857_35113# a_1770_35015# a_1775_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6073 a_46886_51433# _1196_.B1 a_46804_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6074 a_40650_18496# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6075 a_40554_24918# VSS a_40158_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6076 a_28602_60508# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6077 VSS _0467_ a_16965_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6078 VDD a_12219_63303# a_12076_62839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6079 a_18546_14510# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X608 a_1757_26159# a_1591_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6080 a_50198_14918# pmat.row_n[6] a_50690_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6081 VDD a_10055_31591# pmat.rowoff_n[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6082 a_51202_18934# a_18162_18528# a_51294_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6083 a_33130_24958# VDD a_33622_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6084 VSS a_9411_2215# a_31307_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6085 VSS a_1643_65301# a_1591_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6086 a_9112_65161# a_8031_64789# a_8765_64757# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6087 a_23090_57134# a_18162_57174# a_23182_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6088 vcm a_18162_20536# a_19166_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6089 a_6803_77269# a_6628_77295# a_6982_77295# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X609 vcm a_18162_15516# a_33222_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6090 VSS pmat.row_n[9] a_39550_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6091 VSS a_6553_53047# a_5784_52423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6092 a_3491_19465# a_3045_19093# a_3395_19465# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X6093 a_43566_15882# pmat.rowoff_n[7] a_43170_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6094 a_26498_67214# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6095 VDD a_28867_40871# a_13909_39605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X6096 a_6750_60470# a_4351_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X6097 VSS pmat.row_n[9] a_30514_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6098 VDD a_2972_9991# a_2973_10089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6099 vcm a_18162_24552# a_45270_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X61 a_40158_55126# a_18162_55166# a_40250_55126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X610 a_8091_54281# a_7645_53909# a_7995_54281# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X6100 VDD a_43720_32143# a_46978_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6101 VDD nmat.rowon_n[6] a_30118_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6102 a_5173_45993# a_2389_45859# a_5173_45743# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6103 vcm a_18162_66210# a_44266_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6104 a_44666_58500# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6105 VSS pmat.row_n[1] a_20474_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6106 a_11995_20291# a_11803_20535# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6107 a_47582_14878# nmat.rowon_n[9] a_47186_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6108 VSS pmat.row_n[3] a_44570_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6109 VDD a_10515_61839# a_14379_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X611 a_7799_59887# a_5682_56311# a_7436_60039# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6110 VSS pmat.row_n[0] a_33526_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6111 VDD a_1899_35051# a_5353_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X6112 VDD a_23821_35279# a_29051_37607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6113 a_27106_15922# pmat.row_n[7] a_27598_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6114 VSS pmat.row_n[13] a_27502_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6115 a_22178_24552# a_18546_24550# a_22086_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6116 a_13763_67191# a_3615_71631# a_13909_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X6117 a_21174_66170# a_18546_66212# a_21082_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6118 a_31614_13476# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6119 a_4767_24310# a_4339_27804# a_4308_24135# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X612 a_39169_47741# a_39125_47349# a_39003_47753# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6120 a_15747_50069# a_16083_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6121 VDD pmat.rowon_n[2] a_21082_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6122 VSS pmat.row_n[1] a_50594_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6123 a_48190_8894# pmat.row_n[0] a_48682_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6124 VDD a_20173_32117# a_20063_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6125 a_14458_4399# ANTENNA__1190__B1.DIODE a_14289_4649# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6126 VDD a_5768_9527# a_5445_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6127 a_21478_11866# nmat.rowon_n[12] a_21082_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6128 VSS a_5749_30265# a_5683_30333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6129 a_46950_43719# a_46936_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X613 a_9773_47753# a_8583_47381# a_9664_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6130 a_25190_65166# a_18546_65208# a_25098_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6131 vcm a_18162_62194# a_22178_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6132 a_25590_69544# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6133 a_22086_66170# pmat.row_n[10] a_22578_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6134 vcm a_18162_17524# a_39246_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6135 a_9414_63695# a_8656_63811# a_8851_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6136 a_13798_22351# a_11337_25071# a_14065_22671# VSS sky130_fd_pr__nfet_01v8 ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u w=650000u l=150000u
X6137 VDD a_15259_31029# a_5535_29980# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6138 VSS config_1_in[4] a_1591_14735# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X6139 a_43262_15516# a_18546_15514# a_43170_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X614 a_10053_15521# a_9835_15279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X6140 vcm a_18162_12504# a_40250_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6141 vcm a_18162_61190# a_35230_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6142 VSS a_14943_26703# a_16131_29429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6143 VDD a_37129_36130# a_36193_35805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X6144 a_10975_67503# a_10499_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X6145 a_43999_52521# a_23395_53135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X6146 VSS a_42024_46805# a_42703_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X6147 a_21365_27247# a_11927_27399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X6148 a_47278_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6149 a_26102_65166# pmat.row_n[9] a_26594_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X615 VSS a_4976_16091# a_9237_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X6150 VDD a_10239_14183# pmat.rowon_n[11] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6151 VDD a_27947_41245# a_27973_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6152 VDD a_13503_43421# a_13529_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X6153 VDD nmat.rowon_n[15] a_35138_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6154 a_47582_71230# pmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6155 a_33526_58178# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6156 vcm a_18162_11500# a_44266_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6157 a_45178_24958# a_18162_24552# a_45270_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6158 VSS a_24719_39605# a_14589_40726# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6159 VSS a_5423_69367# a_4265_71543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X616 a_45270_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6160 a_7068_11703# a_7276_11739# a_7210_11837# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6161 a_41558_8854# nmat.rowon_n[15] a_41162_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6162 a_20570_55488# pmat.en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6163 a_26498_20902# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6164 a_48190_60146# a_18162_60186# a_48282_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6165 vcm a_18162_23548# a_21174_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6166 VSS pmat.row_n[5] a_41558_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6167 a_29114_56130# pmat.row_n[0] a_29606_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6168 a_2972_9991# a_4865_8181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6169 a_38242_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X617 VDD a_4843_54826# a_4675_54599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X6170 a_7085_15055# a_5266_17143# a_7001_15055# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X6171 a_19746_28111# a_12987_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6172 VSS pmat.row_n[15] a_24490_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6173 a_21174_11500# a_18546_11498# a_21082_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6174 a_33622_8456# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6175 a_21124_39655# a_19965_39867# a_21028_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X6176 a_12375_42895# a_12198_42895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6177 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X6178 VDD nmat.rowon_n[12] a_38150_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6179 vcm a_18162_22544# a_34226_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X618 a_2847_8511# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6180 a_22178_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6181 a_49194_23954# a_18162_23548# a_49286_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6182 a_38905_28853# a_38727_32447# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6183 VSS pmat.row_n[2] a_20474_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6184 a_34226_10496# a_18546_10494# a_34134_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6185 VSS a_2319_67740# a_2250_67869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6186 a_10751_71543# a_10699_72943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X6187 vcm a_18162_59182# a_42258_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6188 VDD a_8695_63937# a_8656_63811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6189 a_35244_32411# a_46130_34319# a_46994_34639# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X619 VDD a_36571_44527# a_36677_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6190 VSS pmat.row_n[4] a_45574_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6191 a_42562_16886# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6192 VSS pmat.row_n[11] a_45574_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6193 VDD a_2672_18377# a_2847_18303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6194 VDD a_18169_31353# a_18199_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6195 VSS pmat.row_n[14] a_28506_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6196 a_40158_10902# a_18162_10496# a_40250_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6197 a_2025_5059# a_1761_2767# a_1953_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6198 a_26194_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6199 a_23090_20942# a_18162_20536# a_23182_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X62 VDD a_2847_18303# a_3305_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X620 a_42166_9898# pmat.row_n[1] a_42658_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6200 a_6895_48981# a_6720_49007# a_7074_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6201 a_9240_60751# a_5651_66975# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=0p ps=0u w=650000u l=150000u M=2
X6202 VSS a_13973_66933# a_13919_65871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6203 vcm a_18162_58178# a_46274_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6204 a_12605_29199# a_10957_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X6205 VDD pmat.rowon_n[15] a_50198_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6206 ANTENNA__1197__A.DIODE a_47407_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6207 a_34063_27791# a_34204_27765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X6208 a_2215_43023# a_1591_43029# a_2107_43401# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X6209 a_20170_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X621 a_1642_26935# a_1738_26677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6210 VDD pmat.rowon_n[5] a_46182_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6211 a_31976_39655# a_30913_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6212 VDD a_44870_48437# a_21279_48999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.65e+12p ps=1.53e+07u w=1e+06u l=150000u M=4
X6213 a_22482_60186# pmat.rowon_n[4] a_22086_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6214 a_19166_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6215 a_22482_19898# nmat.rowon_n[4] a_22086_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6216 a_2939_45503# a_2764_45577# a_3118_45565# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6217 a_50290_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6218 a_28506_17890# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6219 a_33222_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X622 VDD a_15101_29423# a_28803_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.64e+12p ps=1.528e+07u w=1e+06u l=150000u M=2
X6220 a_19166_71190# a_18546_71232# a_19074_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6221 VSS pmat.row_n[7] a_32522_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6222 a_42029_47919# a_33467_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=2.99e+06u as=0p ps=0u w=650000u l=150000u
X6223 VSS a_27947_41245# a_27913_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X6224 a_13549_8181# a_13331_8585# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6225 a_38150_68178# a_18162_68218# a_38242_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6226 VDD VSS a_19074_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6227 a_12431_69367# a_12789_68021# a_12581_69455# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X6228 a_2744_25223# a_2683_22089# a_2886_25398# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X6229 VDD a_13091_28327# a_23033_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X623 VDD a_7663_27247# a_7840_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6230 a_23182_58138# a_18546_58180# a_23090_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6231 vcm a_18162_55166# a_20170_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6232 a_44174_11906# a_18162_11500# a_44266_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6233 a_10781_76029# a_9581_73487# a_10675_76029# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.596e+11p ps=1.6e+06u w=420000u l=150000u
X6234 a_20078_59142# pmat.row_n[3] a_20570_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6235 VDD a_40125_31029# a_37820_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u M=2
X6236 a_5012_10927# a_4989_11079# a_4998_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6237 a_6883_51335# a_6979_51157# a_7281_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6238 a_33130_58138# pmat.row_n[2] a_33622_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6239 a_33526_11866# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X624 a_42166_24958# VDD a_42658_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6240 a_1643_74005# a_1846_74283# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6241 VDD VDD a_27106_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6242 VSS pmat.row_n[12] a_35534_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6243 a_17478_46805# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6244 VDD ANTENNA__1195__A1.DIODE a_26425_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X6245 a_21174_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6246 a_6829_47375# a_6787_47607# a_6723_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6247 a_4149_44431# a_2659_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X6248 a_14287_10927# a_10239_14183# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X6249 VSS pmat.row_n[11] a_48586_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X625 VDD pmat.rowon_n[13] a_48190_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6250 a_45574_64202# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6251 a_7206_5853# a_6487_5629# a_6643_5724# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X6252 a_44082_31599# a_35244_32411# a_43913_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6253 a_43170_21946# pmat.row_n[13] a_43662_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6254 a_43170_17930# a_18162_17524# a_43262_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6255 VDD a_3981_6005# a_3871_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X6256 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X6257 a_2509_34863# a_2467_35015# a_1770_35015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X6258 a_8914_54269# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6259 a_9668_10651# a_9655_6335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X626 a_46229_37583# a_45187_38129# ANTENNA__1395__B1.DIODE VDD sky130_fd_pr__pfet_01v8_hvt ad=2.44e+12p pd=2.288e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=8
X6260 a_50198_63158# a_18162_63198# a_50290_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6261 a_23788_38341# a_22725_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6262 a_37680_42919# a_36345_42567# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6263 VSS pmat.row_n[3] a_38546_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6264 a_10383_75637# a_10697_75218# a_10781_76029# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6265 a_44849_45717# a_29937_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6266 a_40250_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6267 a_42562_57174# pmat.rowon_n[1] a_42166_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6268 VSS a_19413_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X6269 a_4429_76751# a_3951_77055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X627 a_1643_31573# a_1846_31851# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6270 a_36634_16488# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6271 a_18546_22542# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X6272 a_20627_38825# a_19509_39638# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6273 a_24861_52047# a_13459_28111# a_24643_51959# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6274 a_25494_67214# pmat.rowon_n[11] a_25098_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6275 a_2163_56765# a_1586_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6276 VSS pmat.row_n[8] a_22482_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6277 vcm a_18162_15516# a_32218_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6278 VDD a_18243_28327# a_41703_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6279 VSS a_43548_30287# a_43776_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X628 a_24867_53135# a_46211_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X6280 a_49686_15484# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6281 a_45557_52521# _1224_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X6282 a_11893_71427# a_8491_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6283 a_36722_27791# a_25695_28111# a_36419_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X6284 a_42701_31849# a_26479_32117# a_42955_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X6285 a_3303_33609# a_2953_33237# a_3208_33597# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X6286 a_10249_64239# a_5363_70543# a_10167_64239# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6287 a_23090_65166# a_18162_65206# a_23182_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6288 VDD a_10239_14183# a_14289_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X6289 a_14195_11791# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X629 a_4025_54965# a_6559_53903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6290 a_39550_55166# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6291 VSS a_4259_31375# a_9084_51843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6292 a_1927_43541# a_2263_43719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X6293 a_6747_25731# a_6641_25731# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6294 VSS a_20475_49783# a_32411_49559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6295 a_8907_48437# a_9839_47679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6296 a_33765_38053# a_30431_37683# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X6297 a_10494_77547# a_10772_77563# a_10728_77661# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6298 VDD pmat.rowoff_n[7] a_26102_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6299 a_4441_74281# a_4601_74005# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_26194_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X630 a_83217_4649# _1224_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X6300 VDD a_11115_71285# a_11054_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X6301 a_41162_24958# VDD a_41654_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6302 VDD a_10478_25045# a_9075_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6303 VSS a_28812_29575# a_29968_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6304 a_44266_62154# a_18546_62196# a_44174_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6305 a_12471_40214# a_12289_40214# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6306 VDD pmat.rowon_n[13] a_47186_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6307 a_44666_66532# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6308 a_29455_31293# a_30603_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6309 a_3859_23699# a_2835_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X631 a_44789_39215# a_30663_50087# a_44371_39215# VSS sky130_fd_pr__nfet_01v8 ad=8.71e+11p pd=9.18e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X6310 a_19470_58178# pmat.rowon_n[2] a_19074_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6311 a_42658_9460# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6312 VDD a_35499_28023# nmat.col_n[15] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X6313 a_44174_56130# a_18162_56170# a_44266_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6314 a_6971_60797# a_6451_67655# a_6608_60663# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6315 VSS a_10287_24759# a_9777_26935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X6316 a_30514_61190# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6317 VDD a_9463_8439# a_8243_7290# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X6318 a_27106_66170# a_18162_66210# a_27198_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6319 a_41274_28995# a_24747_29967# a_41192_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X632 a_48282_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6320 a_27598_11468# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6321 VSS a_2648_29397# a_6641_8527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6322 a_20170_7484# a_18546_7482# a_20078_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6323 a_11345_70773# a_11115_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6324 VDD pmat.rowon_n[10] a_21082_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6325 a_48682_65528# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6326 a_45178_62154# pmat.row_n[6] a_45670_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6327 a_77882_40202# a_77978_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6328 VDD nmat.rowon_n[14] a_28110_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6329 a_3045_19093# a_2879_19093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X633 a_45178_56130# a_18162_56170# a_45270_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6330 VDD a_22085_38550# a_23420_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6331 VDD a_7343_16042# a_6679_15492# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X6332 a_21174_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6333 a_82998_2473# _1224_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.3e+11p pd=5.26e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6334 a_22657_50345# a_22499_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6335 VSS pmat.row_n[13] a_35534_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6336 a_34530_60186# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6337 a_34530_19898# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6338 a_41663_47893# a_42191_48071# a_42029_47919# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X6339 vcm a_18162_70226# a_22178_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X634 a_4043_59861# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X6340 a_1846_56875# a_2124_56891# a_2080_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6341 a_38642_57496# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6342 VDD VSS a_42166_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6343 a_30913_38779# a_29864_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X6344 VSS pmat.row_n[12] a_48586_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6345 vcm a_18162_20536# a_40250_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6346 a_43262_23548# a_18546_23546# a_43170_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6347 VDD pmat.rowon_n[9] a_25098_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6348 a_39246_13508# a_18546_13506# a_39154_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6349 a_8179_71689# a_7829_71317# a_8084_71677# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X635 VSS a_2411_33749# a_9701_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6350 a_22578_62516# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6351 VSS a_1739_47893# a_1769_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6352 a_46578_71230# pmat.rowon_n[15] a_46182_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6353 a_10898_77661# a_10772_77563# a_10494_77547# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6354 a_25190_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6355 VDD a_14719_37737# a_15737_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X6356 a_44453_53135# _1224_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6357 VSS pmat.row_n[4] a_38546_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6358 a_21028_39655# a_19965_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6359 a_5518_60431# a_4843_54826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X636 a_34887_40183# a_33765_40229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X6360 a_26283_42325# a_11041_40948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6361 a_42562_10862# nmat.rowon_n[13] a_42166_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6362 a_16837_42043# a_15420_41831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X6363 a_25590_14480# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6364 a_25494_20902# pmat.rowoff_n[12] a_25098_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6365 a_38531_51348# a_38575_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6366 a_31393_31055# a_31210_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6367 a_10811_77437# a_7658_71543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6368 a_23700_39655# a_22541_39867# a_23663_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X6369 a_9221_65161# a_8031_64789# a_9112_65161# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X637 a_28110_66170# a_18162_66210# a_28202_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6370 VDD pmat.rowon_n[0] a_28110_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6371 a_20474_69222# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6372 VDD a_7163_53333# a_7067_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6373 a_13546_5263# ANTENNA__1187__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X6374 VDD a_34553_42658# a_33617_42333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X6375 a_51694_18496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6376 a_51598_24918# VSS a_51202_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6377 a_20874_30511# a_1858_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6378 a_6608_60663# a_6451_67655# a_6750_60470# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X6379 pmat.col[7] a_16311_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X638 a_14947_26159# a_14696_26409# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6380 VSS a_30140_43781# a_30103_43447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6381 VSS a_1643_58773# a_1591_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6382 a_10957_14191# a_10791_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6383 VDD a_23700_44869# a_23604_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6384 a_26102_10902# pmat.row_n[2] a_26594_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6385 VSS pmat.row_n[10] a_37542_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6386 a_4549_34685# a_4514_34451# a_4227_34293# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6387 a_41558_58178# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6388 a_20170_61150# a_18546_61192# a_20078_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6389 a_41558_16886# nmat.rowon_n[7] a_41162_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X639 VSS pmat.sample a_18546_72236# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X6390 a_2944_56872# a_3514_57167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6391 a_28770_29673# a_28704_29568# a_28456_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=8.5e+11p ps=5.7e+06u w=1e+06u l=150000u
X6392 a_24490_68218# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6393 a_6583_61519# a_5535_57993# a_6777_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X6394 VDD pmat.rowon_n[2] a_19074_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6395 VDD a_26459_42657# a_26283_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6396 VDD a_7387_33231# a_6283_31591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X6397 vcm a_18162_67214# a_42258_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6398 a_19470_11866# nmat.rowon_n[12] a_19074_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6399 a_9089_12925# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X64 VDD a_41427_31599# a_41427_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X640 a_28602_9460# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6400 a_9919_10422# a_9668_10651# a_9460_10615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X6401 a_33785_30287# a_13641_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X6402 a_2107_41225# a_1591_40853# a_2012_41213# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X6403 vcm a_18162_57174# a_38242_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6404 a_37146_7890# VDD a_37638_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6405 a_10979_42390# a_10949_42364# a_10907_42390# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X6406 a_42258_55126# a_18546_55168# a_42166_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6407 a_39154_70186# a_18162_70226# a_39246_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6408 a_42658_59504# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6409 a_38546_14878# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X641 VSS a_27603_34191# a_30857_39425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6410 a_27049_35515# a_26552_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X6411 a_47678_7452# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6412 a_43566_7850# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6413 a_27502_59182# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6414 VDD a_12934_35823# a_16147_36911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6415 a_6403_37252# a_6061_38377# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6416 VSS a_42024_46805# a_41968_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6417 a_21082_61150# pmat.row_n[5] a_21574_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6418 a_2215_15823# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6419 VSS pmat.row_n[1] a_31518_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X642 a_46182_23954# pmat.row_n[15] a_46674_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6420 a_25098_16926# pmat.row_n[8] a_25590_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6421 VDD a_6664_26159# a_19439_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6422 VDD a_32871_49007# a_9411_2215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X6423 a_8653_12925# a_8175_12533# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6424 a_19470_7850# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6425 VSS a_46263_52245# pmat.col[27] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6426 VSS a_10391_62911# a_10325_62985# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6427 a_32218_66170# a_18546_66212# a_32126_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6428 VDD a_9869_62581# a_9759_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6429 VDD a_12353_16609# a_12243_16733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X643 nmat.col[7] ANTENNA__1190__B1.DIODE a_14471_4943# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X6430 a_9831_74183# a_10515_75895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6431 VDD nmat.rowon_n[4] a_32126_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6432 VSS VDD a_29510_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6433 a_45673_31599# a_38851_28327# a_45589_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X6434 a_7167_52105# a_6817_51733# a_7072_52093# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X6435 a_4583_68021# a_7674_69135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X6436 VSS a_13091_52047# a_20316_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6437 vcm a_18162_68218# a_19166_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6438 VDD a_25681_28879# a_26355_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6439 a_41162_8894# a_18162_8488# a_41254_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X644 a_46182_19938# a_18162_19532# a_46274_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6440 vcm a_18162_63198# a_20170_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6441 VSS a_8735_54207# a_8669_54281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6442 VSS pmat.row_n[15] a_50594_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6443 VSS a_37471_49551# _1154_.A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X6444 a_20078_67174# pmat.row_n[11] a_20570_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6445 VSS a_21371_50087# a_24775_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X6446 vcm a_18162_18528# a_37238_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6447 a_41254_16520# a_18546_16518# a_41162_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6448 a_50198_56130# pmat.row_n[0] a_50690_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6449 a_19166_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X645 a_50198_72194# VDD a_50690_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6450 VDD a_1957_43567# a_14792_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6451 VSS config_1_in[2] a_1591_11471# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6452 vcm a_18162_62194# a_33222_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6453 VSS a_2411_16101# a_2369_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6454 VSS a_2046_30184# a_2787_33237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6455 a_51294_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6456 a_33130_66170# pmat.row_n[10] a_33622_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6457 a_36538_17890# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6458 a_15439_48071# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6459 VSS pmat.row_n[7] a_40554_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X646 a_4337_41935# a_4253_42729# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=0p ps=0u w=840000u l=150000u
X6460 VDD a_7527_30676# a_7047_31226# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X6461 a_18162_66210# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X6462 a_9759_70045# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X6463 a_5331_53511# a_4259_31375# a_5505_53387# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6464 a_20474_22910# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6465 a_3978_48071# a_3987_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6466 VDD a_1674_57711# a_11711_58261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6467 a_12703_31055# a_12079_31061# a_12595_31433# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X6468 a_33382_46983# a_32687_46607# a_33519_46831# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X6469 a_38552_32521# a_37637_32149# a_38205_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X647 a_30210_7484# a_18546_7482# a_30118_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6470 a_7013_34863# a_5823_34863# a_6904_34863# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6471 a_45574_72234# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6472 VDD VDD a_32126_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6473 a_27198_17524# a_18546_17522# a_27106_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6474 a_41162_58138# pmat.row_n[2] a_41654_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6475 a_10878_58487# a_11711_56079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6476 a_30219_29967# a_29968_30083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X6477 a_41558_11866# nmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6478 a_21478_9858# nmat.rowon_n[14] a_21082_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6479 VSS a_11927_27399# a_11987_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.565e+11p ps=5.92e+06u w=650000u l=150000u
X648 a_50690_21508# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6480 a_20811_39095# a_19689_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X6481 a_24490_21906# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6482 VSS a_42240_29423# a_43351_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6483 a_35224_50613# _1154_.X a_35447_50959# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X6484 a_1644_74549# a_1823_74557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6485 VDD config_1_in[5] a_1591_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X6486 a_27106_57134# pmat.row_n[1] a_27598_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6487 a_36234_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6488 a_38546_55166# VSS a_38150_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6489 VDD a_40105_47375# a_47035_43817# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X649 a_49686_65528# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6490 a_31614_55488# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6491 VSS VDD a_22482_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6492 a_14471_27247# a_12987_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u
X6493 vcm a_18162_23548# a_32218_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6494 VSS a_19689_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X6495 a_10117_54697# a_9213_53903# a_10045_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X6496 vcm a_18162_13508# a_28202_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6497 a_7527_30676# a_7619_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6498 a_49286_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6499 a_2319_61493# a_2163_61761# a_2464_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X65 a_12175_55535# a_10497_54697# a_12038_55687# VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X650 a_50290_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6500 a_8175_12533# a_8378_12691# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6501 a_32218_11500# a_18546_11498# a_32126_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6502 VSS a_4443_27247# a_4339_27804# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X6503 VSS a_12345_36924# a_22043_35041# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6504 VDD VSS a_40158_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6505 a_11275_40214# a_11093_40214# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6506 a_27502_12870# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6507 a_39550_63198# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6508 VSS a_5320_27023# a_6406_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6509 VSS pmat.row_n[2] a_31518_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X651 VSS a_7436_60039# a_6816_60699# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6510 a_5941_13103# a_5173_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6511 VDD a_26889_47073# a_26779_47197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6512 a_13547_48169# a_13462_48071# a_13329_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6513 a_17927_48437# a_17397_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X6514 VDD a_1781_9308# a_1725_11254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6515 a_10223_26703# a_9779_26819# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6516 a_5455_72719# a_5363_73807# a_5361_72719# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X6517 VSS pmat.sample_n a_18162_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X6518 VDD a_19584_52423# a_21647_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6519 a_30118_7890# a_18162_7484# a_30210_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X652 a_26364_40517# a_25301_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6520 a_47298_29673# a_37291_29397# a_47212_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X6521 a_2203_39049# a_1757_38677# a_2107_39049# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X6522 a_6017_6575# a_5654_9527# a_5935_6575# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6523 vcm.sky130_fd_sc_hd__nand2_1_0.Y vcm.sky130_fd_sc_hd__buf_4_3.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6524 a_44266_70186# a_18546_70228# a_44174_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6525 a_37146_22950# pmat.row_n[14] a_37638_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6526 a_2215_36495# a_1591_36501# a_2107_36873# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X6527 a_36234_9492# a_18546_9490# a_36142_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6528 a_41654_20504# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6529 VDD pmat.rowoff_n[15] a_44174_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X653 a_6971_70589# a_5687_71829# a_6608_70455# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6530 nmat.col_n[27] a_17139_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6531 a_22039_36950# a_21857_36950# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6532 a_41254_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6533 VDD a_3746_58487# a_9217_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6534 a_44174_64162# a_18162_64202# a_44266_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6535 VDD a_7263_42453# a_4128_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6536 a_13437_26703# a_9217_23983# a_13319_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=3.04e+06u as=4.4e+11p ps=2.88e+06u w=1e+06u l=150000u
X6537 a_37519_46983# a_37791_46811# a_37749_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6538 a_13917_72373# a_13699_72777# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X6539 VSS pmat.row_n[6] a_29510_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X654 VDD a_14887_46377# a_34768_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X6540 a_14641_57711# a_14287_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6541 a_31214_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6542 a_33526_60186# pmat.rowon_n[4] a_33130_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6543 VDD pmat.rowoff_n[7] a_34134_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6544 a_7847_24233# a_6173_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X6545 a_33526_19898# nmat.rowon_n[4] a_33130_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6546 VDD a_7079_34837# a_7066_35229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6547 a_24737_30485# a_23933_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X6548 a_4265_40303# a_3659_39733# a_4193_40303# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6549 vcm a_18162_9492# a_34226_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X655 VSS a_12993_66415# a_14289_66421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6550 a_45178_70186# pmat.row_n[14] a_45670_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6551 VDD nmat.rowon_n[9] a_47186_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6552 result_out[2] a_1644_56053# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6553 a_45270_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6554 a_42166_12910# a_18162_12504# a_42258_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6555 a_6128_59887# a_5497_62839# a_6037_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6556 a_45325_38127# a_45047_38155# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6557 a_21174_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6558 VSS pmat.row_n[13] a_42562_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6559 a_25505_32143# a_23933_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.25e+11p pd=2.65e+06u as=0p ps=0u w=1e+06u l=150000u
X656 a_22178_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6560 a_34226_58138# a_18546_58180# a_34134_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6561 VDD a_9411_2215# a_28543_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X6562 a_31596_34191# a_31419_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6563 a_21478_71230# pmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6564 VSS a_45019_38645# a_45589_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6565 a_29233_47741# a_29189_47349# a_29067_47753# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6566 a_7431_11837# a_7283_11484# a_7068_11703# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6567 a_35630_11468# nmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6568 VSS a_1858_25615# a_12857_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6569 a_11545_18517# a_4383_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X657 a_13013_27023# a_13145_26935# VSS VSS sky130_fd_pr__nfet_01v8 ad=6.24e+11p pd=5.82e+06u as=0p ps=0u w=650000u l=150000u
X6570 a_50690_9460# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6571 VSS a_23884_40517# a_23847_40183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X6572 a_39197_38567# a_39505_38780# a_22153_37179# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X6573 VDD a_16966_29673# nmat.en_bit_n[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X6574 a_18162_17524# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X6575 a_22578_70548# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6576 vcm a_18162_10496# a_31214_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6577 a_39246_21540# a_18546_21538# a_39154_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6578 VSS ANTENNA__1184__B1.DIODE a_40317_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6579 a_25325_29125# a_23933_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X658 a_49194_55126# a_18162_55166# a_49286_55126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6580 a_40771_50959# a_24867_53135# pmat.col[21] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6581 a_48682_10464# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6582 a_3763_6409# a_3247_6037# a_3668_6397# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X6583 a_25190_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6584 a_22086_60146# a_18162_60186# a_22178_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6585 VSS a_1923_31743# a_3320_30333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6586 VSS pmat.row_n[12] a_46578_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6587 a_43566_65206# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6588 a_32218_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6589 VDD a_1957_43567# a_10795_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 a_39550_24918# VSS a_39154_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6590 VSS a_40105_47375# a_46684_43343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X6591 VSS a_30641_44743# a_32035_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X6592 VSS a_4259_31375# a_6925_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X6593 VSS a_35559_30209# a_35520_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6594 a_19074_13914# a_18162_13508# a_19166_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6595 VDD nmat.rowon_n[13] a_25098_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6596 VSS a_7415_29397# a_19611_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6597 a_40554_58178# pmat.rowon_n[2] a_40158_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6598 a_13718_68591# a_13279_68841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X6599 a_39154_63158# pmat.row_n[7] a_39646_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X66 a_4445_64239# a_2879_57487# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X660 clk_dig a_25667_35253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6600 VDD a_25681_28879# a_27605_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6601 a_25839_49783# a_30687_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6602 a_23486_68218# pmat.rowon_n[12] a_23090_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6603 VSS pmat.row_n[3] a_49590_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6604 a_3325_36495# a_2847_36799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6605 a_43662_61512# pmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6606 vcm a_18162_16520# a_30210_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6607 a_33222_19532# a_18546_19530# a_33130_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6608 a_51294_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6609 a_47678_16488# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X661 a_35534_60186# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6610 a_37238_69182# a_18546_69224# a_37146_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6611 a_14533_39631# a_14107_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6612 VDD a_6611_57399# a_6559_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X6613 a_36234_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6614 a_5357_62779# a_6583_61519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X6615 VSS nmat.sample_n a_18162_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X6616 VDD a_4043_22869# a_2835_13077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X6617 a_1757_50095# a_1591_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6618 a_4075_50087# a_4167_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X6619 a_33607_31599# a_29163_29423# a_33501_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X662 a_36142_15922# pmat.row_n[7] a_36634_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6620 a_3641_59709# a_3262_59343# a_3569_59709# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6621 VDD a_44774_40821# a_45164_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X6622 a_14558_24233# a_13768_22325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6623 a_35382_34191# a_35205_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6624 a_2785_38127# a_2743_38279# a_2283_39189# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X6625 a_34828_40517# a_33765_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6626 a_1644_64213# a_1823_64213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6627 a_3203_25398# a_2952_25045# a_2744_25223# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6628 VDD pmat.rowon_n[10] a_19074_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6629 a_26498_59182# pmat.rowon_n[3] a_26102_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X663 VSS pmat.row_n[13] a_36538_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6630 VDD pmat.rowon_n[5] a_20078_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6631 a_5897_38127# a_4533_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X6632 VSS a_33423_47695# a_45201_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6633 vcm a_18162_65206# a_38242_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6634 a_2951_11471# a_2327_11477# a_2843_11849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6635 a_34134_9898# a_18162_9492# a_34226_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6636 a_38150_69182# pmat.row_n[13] a_38642_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6637 a_42258_63158# a_18546_63200# a_42166_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6638 a_4553_18297# a_3576_17143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6639 a_42658_67536# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X664 a_35534_19898# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6640 a_46934_52047# ANTENNA__1395__B1.DIODE a_46765_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X6641 a_42166_57134# a_18162_57174# a_42258_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6642 a_6568_59887# a_5939_60137# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6643 a_12311_54135# a_12003_52815# a_12709_54223# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X6644 VDD a_14011_19087# a_10515_61839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X6645 a_25098_67174# a_18162_67214# a_25190_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6646 VDD pmat.rowon_n[4] a_24094_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6647 VSS VDD a_27502_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6648 a_44879_46070# a_44628_45717# a_44420_45895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X6649 a_46522_34293# a_32405_32463# a_46779_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X665 a_2419_53351# a_3707_53903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6650 VDD a_9583_10121# a_11731_8751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6651 a_37680_41831# a_11113_40835# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6652 VSS pmat.row_n[14] a_42562_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6653 a_39246_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6654 a_6661_29199# a_4068_25615# a_6579_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6655 a_7027_29673# a_6981_28879# a_7109_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X6656 a_8333_24847# a_8307_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6657 VDD a_26460_40517# a_26364_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6658 a_10216_69679# a_9135_69679# a_9869_69921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X6659 a_11545_18517# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X666 VSS a_3615_71631# a_13102_71631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6660 a_35534_17890# nmat.rowon_n[6] a_35138_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6661 VDD a_14287_28995# a_14466_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6662 VSS a_11837_68591# a_13279_68841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6663 VSS a_34002_44527# a_34547_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6664 a_32218_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6665 a_49590_24918# VSS a_49194_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6666 a_30687_48071# a_29076_48695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X6667 a_46182_15922# pmat.row_n[7] a_46674_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6668 a_39550_7850# VDD a_39154_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6669 VSS pmat.row_n[13] a_46578_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X667 a_40650_13476# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6670 a_51598_7850# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X6671 a_41254_24552# a_18546_24550# a_41162_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6672 a_50690_13476# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6673 a_40250_66170# a_18546_66212# a_40158_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6674 a_25423_32463# a_11067_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=0p ps=0u w=650000u l=150000u
X6675 vcm a_18162_70226# a_33222_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6676 a_49686_57496# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6677 a_37238_14512# a_18546_14510# a_37146_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6678 VDD a_3891_25623# a_4068_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6679 a_19746_28111# a_20310_28029# a_20164_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X668 a_2012_18365# a_1895_18170# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6680 a_36234_56130# a_18546_56172# a_36142_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6681 VDD vcm.sky130_fd_sc_hd__nand2_1_1.A a_77980_40594# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6682 a_45829_35407# a_45475_35520# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6683 a_19074_58138# a_18162_58178# a_19166_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6684 a_16911_52423# a_17183_52251# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6685 VSS pmat.row_n[1] a_44570_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6686 a_30118_20942# pmat.row_n[12] a_30610_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6687 a_33622_23516# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6688 a_24602_47919# a_19541_28879# a_24602_48169# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X6689 a_33222_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X669 vcm a_18162_70226# a_23182_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6690 VSS a_8305_20871# a_7847_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.565e+11p ps=5.92e+06u w=650000u l=150000u
X6691 a_16478_29423# a_16131_29429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X6692 a_12163_62723# a_12076_62839# a_12081_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6693 a_2603_58368# a_2727_58470# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6694 a_30118_16926# a_18162_16520# a_30210_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6695 VDD pmat.rowon_n[2] a_40158_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6696 a_39550_16886# nmat.rowon_n[7] a_39154_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6697 VSS pmat.row_n[5] a_36538_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6698 VDD a_19834_34191# a_20711_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6699 a_40554_11866# nmat.rowon_n[12] a_40158_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X67 a_43662_17492# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X670 VSS pmat.row_n[10] a_25494_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6700 a_83094_10089# ANTENNA__1184__B1.DIODE a_82788_9991# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X6701 a_10227_60751# a_10190_60663# a_10058_60431# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6702 a_19074_17930# pmat.row_n[9] a_19566_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6703 VSS pmat.row_n[15] a_19470_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6704 VSS a_39321_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X6705 a_39472_48841# a_38557_48469# a_39125_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X6706 a_23582_15484# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6707 VSS pmat.row_n[4] a_49590_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6708 a_20078_12910# pmat.row_n[4] a_20570_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6709 a_23486_21906# nmat.rowon_n[2] a_23090_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X671 a_39646_57496# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6710 VSS cgen.dlycontrol4_in[3] a_33395_43455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6711 vcm a_18162_62194# a_41254_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6712 VDD pmat.rowon_n[1] a_26102_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6713 a_17317_31849# pmat.rowon_n[7] nmat.rowon_n[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X6714 a_10245_51335# a_9995_52299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6715 a_41162_66170# pmat.row_n[10] a_41654_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6716 VDD a_20164_27791# a_20616_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X6717 a_34134_15922# a_18162_15516# a_34226_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6718 a_6623_22057# a_2683_22089# a_6551_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6719 a_46684_43343# a_7109_29423# a_46013_42997# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X672 a_22199_49667# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X6720 a_26498_12870# pmat.rowoff_n[4] a_26102_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6721 a_38546_63198# pmat.rowon_n[7] a_38150_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6722 a_24094_11906# pmat.row_n[3] a_24586_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6723 a_10845_12559# a_10443_12879# a_10681_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X6724 VSS a_41731_49525# a_45405_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6725 a_35230_17524# a_18546_17522# a_35138_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6726 vcm a_18162_21540# a_28202_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6727 VDD a_11711_56079# a_10878_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6728 a_13459_4943# _1187_.A2 nmat.col[10] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6729 a_2250_74397# a_2124_74299# a_1846_74283# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X673 a_9655_6335# a_9480_6409# a_9834_6397# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6730 a_31214_61150# a_18546_61192# a_31122_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6731 vcm a_18162_68218# a_40250_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6732 a_35534_68218# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6733 VDD nmat.rowon_n[1] a_36142_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6734 a_9089_64061# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6735 VDD a_11807_51157# a_4991_69831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X6736 a_3609_9295# a_3415_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6737 nmat.col[8] a_10883_3303# a_27618_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X6738 a_23486_8854# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6739 a_27598_8456# nmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X674 a_15749_28111# a_13479_26935# a_15667_28111# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6740 a_11902_56775# a_12311_54135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6741 vcm a_18162_13508# a_36234_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6742 a_40250_11500# a_18546_11498# a_40158_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6743 VSS pmat.row_n[15] a_43566_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6744 a_13529_34951# a_13801_34427# a_14923_34473# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X6745 a_3431_39759# a_2935_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X6746 vcm a_18162_12504# a_49286_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6747 a_32126_61150# pmat.row_n[5] a_32618_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6748 a_41254_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6749 VSS a_16635_31573# a_4707_32156# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X675 VDD VSS a_43170_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6750 a_40250_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6751 VDD a_21981_34191# a_25647_38695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6752 a_37238_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6753 a_33309_42693# a_33617_42333# a_33283_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X6754 a_14471_29673# a_12461_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6755 VDD a_4443_27247# a_4339_27804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X6756 a_23090_19938# pmat.row_n[11] a_23582_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6757 a_8653_64061# a_8175_63669# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6758 a_44266_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6759 inn_analog clk_ena ctopn VDD sky130_fd_pr__pfet_01v8 ad=1.102e+12p pd=8.76e+06u as=0p ps=0u w=1.9e+06u l=220000u M=4
X676 a_49194_14918# pmat.row_n[6] a_49686_14480# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6760 a_6523_42479# a_6173_42479# a_6428_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X6761 VDD a_37820_30485# a_41335_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6762 a_25590_56492# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6763 a_8782_12559# a_8695_12801# a_8378_12691# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6764 a_27198_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6765 a_20474_71230# pmat.rowon_n[15] a_20078_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6766 a_30210_22544# a_18546_22542# a_30118_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6767 VSS a_1957_43567# a_13685_55357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6768 a_11711_60751# a_10049_60663# a_12155_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6769 a_26194_12504# a_18546_12502# a_26102_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X677 VSS pmat.row_n[12] a_49590_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6770 a_1586_18231# a_3944_28853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6771 VDD a_2791_57703# a_2603_58368# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6772 VDD a_14653_53458# a_14655_53359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6773 a_42166_20942# a_18162_20536# a_42258_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6774 a_45270_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6775 a_25209_42043# a_23700_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X6776 VSS a_1923_61759# a_1881_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6777 VDD a_78165_40202# a_77978_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6778 VSS a_39359_49172# a_38695_48634# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6779 vcm a_18162_18528# a_48282_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X678 a_20078_20942# pmat.row_n[12] a_20570_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6780 a_6664_26159# a_7072_26311# a_6323_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6781 a_4312_74005# a_4697_74005# a_4441_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X6782 a_9749_19061# a_8305_20871# a_10129_19203# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6783 a_37737_50095# a_26891_28327# a_34942_51701# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6784 VDD a_7419_14379# a_7377_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6785 a_25384_48169# a_15899_47939# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X6786 a_4745_45519# a_4700_44655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X6787 a_13655_26703# a_13437_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X6788 a_12445_58229# a_12227_58633# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6789 a_24490_70226# pmat.rowon_n[14] a_24094_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X679 a_23582_23516# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6790 a_47582_17890# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6791 a_2163_31741# a_2046_30184# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6792 a_12252_55785# a_10955_55687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X6793 VSS a_13091_52047# a_17459_49641# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6794 a_38242_71190# a_18546_71232# a_38150_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6795 VSS pmat.row_n[7] a_51598_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6796 a_39472_48841# a_38391_48469# a_39125_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6797 VDD a_9871_48463# a_6787_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X6798 vcm a_18162_8488# a_48282_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6799 a_19417_43990# a_19689_44581# a_20811_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X68 a_43566_23914# pmat.rowoff_n[15] a_43170_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X680 a_14336_48071# a_14486_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6800 a_12131_71829# a_12249_71311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X6801 VDD a_46811_33927# a_45908_33749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6802 a_18176_42693# a_18272_42693# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6803 a_6325_77295# a_6281_77537# a_6159_77295# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6804 a_11193_42390# a_11021_42619# a_10979_42390# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X6805 a_28110_21946# a_18162_21540# a_28202_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6806 VDD pmat.rowon_n[7] a_38150_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6807 vcm.sky130_fd_sc_hd__buf_4_1.X a_77980_40594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6808 VSS a_15899_47939# a_24602_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6809 a_42240_29423# a_41703_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X681 a_23182_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6810 a_11209_17782# a_9528_20407# a_10995_17782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X6811 a_27502_61190# pmat.rowon_n[5] a_27106_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6812 VSS pmat.row_n[9] a_24490_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6813 VDD a_3339_70759# a_7605_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6814 a_9943_15645# a_9319_15279# a_9835_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6815 VSS a_3325_36495# a_4073_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X6816 a_47591_51183# _1194_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6817 a_49194_10902# a_18162_10496# a_49286_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6818 VSS a_19689_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X6819 a_39154_71190# pmat.row_n[15] a_39646_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X682 a_44266_23548# a_18546_23546# a_44174_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6820 VDD a_5935_6575# a_6337_6825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6821 a_18272_42693# a_17113_42405# a_18235_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X6822 VDD a_1957_43567# a_13739_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6823 a_35534_21906# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6824 vcm a_18162_24552# a_30210_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6825 a_4951_76983# a_5047_76983# a_5349_77071# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X6826 a_40250_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6827 a_10471_12791# a_10839_11989# a_10785_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6828 a_47278_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6829 a_28202_59142# a_18546_59184# a_28110_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X683 a_20078_16926# a_18162_16520# a_20170_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6830 vcm a_18162_56170# a_25190_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6831 VSS pmat.row_n[8] a_28506_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6832 a_25494_13874# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6833 a_32522_14878# nmat.rowon_n[9] a_32126_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6834 a_2080_70045# a_1643_69653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6835 a_26194_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6836 a_19143_41085# a_18963_41085# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6837 a_37238_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6838 VDD VSS a_51202_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6839 a_2847_63999# a_2672_64073# a_3026_64061# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X684 _1183_.A2 a_47357_38127# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X6840 a_38714_32143# a_37637_32149# a_38552_32521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6841 VSS a_8693_11769# a_8627_11837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6842 a_9552_67191# a_9545_66567# a_9783_67075# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6843 a_17191_48981# a_17139_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X6844 a_37542_66210# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6845 a_2526_13647# a_2400_13763# a_2122_13779# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6846 a_2012_26159# a_1895_26372# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6847 vcm a_18162_55166# a_29206_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6848 a_27579_34967# a_27687_34967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6849 a_44570_67214# pmat.rowon_n[11] a_44174_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X685 VDD pmat.rowon_n[9] a_26102_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6850 VSS pmat.row_n[8] a_41558_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6851 a_9642_6031# a_8565_6037# a_9480_6409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6852 cgen.dlycontrol4_in[5] a_1591_23983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6853 a_29114_59142# pmat.row_n[3] a_29606_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6854 vcm a_18162_15516# a_51294_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6855 a_27421_41814# a_26773_40955# a_27895_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X6856 a_33222_8488# a_18546_8486# a_33130_8894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6857 VSS a_4312_74005# a_4048_74549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X6858 a_10400_15279# a_9319_15279# a_10053_15521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X6859 a_26283_42325# a_26459_42657# a_26411_42717# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X686 a_5904_55311# a_4351_55527# a_5329_54965# VSS sky130_fd_pr__nfet_01v8 ad=1.6575e+11p pd=1.81e+06u as=5.72e+11p ps=4.36e+06u w=650000u l=150000u
X6860 a_42166_65166# a_18162_65206# a_42258_65166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6861 a_2969_55785# a_1591_54991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X6862 a_48190_22950# pmat.row_n[14] a_48682_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6863 a_38150_55126# a_18162_55166# a_38242_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6864 a_7445_29673# a_2952_25045# a_7803_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X6865 a_34530_59182# pmat.rowon_n[3] a_34134_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6866 a_7186_25615# a_6747_25731# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X6867 VSS a_43971_28487# a_27763_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6868 VSS pmat.row_n[7] a_27502_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6869 VSS a_13479_26935# a_14751_28341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X687 VSS a_4383_7093# a_11216_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6870 a_11138_50347# a_11416_50363# a_11372_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6871 a_9913_62973# a_9869_62581# a_9747_62985# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6872 vcm a_18162_17524# a_24186_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6873 a_38150_14918# pmat.row_n[6] a_38642_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6874 a_39939_29967# a_39666_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6875 a_39154_18934# a_18162_18528# a_39246_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6876 VDD pmat.rowoff_n[7] a_45178_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6877 a_42658_12472# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6878 nmat.col_n[30] a_84028_9615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X6879 a_40592_31599# a_39939_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X688 a_51202_13914# a_18162_13508# a_51294_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6880 a_40158_13914# a_18162_13508# a_40250_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6881 VSS a_10195_30186# a_9899_30724# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6882 a_25755_38695# cgen.dlycontrol3_in[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6883 a_18487_50069# a_18823_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X6884 VSS pmat.en_bit_n[2] a_35534_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6885 a_9466_65149# a_1923_61759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6886 a_32218_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6887 a_3675_15113# a_3229_14741# a_3579_15113# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X6888 a_46182_66170# a_18162_66210# a_46274_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6889 a_18546_60188# pmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X689 VDD a_2563_34837# a_4785_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6890 a_13688_47893# a_12044_49641# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X6891 a_17927_47349# a_18083_47593# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X6892 a_32522_71230# pmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6893 a_36234_64162# a_18546_64204# a_36142_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6894 a_46674_11468# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6895 a_24719_35253# a_24895_35253# a_24847_35279# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X6896 a_36634_68540# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6897 a_30118_24958# a_18162_24552# a_30210_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6898 VDD ANTENNA__1187__B1.DIODE pmat.col_n[20] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X6899 VSS ANTENNA__1190__B1.DIODE nmat.col[7] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X69 a_40158_14918# pmat.row_n[6] a_40650_14480# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X690 a_30210_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6900 a_29606_21508# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6901 VDD pmat.rowon_n[10] a_40158_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6902 a_29206_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6903 a_40250_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6904 VSS a_14071_74879# a_14005_74953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6905 a_33130_60146# a_18162_60186# a_33222_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6906 a_25802_48169# a_19541_28879# a_25384_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X6907 a_23182_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6908 a_16833_51183# a_13091_52047# a_16761_51183# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6909 a_19566_13476# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X691 a_21739_29415# a_43659_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6910 VDD a_10216_69679# a_10391_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6911 vcm a_18162_70226# a_41254_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6912 VDD nmat.rowon_n[12] a_23090_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6913 vcm a_18162_60186# a_37238_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6914 a_20752_36165# a_19689_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6915 VDD a_1586_63927# a_12723_64789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6916 a_14158_65149# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6917 a_3325_40847# a_2847_41151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6918 a_37146_64162# pmat.row_n[8] a_37638_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6919 a_34134_23954# a_18162_23548# a_34226_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X692 a_13553_50461# a_13290_50095# a_13140_50247# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6920 a_12383_39631# a_12235_39913# a_12020_39783# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6921 VDD pmat.rowon_n[9] a_44174_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6922 a_41654_62516# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6923 VDD a_3868_33609# a_4043_33535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6924 a_24765_28111# a_13091_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6925 VDD a_18563_27791# a_37795_29111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6926 a_51598_58178# pmat.rowon_n[2] a_51202_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6927 a_23663_43177# a_22541_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6928 a_26498_62194# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6929 VSS pmat.row_n[4] a_30514_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X693 a_26194_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6930 a_6417_49007# a_6373_49249# a_6251_49007# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6931 VSS pmat.row_n[11] a_30514_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6932 VDD pmat.rowon_n[1] a_34134_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6933 a_44570_20902# pmat.rowoff_n[12] a_44174_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6934 a_13814_59663# a_9963_13967# a_13645_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6935 vcm a_18162_71230# a_27198_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6936 VDD nmat.rowon_n[14] a_21082_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6937 a_2325_17973# a_2107_18377# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X6938 VDD pmat.rowon_n[0] a_47186_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6939 VSS a_22522_50247# a_22475_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X694 VSS pmat.row_n[4] a_39550_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6940 vcm a_18162_58178# a_31214_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6941 a_27598_63520# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6942 a_5233_40553# a_4705_39759# a_5161_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6943 a_40967_30511# a_28704_29568# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6944 VDD pmat.rowon_n[5] a_31122_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6945 a_34530_12870# pmat.rowoff_n[4] a_34134_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6946 a_46968_45743# a_47147_44655# a_46797_45993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6947 VSS a_28116_37479# a_28079_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X6948 a_9182_7119# a_8105_7125# a_9020_7497# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6949 a_40158_58138# a_18162_58178# a_40250_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X695 VSS a_12345_36924# a_12289_36950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6950 vcm a_18162_21540# a_36234_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6951 VSS a_7693_22365# a_12212_22467# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6952 a_3944_28853# clk_dig VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6953 VSS a_45405_30511# ANTENNA__1183__B1.DIODE VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.64e+11p ps=3.72e+06u w=650000u l=150000u M=4
X6954 a_23090_68178# a_18162_68218# a_23182_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6955 a_34002_34191# a_33825_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6956 vcm a_18162_20536# a_49286_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6957 a_82787_54421# _1154_.A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6958 a_40158_17930# pmat.row_n[9] a_40650_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6959 a_37238_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X696 a_26649_34219# a_26583_34343# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6960 VSS a_12020_39783# a_11565_39061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6961 VDD nmat.rowon_n[15] a_37146_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6962 a_44697_48783# a_44774_48695# a_45152_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6963 a_23847_38007# a_23329_37462# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X6964 a_44423_36815# a_44811_36469# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6965 a_2559_46261# a_2347_46070# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6966 VSS a_5081_53135# a_6242_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6967 VSS a_23395_53135# a_43347_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X6968 a_43566_8854# nmat.rowon_n[15] a_43170_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6969 a_32371_47349# a_30999_48071# a_32589_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X697 a_2617_35113# a_2563_34837# a_1770_35015# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6970 VSS pmat.row_n[12] a_20474_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6971 a_46578_59182# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6972 a_26194_20536# a_18546_20534# a_26102_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6973 a_8565_6037# a_8399_6037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6974 VDD a_9427_50095# a_10299_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6975 a_32035_38007# a_30913_38053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6976 VSS pmat.row_n[1] a_50594_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6977 VSS a_9581_56079# a_12353_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X6978 a_46578_17890# nmat.rowon_n[6] a_46182_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6979 a_44174_16926# pmat.row_n[8] a_44666_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X698 result_out[10] a_1644_68565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6980 a_19470_8854# nmat.rowon_n[15] a_19074_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6981 a_29510_69222# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6982 VDD a_2935_38279# a_2893_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6983 a_31518_8854# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6984 VSS pmat.row_n[11] a_33526_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6985 a_30514_64202# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6986 VSS pmat.rowon_n[7] pmat.rowoff_n[10] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6987 VDD a_22787_34709# a_12197_38306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6988 a_6553_53047# a_5566_44905# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.1275e+11p pd=3.87e+06u as=0p ps=0u w=650000u l=150000u
X6989 VSS a_7037_70521# a_6971_70589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X699 a_8765_64757# a_8547_65161# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X6990 a_46949_28585# a_38851_28327# a_46863_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X6991 a_4699_28701# a_4075_28335# a_4591_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X6992 a_7644_16341# a_10575_15253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6993 a_13686_13967# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6994 nmat.col[19] _1154_.X a_83630_3311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X6995 a_51294_66170# a_18546_66212# a_51202_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6996 a_35230_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6997 a_47278_56130# a_18546_56172# a_47186_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6998 VSS pmat.row_n[3] a_23486_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6999 a_20474_56170# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7 a_12531_34743# a_11409_34789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=3.13473e+15p ps=2.99317e+10u w=800000u l=150000u
X70 a_6574_5853# a_6487_5629# a_6170_5739# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X700 VDD a_25815_43957# a_25639_43957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7000 a_44976_47349# a_33467_46261# a_45368_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X7001 VDD pmat.rowon_n[2] a_51202_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7002 VSS pmat.row_n[5] a_47582_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7003 a_21574_16488# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7004 a_17635_39605# a_17811_39605# a_17763_39631# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X7005 a_6800_69251# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7006 a_14125_13647# a_11435_58791# pmat.rowon_n[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7007 a_51598_11866# nmat.rowon_n[12] a_51202_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7008 VDD pmat.rowon_n[15] a_38150_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7009 a_23788_40517# a_23884_40517# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X701 a_43566_10862# nmat.rowon_n[13] a_43170_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7010 a_9861_26819# a_9777_26935# a_9779_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7011 a_9779_26819# a_9777_26935# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X7012 VSS a_11921_41814# a_10985_42044# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X7013 a_34626_15484# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7014 VSS pmat.sw ANTENNA_fanout52_A.DIODE VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X7015 a_2200_10927# a_1761_9839# a_1979_11254# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7016 VSS a_10959_23983# a_12449_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7017 a_38242_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7018 ANTENNA__1184__B1.DIODE a_47212_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u M=4
X7019 VSS a_1717_13647# a_6879_10473# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X702 a_24591_28327# a_40567_32403# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7020 a_5510_14013# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7021 a_35007_44527# a_34830_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7022 a_24490_55166# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7023 a_11067_30287# a_21279_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7024 a_1644_56053# a_1591_56623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7025 pmat.col_n[29] ANTENNA__1196__A2.DIODE a_46027_52047# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7026 a_6428_42479# a_6311_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7027 a_36142_21946# a_18162_21540# a_36234_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7028 a_5537_22057# a_3351_27249# a_5455_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7029 a_19689_39141# a_18272_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X703 a_2203_33775# a_1757_33775# a_2107_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X7030 a_11149_40188# a_33255_43777# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X7031 a_28202_67174# a_18546_67216# a_28110_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7032 vcm a_18162_64202# a_25190_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7033 VSS a_7497_11769# a_7431_11837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7034 a_35138_11906# pmat.row_n[3] a_35630_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7035 VDD VDD a_26102_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7036 VSS VDD a_22482_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7037 a_25098_68178# pmat.row_n[12] a_25590_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7038 a_36538_66210# pmat.rowon_n[10] a_36142_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7039 VSS a_23815_50069# pmat.row_n[6] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X704 a_8356_23671# a_2683_22089# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X7040 VDD pmat.rowon_n[13] a_32126_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7041 a_46274_17524# a_18546_17522# a_46182_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7042 VDD pmat.rowon_n[3] a_28110_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7043 cgen.dlycontrol3_in[2] a_1591_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7044 VSS a_36380_34191# a_36486_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7045 VDD a_2659_35015# a_4253_42729# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7046 VSS a_1586_8439# a_7939_7125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7047 a_46182_57134# pmat.row_n[1] a_46674_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7048 vcm a_18162_63198# a_29206_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7049 VSS VDD a_41558_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X705 a_26594_14480# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7050 VDD a_35099_34191# a_35205_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7051 a_4308_21495# a_4516_21531# a_4450_21629# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7052 a_29114_67174# pmat.row_n[11] a_29606_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7053 vcm a_18162_23548# a_51294_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7054 a_35039_29941# a_35242_30099# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7055 VDD a_38205_32117# a_38095_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7056 a_10579_76029# a_10515_75895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7057 a_33622_65528# pmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7058 a_30118_62154# pmat.row_n[6] a_30610_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7059 vcm a_18162_13508# a_47278_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X706 VDD nmat.rowon_n[6] a_29114_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7060 a_20170_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7061 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7062 a_51294_11500# a_18546_11498# a_51202_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7063 a_38150_63158# a_18162_63198# a_38242_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7064 VSS a_9195_58951# a_8193_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7065 a_46578_12870# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7066 VSS pmat.row_n[13] a_20474_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7067 VSS pmat.row_n[2] a_50594_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7068 a_23582_57496# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7069 a_29510_22910# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X707 a_26498_20902# pmat.rowoff_n[12] a_26102_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7070 a_4043_22869# a_2007_25597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X7071 VSS a_15753_28879# a_24524_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7072 vcm a_18162_7484# a_37238_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7073 VSS pmat.row_n[12] a_33526_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7074 VSS a_1923_53055# a_1881_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7075 a_24186_13508# a_18546_13506# a_24094_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7076 a_18546_58180# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7077 a_31518_71230# pmat.rowon_n[15] a_31122_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7078 VDD a_4680_63669# a_3751_64757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7079 a_19487_49159# a_19759_48987# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X708 VDD ANTENNA__1395__A1.DIODE a_45471_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X7080 a_12225_74575# a_11823_74895# a_12061_74895# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X7081 a_47278_7484# a_18546_7482# a_47186_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7082 VDD a_13795_10687# a_13782_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7083 a_10954_73195# a_11232_73211# a_11188_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7084 VSS pmat.row_n[4] a_23486_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7085 VSS pmat.row_n[7] a_35534_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7086 VDD a_22153_37179# a_39197_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7087 a_4241_7663# a_3663_9269# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X7088 VDD a_10781_42364# a_11193_42390# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7089 a_13012_57487# a_6927_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=0p ps=0u w=650000u l=150000u M=2
X709 a_4511_71631# a_2727_58470# a_4415_71631# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X7090 VDD a_43533_30761# a_44647_35520# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7091 a_2467_35925# a_4031_37191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7092 a_34924_37253# a_33765_36965# a_34828_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7093 VSS pmat.row_n[6] a_48586_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7094 a_45574_18894# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7095 a_50290_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7096 VDD _1154_.A a_46886_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7097 a_36234_72194# a_18546_72236# a_36142_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7098 vcm a_18162_9492# a_28202_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7099 VDD a_10400_15279# a_10575_15253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X71 a_41162_18934# a_18162_18528# a_41254_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X710 a_24094_15922# a_18162_15516# a_24186_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7100 a_17969_50755# a_16800_47213# a_17874_50755# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X7101 a_19965_36603# a_17996_36391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X7102 a_49286_71190# a_18546_71232# a_49194_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7103 VDD pmat.rowon_n[8] a_36142_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7104 VSS a_2411_43301# a_2369_43389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7105 a_40250_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7106 VDD VSS a_49194_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7107 a_10873_40693# a_30403_40747# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X7108 VSS a_12437_28879# a_17830_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7109 VDD a_2944_56872# a_2882_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X711 VDD pmat.rowoff_n[4] a_30118_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7110 a_20078_71190# a_18162_71230# a_20170_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7111 a_25494_62194# pmat.rowon_n[6] a_25098_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7112 a_50198_59142# pmat.row_n[3] a_50690_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7113 VSS pmat.row_n[10] a_22482_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7114 a_44666_9460# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7115 a_37146_72194# VDD a_37638_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7116 a_7088_42479# a_6007_42479# a_6741_42721# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X7117 a_10781_75119# a_10697_75218# a_10699_75119# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7118 a_9414_12559# a_8656_12675# a_8851_12533# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7119 a_41654_70548# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X712 vcm a_18162_61190# a_44266_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7120 a_37638_60508# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7121 a_32072_42919# a_30913_43131# a_32035_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7122 a_41162_60146# a_18162_60186# a_41254_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7123 vcm a_18162_57174# a_23182_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7124 a_11711_50959# a_40949_48437# a_40897_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7125 VSS pmat.sample_n a_18162_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X7126 a_51294_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7127 a_24094_70186# a_18162_70226# a_24186_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7128 a_23486_14878# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7129 VSS a_26659_34967# a_12069_36341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X713 a_15048_41605# a_11021_42619# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X7130 a_14097_55369# a_12907_54997# a_13988_55369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X7131 VSS a_9184_51335# a_6979_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7132 VDD nmat.rowon_n[13] a_44174_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7133 VSS a_14839_54599# a_14839_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7134 a_33797_47081# a_33423_47695# a_33382_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7135 a_27598_71552# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7136 VDD a_4737_23957# a_4767_24310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7137 VDD pmat.rowoff_n[12] a_27106_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7138 a_42562_68218# pmat.rowon_n[12] a_42166_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7139 a_8338_20291# a_7644_16341# a_8256_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X714 a_37525_27221# a_24591_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X7140 a_12557_30485# a_6467_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7141 a_27106_61150# a_18162_61190# a_27198_61150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7142 a_48586_66210# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7143 a_25639_43957# a_11041_39860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7144 nmat.rowon_n[7] a_16219_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7145 a_5699_18543# a_5253_18543# a_5603_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X7146 a_18963_41085# a_18975_40871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7147 a_9374_7485# a_2199_13887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7148 a_13102_71311# a_13158_71285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X7149 VDD ANTENNA__1195__A1.DIODE a_42709_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X715 VSS a_3305_17999# a_6651_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7150 a_10455_53387# a_9213_53903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7151 a_35630_63520# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7152 a_46566_52521# _1192_.A2 a_46263_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7153 vcm a_18162_18528# a_22178_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7154 a_11183_35862# a_11001_35862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7155 a_17763_39631# a_12969_40175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7156 a_45574_59182# pmat.rowon_n[3] a_45178_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7157 VSS pmat.row_n[0] a_42562_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7158 a_39646_18496# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7159 a_28202_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X716 _1183_.A2 a_47357_38127# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X7160 a_2215_63695# a_1591_63701# a_2107_64073# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X7161 a_28110_9898# a_18162_9492# a_28202_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7162 a_17900_44007# a_16837_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X7163 VDD nmat.rowon_n[7] a_43170_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7164 a_28506_69222# pmat.rowon_n[13] a_28110_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7165 a_17625_42902# a_17113_41317# a_18235_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7166 VSS a_32411_49559# a_28915_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X7167 vcm a_18162_17524# a_35230_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7168 a_9183_76359# a_6975_76823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X7169 a_21478_17890# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X717 VDD a_46522_34293# a_46912_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X7170 VSS a_2983_48071# a_3983_49911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7171 VSS a_12263_50959# a_18429_51189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X7172 pmat.rowon_n[1] a_14839_54447# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7173 VSS a_4396_69109# a_4340_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7174 VSS a_5331_13951# a_5265_14025# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X7175 a_44174_67174# a_18162_67214# a_44266_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7176 a_49590_58178# pmat.rowon_n[2] a_49194_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7177 VSS VDD a_46578_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7178 a_4712_27023# a_3305_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X7179 VDD a_11067_64015# a_13915_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X718 a_40256_41831# a_40352_41831# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X7180 a_30514_72234# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7181 VSS a_1586_33927# a_1591_40853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7182 VDD a_1586_50247# a_8583_47381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7183 VDD a_6884_74183# a_5931_74183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7184 VSS pmat.row_n[9] a_29510_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7185 VDD a_10391_62911# a_10049_60663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X7186 a_27198_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7187 VSS a_20848_39429# a_20811_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X7188 a_47278_64162# a_18546_64204# a_47186_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7189 a_20848_41605# a_19689_41317# a_20752_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X719 VDD a_10055_31591# a_14747_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X7190 a_40105_47375# a_39647_47679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7191 a_47678_68540# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7192 a_39154_7890# VDD a_39646_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7193 VDD pmat.rowon_n[10] a_51202_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7194 VSS a_6559_6031# a_7206_5853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7195 a_35465_32441# a_7717_14735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7196 VSS pmat.row_n[1] a_19470_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7197 a_21174_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7198 a_23486_55166# VSS a_23090_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7199 a_51294_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X72 VSS a_9785_28879# a_32687_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X720 a_8511_10422# a_8481_10396# a_8439_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7200 a_44984_48783# a_44774_48695# a_44697_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7201 a_49686_7452# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7202 a_45574_7850# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7203 a_12368_35823# a_12191_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7204 VDD pmat.rowon_n[5] a_29114_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7205 a_23844_52271# ANTENNA__1395__A1.DIODE a_23541_52245# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X7206 a_11497_40719# a_11071_41046# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7207 a_34226_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7208 VSS a_43315_48437# a_43261_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7209 a_3687_14735# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X721 a_29225_39659# a_29159_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7210 a_37739_37737# a_36617_37691# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7211 a_8723_67191# a_8491_47911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7212 vcm a_18162_60186# a_48282_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7213 a_48190_64162# pmat.row_n[8] a_48682_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7214 a_24490_63198# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7215 a_13354_2223# a_9411_2215# a_13268_2223# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X7216 VSS a_1586_18231# a_9411_15831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7217 VDD a_44774_48695# a_21279_48999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7218 VSS a_39089_27765# nmat.col[20] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7219 a_34553_42658# a_33489_43131# a_34611_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X722 a_3981_6005# a_3763_6409# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7220 VSS pmat.row_n[15] a_38546_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7221 a_16837_35515# a_16381_35286# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X7222 VSS a_10985_35516# a_10677_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7223 a_42562_21906# nmat.rowon_n[2] a_42166_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7224 vcm a_18162_72234# a_25190_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7225 a_38150_56130# pmat.row_n[0] a_38642_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7226 a_22361_41479# a_22357_43493# a_23420_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7227 a_11807_51157# a_12242_51435# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7228 VDD pmat.rowon_n[1] a_45178_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7229 a_22086_22950# pmat.row_n[14] a_22578_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X723 a_77528_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7230 VSS a_2199_13887# a_7258_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7231 vcm a_18162_22544# a_43262_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7232 VDD pmat.rowon_n[11] a_28110_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7233 VSS a_2099_25236# a_1895_26372# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7234 a_50594_69222# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7235 VDD a_18272_39429# a_18176_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X7236 a_9301_62613# a_9135_62613# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7237 a_28202_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7238 VDD a_47915_46506# nmat.col[31] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7239 a_46848_53135# ANTENNA__1395__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X724 a_19351_28879# a_14365_22351# a_19267_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7240 a_38972_39655# a_37813_39867# a_38876_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7241 a_45574_12870# pmat.rowoff_n[4] a_45178_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7242 VDD a_2419_53351# a_4885_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7243 a_14185_16189# a_11067_16359# a_14103_15936# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7244 VDD a_39125_48437# a_39015_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7245 a_28506_22910# nmat.rowon_n[1] a_28110_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7246 VSS pmat.row_n[14] a_37542_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7247 a_26102_21946# pmat.row_n[13] a_26594_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7248 VDD a_30765_37692# a_30371_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7249 a_11071_41046# a_11113_40835# a_11071_40719# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X725 VDD a_1586_18231# a_2879_19093# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7250 a_30118_70186# pmat.row_n[14] a_30610_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7251 VDD nmat.rowon_n[9] a_32126_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7252 VSS a_6316_8903# a_5654_9527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7253 a_26102_17930# a_18162_17524# a_26194_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7254 vcm a_18162_21540# a_47278_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7255 VDD a_45915_29941# a_22199_30287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X7256 a_46765_36201# a_43776_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X7257 a_10494_77547# a_10811_77437# a_10769_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7258 VSS a_19970_46287# a_20076_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7259 a_30210_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X726 VSS a_12585_37179# a_18235_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X7260 a_43451_30511# a_41227_29423# a_43869_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7261 a_21124_42919# a_19965_43131# a_21087_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7262 a_50290_61150# a_18546_61192# a_50198_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7263 VSS a_2467_46506# a_1987_45370# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7264 a_21279_48999# a_45370_48169# a_45502_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7265 VSS VDD a_30514_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7266 VSS a_25647_34343# a_12345_36924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7267 VDD pmat.rowon_n[2] a_49194_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7268 a_11561_36950# a_10651_37683# a_11347_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X7269 a_49590_11866# nmat.rowon_n[12] a_49194_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X727 a_27106_10902# pmat.row_n[2] a_27598_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7270 a_20570_11468# nmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7271 a_23486_9858# nmat.rowon_n[14] a_23090_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7272 VSS a_6082_46831# a_6553_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7273 a_9112_65161# a_8197_64789# a_8765_64757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X7274 a_19566_55488# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7275 a_19860_30511# a_9307_31068# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7276 VDD a_12895_53359# a_13139_54599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7277 a_29114_12910# pmat.row_n[4] a_29606_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7278 VDD a_3615_71631# a_13102_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7279 a_24186_21540# a_18546_21538# a_24094_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X728 a_42562_58178# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7280 a_42258_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7281 a_33622_10464# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7282 a_2834_17999# a_1757_18005# a_2672_18377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7283 a_18162_61190# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X7284 a_5156_14025# a_4075_13653# a_4809_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7285 VSS pmat.row_n[12] a_31518_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7286 a_51202_61150# pmat.row_n[5] a_51694_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7287 vcm a_18162_69222# a_45270_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7288 VSS pmat.row_n[2] a_19470_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7289 VSS a_9287_77055# a_9221_77129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X729 a_21174_61150# a_18546_61192# a_21082_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7290 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7291 a_42166_19938# pmat.row_n[11] a_42658_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7292 a_28901_48437# a_31152_48071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7293 VSS a_10090_58093# a_9919_57863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7294 a_35646_29967# a_35559_30209# a_35242_30099# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7295 a_15144_36165# a_13985_35877# a_15107_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7296 VSS a_4703_24527# a_9135_22057# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7297 a_22193_48579# a_21279_48999# a_22097_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7298 a_46274_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7299 cgen.dlycontrol4_in[3] a_1591_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X73 a_17900_35303# a_17996_35303# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=8.42088e+14p ps=8.51553e+09u w=420000u l=150000u M=2
X730 VDD pmat.rowon_n[12] a_24094_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7300 a_4075_68583# a_4399_51157# a_4357_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7301 a_2467_46506# a_2559_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7302 a_15899_47939# a_23823_47679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7303 a_24094_63158# pmat.row_n[7] a_24586_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7304 VDD a_37820_30485# a_45719_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7305 a_32126_7890# a_18162_7484# a_32218_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7306 VDD a_20315_29098# nmat.col[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7307 VSS pmat.row_n[3] a_34530_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7308 a_45270_12504# a_18546_12502# a_45178_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7309 VDD VDD a_36142_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X731 a_25494_68218# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7310 a_2893_59709# a_2858_59475# a_2655_59317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7311 a_28110_18934# pmat.row_n[10] a_28602_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7312 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7313 a_22178_69182# a_18546_69224# a_22086_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7314 a_32618_16488# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7315 vcm a_18162_68218# a_49286_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7316 a_7342_37405# a_6265_37039# a_7180_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7317 VSS a_3339_59879# a_8809_77117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7318 a_36234_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7319 a_38242_9492# a_18546_9490# a_38150_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X732 a_2369_18365# a_2325_17973# a_2203_18377# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X7320 vcm a_18162_63198# a_50290_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7321 a_28621_47381# a_28455_47381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7322 a_50198_67174# pmat.row_n[11] a_50690_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7323 VDD a_10053_15521# a_9943_15645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7324 a_19166_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7325 VSS a_3267_74817# a_3228_74691# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7326 a_2802_51727# a_2715_51969# a_2398_51859# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7327 a_49286_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7328 VDD a_8477_57141# a_4843_54826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X7329 a_3970_55311# a_4025_54965# a_3801_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X733 a_19828_27791# a_12987_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7330 a_12219_63303# a_12217_66389# a_12453_63151# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7331 a_26194_68178# a_18546_68220# a_26102_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7332 vcm a_18162_65206# a_23182_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7333 a_50594_22910# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7334 a_47186_21946# a_18162_21540# a_47278_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7335 a_23090_69182# pmat.row_n[13] a_23582_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7336 VSS pmat.sample_n a_18162_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X7337 a_1586_33927# a_1644_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7338 a_12543_40214# a_11565_39061# a_12471_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X7339 a_44266_18528# a_18546_18526# a_44174_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X734 a_6608_70455# a_5687_71829# a_6750_70262# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X7340 a_8013_73493# a_7847_73493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7341 pmat.col_n[12] _1183_.A2 a_31393_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7342 a_6244_40303# a_6127_40516# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7343 a_12227_12937# a_11711_12565# a_12132_12925# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X7344 VSS pmat.row_n[9] a_43566_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7345 VSS a_16837_40955# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X7346 vcm a_18162_10496# a_19166_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7347 clk_comp a_40399_36911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7348 a_29510_71230# pmat.rowon_n[15] a_29114_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7349 VDD a_9827_53379# a_9639_53339# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X735 VDD a_5651_66975# a_12150_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X7350 VDD a_18563_27791# a_41274_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7351 VDD a_5731_17455# a_2564_21959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7352 a_24186_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7353 a_3381_22717# a_3337_22325# a_3215_22729# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X7354 a_10287_61127# a_10286_60405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X7355 VSS a_13763_67191# a_12597_68279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7356 vcm a_18162_14512# a_45270_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7357 vcm a_18162_56170# a_44266_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7358 VSS a_16113_52271# a_16863_52815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X7359 a_20474_17890# nmat.rowon_n[6] a_20078_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X736 VSS cgen.dlycontrol2_in[4] a_29163_38545# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X7360 a_15210_51727# a_14491_51969# a_14647_51701# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X7361 a_44570_13874# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7362 VSS a_27155_31599# a_30121_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7363 VDD a_12345_36924# a_12757_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X7364 a_12431_69367# a_12719_69367# a_12665_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X7365 a_45270_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7366 a_6904_34863# a_5989_34863# a_6557_35105# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7367 a_35630_71552# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7368 a_27502_23914# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7369 a_28079_39913# a_26957_39867# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X737 vcm a_18162_67214# a_43262_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7370 VDD a_2847_38975# a_2834_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7371 VSS a_18203_48981# pmat.row_n[3] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X7372 a_31122_15922# pmat.row_n[7] a_31614_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7373 VSS pmat.row_n[13] a_31518_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7374 a_28202_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7375 a_39246_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7376 a_34626_57496# pmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7377 a_22178_14512# a_18546_14510# a_22086_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7378 a_7257_59049# a_3339_70759# a_6823_58951# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7379 a_21174_56130# a_18546_56172# a_21082_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X738 VDD a_46449_46261# a_45112_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7380 a_22199_30287# a_41731_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7381 VDD a_33719_34191# a_33825_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7382 VDD a_1923_61759# a_8996_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7383 a_23634_32509# a_2007_25597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X7384 a_27198_8488# a_18546_8486# a_27106_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7385 result_out[4] a_1644_59861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7386 a_24490_16886# nmat.rowon_n[7] a_24094_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7387 VSS pmat.row_n[5] a_21478_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7388 a_11091_26311# a_4523_21276# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7389 a_11347_36950# a_10651_37683# a_11347_37277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X739 VDD a_9749_19061# a_7693_22365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7390 a_38242_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7391 a_10515_24233# a_9075_28023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7392 a_24895_36341# a_12069_36341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7393 VDD a_4831_40303# a_5233_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7394 VSS a_11133_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X7395 VSS pmat.row_n[4] a_34530_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7396 VSS pmat.row_n[7] a_46578_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7397 a_4241_44111# a_3325_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7398 a_43566_60186# pmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7399 a_43566_19898# nmat.col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X74 VSS a_6976_32375# a_5963_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X740 a_47186_7890# VDD a_47678_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7400 a_31297_31849# a_31210_31751# a_30412_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7401 VSS a_40349_40726# a_39413_40956# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X7402 a_35306_46831# a_35186_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.9e+11p pd=3.8e+06u as=0p ps=0u w=650000u l=150000u
X7403 a_25190_55126# a_18546_55168# a_25098_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7404 a_5329_54965# a_5730_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7405 a_1644_66933# a_1823_66941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7406 a_25590_59504# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7407 inp_analog pmat.sw ctopp VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7645e+12p ps=2.191e+07u w=1.9e+06u l=220000u M=4
X7408 a_47278_72194# a_18546_72236# a_47186_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7409 a_44666_22512# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X741 a_26239_39095# a_26276_39429# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X7410 a_12132_12925# a_10845_12559# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7411 a_9050_15101# a_4383_7093# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7412 VSS a_2289_29397# a_2237_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7413 pmat.rowon_n[6] a_10515_15055# a_14462_61839# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X7414 a_23486_63198# pmat.rowon_n[7] a_23090_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7415 VDD a_11435_58791# a_14011_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X7416 VDD a_4679_28853# a_4379_28548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7417 a_51294_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7418 a_8581_56053# a_8363_56457# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X7419 VDD a_2648_29397# a_9913_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X742 a_16311_28327# a_45019_38645# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=0p ps=0u w=650000u l=150000u M=8
X7420 a_2405_17455# a_2228_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7421 a_42857_32481# a_42791_32375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7422 a_20170_17524# a_18546_17522# a_20078_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7423 VDD nmat.rowon_n[6] a_37146_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7424 a_30409_48463# a_28901_48437# a_19283_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X7425 a_51598_71230# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7426 a_35230_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7427 a_27623_52521# a_16311_28327# a_27405_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7428 a_14372_14191# a_11435_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7429 a_25319_42359# a_24197_42405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X743 a_36854_44527# a_36677_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7430 pmat.rowon_n[6] a_11067_16359# a_14379_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X7431 a_48190_72194# VDD a_48682_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7432 a_22787_34709# a_22963_35041# a_22915_35101# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X7433 VDD nmat.rowon_n[1] a_21082_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7434 a_48682_21508# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7435 a_48282_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7436 a_45178_14918# a_18162_14512# a_45270_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7437 a_2080_52815# a_1643_52789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7438 vcm a_18162_13508# a_21174_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7439 a_35138_70186# a_18162_70226# a_35230_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X744 a_25190_60146# a_18546_60188# a_25098_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7440 a_38642_13476# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7441 a_8723_11510# a_8472_11739# a_8264_11703# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7442 VDD nmat.rowon_n[12] a_42166_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7443 a_27502_64202# pmat.rowon_n[8] a_27106_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7444 a_36538_9858# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7445 a_46084_42051# a_32405_32463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7446 vcm a_18162_12504# a_34226_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7447 VDD nmat.sample_n a_18162_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X7448 VDD nmat.rowon_n[2] a_25098_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7449 a_22178_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X745 a_25590_64524# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7450 a_49194_13914# a_18162_13508# a_49286_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7451 a_19459_35279# a_19282_35279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7452 a_28202_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7453 a_25098_62154# a_18162_62194# a_25190_62154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7454 VSS pmat.row_n[1] a_46578_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7455 a_25042_31375# a_24160_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X7456 VDD a_4675_54599# a_3199_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7457 a_6244_34863# a_6127_35076# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7458 vcm a_18162_71230# a_46274_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7459 ctopn clk_ena ctopn VSS sky130_fd_pr__nfet_01v8 ad=2.7645e+12p pd=2.191e+07u as=0p ps=0u w=1.9e+06u l=220000u M=2
X746 a_28506_59182# pmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7460 VSS a_10851_30485# a_6927_30503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X7461 VDD pmat.rowoff_n[4] a_28110_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7462 vcm a_18162_19532# a_20170_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7463 a_30210_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7464 VDD a_12368_35823# a_12474_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7465 a_3551_6202# a_4254_7351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X7466 a_26194_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7467 a_13909_66959# a_13327_70741# a_13763_67191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7468 VDD a_2791_57703# a_3123_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7469 VDD pmat.rowon_n[10] a_49194_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X747 vcm a_18162_12504# a_39246_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7470 a_46674_63520# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7471 vcm a_18162_18528# a_33222_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7472 a_44849_45717# a_29937_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7473 VDD pmat.rowon_n[5] a_50198_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7474 a_12646_51549# a_12559_51325# a_12242_51435# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7475 a_12449_40693# a_12116_40871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7476 a_3295_23060# a_3387_22869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X7477 a_32522_17890# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7478 VDD nmat.rowon_n[4] a_41162_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7479 VSS a_7457_62037# a_7072_62037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X748 a_22086_61150# pmat.row_n[5] a_22578_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7480 a_23182_71190# a_18546_71232# a_23090_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7481 a_2325_42997# a_2107_43401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X7482 a_6999_15645# a_2411_16101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X7483 a_9317_47349# a_9099_47753# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7484 a_19166_61150# a_18546_61192# a_19074_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7485 a_42166_68178# a_18162_68218# a_42258_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7486 VSS a_8193_61493# a_7808_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7487 nmat.rowon_n[1] a_14195_7119# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7488 VSS a_4135_37815# a_2839_38101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7489 VDD pmat.rowon_n[7] a_23090_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X749 VSS cgen.dlycontrol1_in[3] a_28247_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X7490 a_43170_8894# pmat.row_n[0] a_43662_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7491 VDD _1194_.B1 a_12081_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X7492 VDD a_8673_7093# a_8563_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7493 a_5320_27023# a_4712_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.8675e+11p pd=3.79e+06u as=0p ps=0u w=650000u l=150000u M=2
X7494 a_5967_5461# a_6170_5739# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7495 a_39580_30287# a_39496_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7496 VDD a_20499_31274# a_9307_31068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7497 a_16131_29429# a_12437_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7498 a_19074_8894# pmat.row_n[0] a_19566_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7499 a_19746_27791# a_10441_21263# a_19828_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X75 VSS a_10245_51335# a_9919_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8025e+11p ps=3.77e+06u w=650000u l=150000u
X750 a_30118_69182# a_18162_69222# a_30210_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7500 a_19526_28335# a_7840_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X7501 a_34134_10902# a_18162_10496# a_34226_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7502 a_24094_71190# pmat.row_n[15] a_24586_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7503 a_45178_59142# a_18162_59182# a_45270_59142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7504 a_38770_50755# a_25879_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7505 a_45270_20536# a_18546_20534# a_45178_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7506 a_25494_8854# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7507 a_29606_8456# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7508 a_28110_69182# a_18162_69222# a_28202_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7509 a_15420_44007# a_14261_44219# a_15324_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X751 VSS pmat.row_n[1] a_32522_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7510 VDD a_31152_48071# a_32371_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7511 VDD pmat.rowon_n[6] a_27106_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7512 a_11645_68619# a_10864_68565# a_11559_68619# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7513 a_32218_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7514 a_11877_56079# a_6927_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X7515 a_13529_37253# a_13837_36893# a_13503_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7516 a_1644_58229# a_1823_58237# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7517 VSS a_41481_52245# pmat.col[22] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7518 nmat.rowoff_n[1] a_14839_7119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X7519 a_11347_40214# a_11317_40188# a_11275_40214# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X752 a_43262_10496# a_18546_10494# a_43170_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7520 a_4349_62313# a_4317_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X7521 a_10839_11989# a_12967_12863# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7522 a_22178_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7523 a_49194_58138# a_18162_58178# a_49286_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7524 a_35534_63198# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7525 a_36142_18934# pmat.row_n[10] a_36634_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7526 VSS nmat.en_bit_n[0] a_36538_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7527 VDD a_5363_70543# a_7953_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7528 a_40650_16488# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7529 VSS pmat.row_n[13] a_25494_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X753 VSS a_10651_35507# a_10591_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X7530 a_22482_66210# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7531 VSS a_7521_47081# a_9367_53511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7532 a_18546_12502# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7533 a_49194_17930# pmat.row_n[9] a_49686_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7534 VSS a_11927_27399# a_11885_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7535 VSS pmat.row_n[15] a_49590_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7536 a_20078_23954# pmat.row_n[15] a_20570_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7537 VSS a_10441_21263# a_19746_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7538 a_20078_19938# a_18162_19532# a_20170_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7539 a_40315_43177# a_39193_43131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X754 a_33467_46261# a_40047_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X7540 a_50198_12910# pmat.row_n[4] a_50690_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7541 a_11834_52931# a_10641_52815# a_11752_52931# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7542 a_17113_39141# a_13503_39069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X7543 a_5991_23983# a_5547_24233# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X7544 a_1781_9308# a_10383_13077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X7545 a_33130_22950# pmat.row_n[14] a_33622_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7546 a_26194_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7547 a_23090_55126# a_18162_55166# a_23182_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7548 a_25850_48981# a_25839_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7549 VSS pmat.row_n[7] a_39550_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X755 a_1846_72107# a_2124_72123# a_2080_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7550 a_4533_38279# a_7355_37013# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7551 a_47975_46831# a_47724_47081# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X7552 a_43566_13874# nmat.rowon_n[10] a_43170_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7553 VDD a_2847_20479# a_2834_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7554 a_26498_65206# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7555 VDD a_11149_36924# a_11561_36950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7556 nmat.col[12] ANTENNA__1184__B1.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=0p ps=0u w=650000u l=150000u M=2
X7557 a_26594_17492# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7558 a_26498_23914# pmat.rowoff_n[15] a_26102_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7559 a_4031_40455# a_2935_38279# a_4265_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X756 a_8851_63669# a_8695_63937# a_8996_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7560 a_23090_14918# pmat.row_n[6] a_23582_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7561 cgen.dlycontrol4_in[5] a_1591_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7562 pmat.col_n[25] _1192_.B1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X7563 VDD pmat.rowoff_n[7] a_30118_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7564 a_24094_18934# a_18162_18528# a_24186_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7565 a_38041_30485# a_7717_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7566 vcm a_18162_64202# a_44266_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7567 a_44174_68178# pmat.row_n[12] a_44666_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7568 a_45009_43817# a_43720_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.25e+11p pd=2.65e+06u as=0p ps=0u w=1e+06u l=150000u
X7569 VDD a_25879_31591# a_39757_50700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X757 a_12196_34215# a_10953_34951# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X7570 VDD pmat.rowon_n[3] a_47186_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7571 a_3305_27791# a_2847_28095# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X7572 VSS pmat.en_C0_n a_20474_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7573 cgen.dlycontrol3_in[4] a_1591_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X7574 VDD a_28915_50959# a_47407_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7575 a_47147_44655# a_46896_44905# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X7576 a_29510_56170# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7577 a_9335_51727# a_9084_51843# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X7578 VDD a_6800_44629# a_6830_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7579 a_31122_66170# a_18162_66210# a_31214_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X758 a_29510_7850# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7580 a_8673_7093# a_8455_7497# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7581 a_1846_55123# a_2124_55107# a_2080_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7582 a_27106_13914# pmat.row_n[5] a_27598_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7583 a_2629_65327# a_2250_65693# a_2557_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7584 a_31614_11468# nmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7585 a_21174_64162# a_18546_64204# a_21082_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7586 a_7072_52093# a_6835_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7587 a_21574_68540# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7588 a_9323_28879# a_9217_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7589 a_7067_70262# a_6292_65479# a_6608_70455# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X759 VDD a_13641_23439# a_31371_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7590 a_14197_67279# a_13327_70741# a_13763_67191# VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X7591 a_26515_41271# a_25393_41317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X7592 a_10913_55535# a_10409_53903# a_10815_55785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X7593 a_22915_35101# a_11041_38772# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7594 VDD a_2319_52789# a_2250_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X7595 a_1846_74283# a_2163_74173# a_2121_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X7596 VDD a_1899_35051# a_6641_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7597 a_25190_63158# a_18546_63200# a_25098_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7598 vcm a_18162_60186# a_22178_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7599 a_25590_67536# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X76 a_23090_24958# VDD a_23582_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X760 pmat.sample a_21815_42351# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X7600 vcm a_18162_15516# a_39246_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7601 a_1757_40853# a_1591_40853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7602 a_22086_64162# pmat.row_n[8] a_22578_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7603 a_29308_44869# a_29404_44869# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7604 a_43262_13508# a_18546_13506# a_43170_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7605 a_12403_24527# a_7026_24527# a_12295_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7606 a_10999_41046# a_10817_41046# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7607 vcm a_18162_10496# a_40250_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7608 VDD a_4859_31274# a_4471_30724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7609 a_10570_69679# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X761 a_3305_27791# a_2847_28095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7610 a_50594_71230# pmat.rowon_n[15] a_50198_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7611 a_35138_63158# pmat.row_n[7] a_35630_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7612 a_14911_31965# a_14287_31599# a_14803_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X7613 a_28525_43655# a_27785_43131# a_28848_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7614 VSS a_10515_15055# a_14287_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7615 a_78165_39738# a_78261_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7616 VSS a_29937_31055# a_46752_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7617 a_20257_49667# a_19283_49783# a_20175_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7618 VSS pmat.row_n[14] a_25494_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7619 VSS a_31695_43439# a_31801_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X762 VDD a_33283_42333# a_33309_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X7620 a_47278_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7621 VSS a_16911_51959# a_14839_66103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X7622 a_3305_15823# a_2847_16127# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7623 VDD a_3173_25045# a_3203_25398# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7624 a_83094_10383# ANTENNA__1190__B1.DIODE a_82788_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7625 a_7301_73487# a_6787_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7626 VDD a_2375_18708# a_1895_18170# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7627 VDD pmat.rowon_n[0] a_32126_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7628 a_7527_11510# a_7276_11739# a_7068_11703# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X7629 a_45178_22950# a_18162_22544# a_45270_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X763 VDD a_2315_44124# a_4070_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X7630 a_6800_22869# a_3351_27249# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X7631 a_42258_19532# a_18546_19530# a_42166_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7632 VSS a_3866_57399# a_5541_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7633 a_9155_17455# a_8305_20871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X7634 a_34593_43493# a_33283_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X7635 a_6381_72105# a_2407_49289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X7636 a_37542_61190# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7637 VDD a_31539_51946# pmat.col[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7638 vcm a_18162_21540# a_21174_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7639 a_44570_62194# pmat.rowon_n[6] a_44174_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X764 VDD a_45019_38645# a_46229_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=8
X7640 VSS pmat.row_n[10] a_41558_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7641 a_29825_52271# a_24867_53135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7642 a_12531_42583# nmat.sw VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7643 a_27502_72234# VDD a_27106_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7644 vcm a_18162_20536# a_34226_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7645 VDD nmat.sample_n a_18162_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X7646 a_36278_29967# a_35520_30083# a_35715_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7647 a_4898_29199# a_2648_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7648 VSS a_45064_44807# a_44628_45717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7649 a_22178_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X765 a_3069_69367# a_2727_58470# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X7650 VSS a_4516_21531# a_6661_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7651 VSS a_4719_30287# a_9176_50345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7652 a_10728_77661# a_10291_77269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7653 a_5361_72719# a_5271_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7654 pmat.row_n[5] a_21883_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X7655 a_2319_72092# a_2163_71997# a_2464_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7656 vcm a_18162_57174# a_42258_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7657 VDD a_18277_37620# a_14712_37429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7658 VDD a_46211_50095# a_24867_53135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X7659 a_12032_59887# a_9135_60967# a_11932_59887# VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X766 VDD nmat.rowon_n[4] a_33130_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7660 VSS a_11487_69653# a_11433_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X7661 VDD a_35186_47375# a_36532_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X7662 VDD a_2215_47375# a_7201_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X7663 a_42562_14878# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7664 a_11133_44581# a_10651_44211# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X7665 a_41515_27497# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7666 a_31518_59182# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7667 pmat.col_n[22] _1187_.A2 a_41335_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X7668 a_25494_24918# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7669 a_31518_17890# nmat.rowon_n[6] a_31122_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X767 a_20170_22544# a_18546_22542# a_20078_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7670 a_13423_55369# a_13073_54997# a_13328_55357# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X7671 nmat.col[28] _1194_.B1 a_83238_4175# VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u M=4
X7672 a_12075_24847# a_11897_21263# a_11987_24847# VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=0p ps=0u w=650000u l=150000u
X7673 VSS a_18597_31599# a_43543_32151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7674 a_12309_36483# a_22357_35877# a_23479_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7675 a_46674_71552# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7676 ctopn nmat.sw inn_analog VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.102e+12p ps=8.76e+06u w=1.9e+06u l=220000u M=4
X7677 a_9221_77129# a_8031_76757# a_9112_77129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X7678 VDD a_7313_74005# a_7343_74358# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7679 VDD ANTENNA__1190__A1.DIODE a_37743_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X768 a_11067_16359# a_18487_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7680 a_12235_62723# a_12199_62621# a_12163_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7681 a_20170_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7682 a_46182_61150# a_18162_61190# a_46274_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7683 a_7436_16519# a_4976_16091# a_7578_16694# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X7684 VSS a_11019_71543# a_11345_70773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7685 a_32218_56130# a_18546_56172# a_32126_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7686 VDD a_2199_13887# a_6788_5853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7687 a_29114_71190# a_18162_71230# a_29206_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7688 a_28506_15882# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7689 a_11949_21237# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X769 comp.adc_comp_circuit_0.adc_comp_buffer_0.in comp.adc_comp_circuit_0.adc_comp_buffer_1.in VSS VSS sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X7690 VSS pmat.row_n[5] a_32522_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7691 nmat.col[12] a_10883_3303# a_14558_3311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X7692 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7693 a_25839_49783# a_30687_48071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X7694 VDD nmat.rowon_n[1] a_19074_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7695 vcm a_18162_58178# a_19166_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7696 VDD pmat.rowon_n[15] a_23090_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7697 VSS a_10045_19677# a_10151_19637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7698 vcm a_18162_18528# a_41254_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7699 VDD nmat.rowon_n[14] a_23090_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X77 a_28849_48783# a_29076_48695# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X770 a_51202_58138# a_18162_58178# a_51294_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7700 VSS a_11703_48156# a_11634_48285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X7701 VDD a_22879_41781# a_11921_41814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7702 a_8178_31421# a_1923_31743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7703 a_23182_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7704 a_47582_69222# pmat.rowon_n[13] a_47186_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7705 VSS pmat.row_n[10] a_44570_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7706 VDD _1184_.A2 a_83196_3561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7707 VDD a_5651_66975# a_11711_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X7708 a_4505_74005# a_4259_73807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X7709 VSS a_10651_37683# a_10591_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X771 pmat.col[1] ANTENNA__1197__B.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7710 VSS a_2021_11043# a_6607_10615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X7711 a_42658_23516# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7712 a_42258_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7713 VDD a_15657_52317# a_15757_52535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X7714 a_83630_3311# _1184_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7715 a_2122_13779# a_2439_13889# a_2397_14013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X7716 a_5537_47081# a_5173_45993# a_5621_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7717 a_21082_21946# a_18162_21540# a_21174_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7718 a_16381_35286# a_16745_34427# a_17808_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7719 a_34978_31599# a_33684_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X772 VDD config_2_in[1] a_1591_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7720 a_24565_34789# a_23700_36391# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X7721 VDD pmat.rowon_n[14] a_27106_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7722 pmat.col[8] a_13091_28327# a_27986_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X7723 VDD nmat.rowon_n[5] a_35138_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7724 VDD a_10811_77437# a_10772_77563# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7725 a_2325_26401# a_2107_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7726 a_21478_66210# pmat.rowon_n[10] a_21082_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7727 VSS pmat.row_n[9] a_48586_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7728 a_31214_17524# a_18546_17522# a_31122_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7729 VDD nmat.rowon_n[6] a_48190_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X773 a_26102_60146# pmat.row_n[4] a_26594_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7730 VDD nmat.rowon_n[15] a_39154_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7731 pmat.row_n[12] a_19491_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X7732 VSS pmat.row_n[0] a_35534_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7733 a_43170_15922# a_18162_15516# a_43262_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7734 a_46274_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7735 a_51202_8894# pmat.row_n[0] a_51694_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7736 a_5331_28309# a_5156_28335# a_5510_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7737 VDD a_1586_18231# a_1591_20181# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7738 a_36142_69182# a_18162_69222# a_36234_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7739 a_2107_18377# a_1591_18005# a_2012_18365# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X774 a_35230_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7740 a_20063_32143# a_19439_32149# a_19955_32521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X7741 VSS pmat.row_n[1] a_38546_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7742 a_45574_8854# nmat.rowon_n[15] a_45178_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7743 VDD vcm.sky130_fd_sc_hd__buf_4_0.A a_77428_40594# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7744 a_31122_57134# pmat.row_n[1] a_31614_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7745 a_40250_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7746 a_42562_55166# VSS a_42166_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7747 a_17702_30287# a_12461_29673# a_17702_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X7748 a_18546_20534# nmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7749 a_18176_39429# a_17113_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X775 a_20695_32447# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7750 a_25494_65206# pmat.rowon_n[9] a_25098_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7751 vcm a_18162_13508# a_32218_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7752 a_39246_66170# a_18546_66212# a_39154_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7753 a_49686_13476# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7754 a_12437_28585# a_12175_27221# a_12521_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X7755 VDD a_10167_64239# a_10569_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7756 VDD nmat.rowon_n[4] a_39154_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7757 VDD pmat.rowon_n[12] a_43170_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7758 a_23090_63158# a_18162_63198# a_23182_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7759 a_31518_12870# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X776 a_34134_68178# a_18162_68218# a_34226_68178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7760 VSS a_20439_27247# a_33785_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7761 a_34148_28111# a_9411_2215# a_33845_27765# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X7762 a_14919_30287# a_13479_26935# a_14465_29575# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X7763 VDD a_43776_30287# a_46023_32937# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X7764 a_28506_56170# pmat.rowon_n[0] a_28110_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7765 a_37146_8894# a_18162_8488# a_37238_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7766 vcm a_18162_72234# a_44266_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7767 VDD nmat.rowon_n[10] a_26102_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7768 a_41162_22950# pmat.row_n[14] a_41654_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7769 comp_latch comp.adc_nor_latch_0.QN a_55610_40254# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X777 pmat.col[29] a_47764_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X7770 VDD a_1591_13103# a_1769_13103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7771 a_44266_60146# a_18546_60188# a_44174_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7772 a_11207_31764# a_11299_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X7773 a_23280_32521# a_22365_32149# a_22933_32117# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X7774 VDD pmat.rowon_n[11] a_47186_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7775 a_44666_64524# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7776 a_7805_55563# a_1769_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7777 VSS pmat.row_n[7] a_20474_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7778 a_47278_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7779 VSS a_3663_9269# a_5173_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X778 VSS a_9463_53511# a_11752_52931# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7780 a_83092_13103# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X7781 a_42658_7452# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7782 VSS a_2944_56872# a_2882_56989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X7783 VSS a_39781_41245# a_39473_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7784 a_34530_23914# pmat.rowoff_n[15] a_34134_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7785 VDD a_10697_75218# a_10699_75119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X7786 VSS pmat.row_n[6] a_33526_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7787 a_30514_18894# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7788 a_2325_36469# a_2107_36873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X7789 a_45589_31599# a_38851_28327# a_45505_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X779 a_27619_36649# a_26497_36603# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X7790 a_21174_72194# a_18546_72236# a_21082_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7791 a_47582_22910# nmat.rowon_n[1] a_47186_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7792 VDD a_32371_50247# a_32319_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7793 VSS a_1923_69823# a_6325_77295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7794 a_15259_31029# a_11067_30287# a_15477_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X7795 a_34226_71190# a_18546_71232# a_34134_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7796 VDD pmat.rowon_n[8] a_21082_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7797 VDD a_13327_70741# a_14347_69831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7798 a_45178_60146# pmat.row_n[4] a_45670_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7799 VDD a_2879_57487# a_4541_64561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X78 VSS vcm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u M=80
X780 a_51202_8894# a_18162_8488# a_51294_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7800 VDD VDD a_28110_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7801 VSS VDD a_24490_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7802 a_42307_31756# a_41949_30761# a_43179_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7803 VSS a_16163_43413# a_15921_38550# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7804 a_7255_71829# a_7431_71829# a_7383_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X7805 a_16324_36911# a_16147_36911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7806 a_38642_55488# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7807 vcm a_18162_23548# a_39246_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7808 a_22086_72194# VDD a_22578_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7809 a_43262_21540# a_18546_21538# a_43170_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X781 VDD VDD a_34134_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7810 VDD a_5363_70543# a_5423_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7811 VSS a_17996_41831# a_17959_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X7812 a_22578_60508# pmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7813 a_39246_11500# a_18546_11498# a_39154_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7814 a_35138_71190# pmat.row_n[15] a_35630_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7815 VSS pmat.row_n[12] a_50594_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7816 a_17900_36391# a_16837_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X7817 a_6772_61839# a_5731_58951# a_6681_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X7818 VSS a_14379_6567# a_14839_7119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7819 VSS pmat.row_n[2] a_38546_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X782 a_51202_17930# pmat.row_n[9] a_51694_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7820 a_9135_26409# a_2952_25045# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X7821 a_47126_29673# a_38851_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X7822 VSS a_3305_27791# a_7023_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7823 a_36538_61190# pmat.rowon_n[5] a_36142_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7824 a_13278_51549# a_12520_51451# a_12715_51420# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7825 a_25590_12472# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7826 VSS a_6283_31591# a_37471_32149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7827 VDD a_1959_12791# a_1959_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7828 VSS a_2411_16101# a_7153_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7829 a_4328_6409# a_3413_6037# a_3981_6005# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X783 VSS pmat.row_n[15] a_51598_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7830 VSS _1184_.A2 a_33227_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X7831 VDD a_24737_30485# a_24160_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7832 a_20474_67214# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7833 a_29206_22544# a_18546_22542# a_29114_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7834 a_2307_45199# a_1683_45205# a_2199_45577# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X7835 vcm a_18162_7484# a_39246_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7836 a_50594_56170# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7837 a_47186_18934# pmat.row_n[10] a_47678_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7838 VSS VDD a_47582_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7839 a_11889_56399# a_11835_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X784 VDD a_11067_64015# a_15163_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X7840 a_41254_69182# a_18546_69224# a_41162_69182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7841 a_51694_16488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7842 a_8861_24527# a_8831_24501# a_8607_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X7843 VSS a_3951_77055# a_3885_77129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X7844 a_33526_66210# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7845 VDD a_25647_37607# a_21219_36885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X7846 a_37238_59142# a_18546_59184# a_37146_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7847 a_49286_7484# a_18546_7482# a_49194_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7848 a_38242_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7849 VDD a_1781_9308# a_2507_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X785 a_4257_49667# a_3983_49911# a_4175_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7850 a_33423_47695# a_6664_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=8
X7851 VSS pmat.row_n[8] a_37542_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7852 a_2325_38645# a_2107_39049# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7853 VSS a_17139_30503# a_24857_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X7854 a_2192_49159# a_1769_13103# a_2334_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7855 a_41558_14878# nmat.rowon_n[9] a_41162_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7856 a_3951_77055# a_1923_69823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7857 VDD a_3325_20175# a_5797_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7858 a_20570_63520# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7859 VDD ANTENNA__1395__A1.DIODE a_33327_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X786 vcm a_18162_18528# a_38242_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7860 VSS a_1923_61759# a_9913_62973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7861 a_8885_67325# a_8819_67197# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7862 a_30514_59182# pmat.rowon_n[3] a_30118_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7863 a_24586_18496# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7864 a_3142_9839# a_2021_9563# a_3056_9839# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X7865 a_45270_68178# a_18546_68220# a_45178_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7866 vcm a_18162_65206# a_42258_65166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7867 a_42166_69182# pmat.row_n[13] a_42658_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7868 pmat.en_bit_n[1] nmat.en_bit_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X7869 VDD a_11159_23145# a_13798_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.6e+11p ps=5.72e+06u w=1e+06u l=150000u
X787 a_48282_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7870 vcm a_18162_55166# a_38242_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7871 a_8013_25615# a_7665_25731# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7872 a_38150_59142# pmat.row_n[3] a_38642_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7873 a_23280_32521# a_22199_32149# a_22933_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7874 a_36142_9898# pmat.row_n[1] a_36634_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7875 a_35138_18934# a_18162_18528# a_35230_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7876 a_3069_53609# a_2419_53351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7877 cgen.dlycontrol4_in[3] a_1591_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7878 a_4653_53359# a_4587_53505# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7879 VSS a_4737_21561# a_4671_21629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X788 a_12295_24527# a_11892_21959# a_12075_24847# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X7880 a_2629_58799# a_2250_59165# a_2557_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7881 a_27502_57174# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7882 a_11133_34427# a_10651_35507# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X7883 VSS VDD a_31518_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7884 a_46674_9460# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7885 a_5725_76207# a_5497_73719# a_5737_76457# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7886 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7887 a_5968_77295# a_5725_76207# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7888 VSS a_25393_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X7889 a_43262_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X789 VSS a_3936_70197# a_3880_70543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7890 a_7066_35229# a_5989_34863# a_6904_34863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7891 vcm a_18162_66210# a_28202_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7892 a_39246_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7893 a_32218_64162# a_18546_64204# a_32126_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7894 a_40685_50639# a_21739_29415# pmat.col[21] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7895 a_28602_19500# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7896 a_32618_68540# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7897 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7898 VDD a_9135_60967# a_9525_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X7899 a_8453_46287# a_8051_46607# a_8289_46607# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X79 a_8511_10749# a_8257_10422# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X790 a_42258_16520# a_18546_16518# a_42166_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7900 a_35108_39655# a_33949_39867# a_35071_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X7901 a_46578_23914# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7902 VDD a_10651_35507# a_10677_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7903 a_9485_27247# a_9137_27253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7904 a_13331_74953# a_12981_74581# a_13236_74941# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X7905 VSS pmat.row_n[13] a_50594_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7906 VDD a_19086_34343# a_19091_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7907 a_20078_65166# pmat.row_n[9] a_20570_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7908 vcm a_18162_16520# a_37238_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7909 a_41254_14512# a_18546_14510# a_41162_14918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X791 VDD a_35786_47893# a_33957_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X7910 a_40250_56130# a_18546_56172# a_40158_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7911 vcm a_18162_60186# a_33222_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7912 a_33130_64162# pmat.row_n[8] a_33622_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7913 a_36538_15882# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7914 a_18546_69224# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7915 VSS pmat.row_n[5] a_40554_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7916 VSS a_2411_43301# a_6417_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7917 a_18162_64202# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X7918 VSS pmat.row_n[15] a_23486_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7919 a_20474_20902# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X792 VSS a_2847_20479# a_2781_20553# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X7920 VSS a_4523_21276# a_14369_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X7921 a_36617_43131# a_35752_43781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X7922 a_83178_13353# _1187_.A2 a_82787_13077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X7923 a_23090_56130# pmat.row_n[0] a_23582_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7924 a_34552_42919# a_33489_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X7925 VDD pmat.rowon_n[1] a_30118_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7926 a_45574_70226# pmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7927 a_33135_27247# _1154_.X nmat.col_n[11] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7928 a_27198_15516# a_18546_15514# a_27106_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7929 VSS a_12987_26159# a_14301_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X793 a_40554_7850# VDD a_40158_7890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7930 VDD a_20572_40517# a_20645_42044# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X7931 a_43170_23954# a_18162_23548# a_43262_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7932 VDD a_15899_47939# a_22063_46519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7933 a_25315_28335# a_22307_27791# a_25226_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X7934 a_29510_17890# nmat.rowon_n[6] a_29114_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7935 VSS a_36193_35805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X7936 a_2163_67645# a_1674_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7937 a_30514_12870# pmat.rowoff_n[4] a_30118_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7938 a_42562_63198# pmat.rowon_n[7] a_42166_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7939 VDD a_13091_52047# a_19759_48987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X794 a_43533_30761# a_28704_29568# a_43869_30511# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.71e+11p ps=9.18e+06u w=650000u l=150000u M=4
X7940 VSS a_39321_42333# a_39013_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7941 a_27106_55126# VDD a_27598_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7942 a_19423_37737# a_13597_37571# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X7943 a_10907_43222# a_10725_43222# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7944 VSS pmat.row_n[14] a_22482_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7945 a_48586_61190# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7946 vcm a_18162_21540# a_32218_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7947 a_50198_71190# a_18162_71230# a_50290_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7948 VSS a_6829_26703# a_9135_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.6875e+11p ps=5.65e+06u w=650000u l=150000u
X7949 vcm a_18162_11500# a_28202_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X795 VDD a_2325_27765# a_2215_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7950 a_2319_65564# a_2163_65469# a_2464_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7951 a_36634_24520# nmat.en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7952 a_30571_50959# a_41427_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7953 VDD nmat.rowon_n[1] a_40158_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7954 vcm a_18162_58178# a_40250_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7955 a_27502_10862# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7956 VDD a_11823_46973# a_11784_47099# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7957 a_13443_39095# a_13837_39069# a_13503_39069# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X7958 a_7383_71855# a_6292_65479# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7959 a_20175_49667# a_19584_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X796 a_37542_17890# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7960 a_39246_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7961 a_34887_41271# a_33765_41317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7962 a_4224_63401# a_3784_62607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7963 a_2983_48071# a_2847_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7964 a_15181_53135# a_10055_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X7965 VDD a_17007_50613# pmat.row_n[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7966 VSS a_36789_52245# pmat.col_n[17] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7967 nmat.col_n[6] a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X7968 a_47582_7850# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7969 a_37146_20942# pmat.row_n[12] a_37638_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X797 VSS pmat.row_n[7] a_41558_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7970 a_44666_72556# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7971 a_37146_16926# a_18162_16520# a_37238_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7972 VSS a_1586_8439# a_8399_6037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7973 a_2493_11477# a_2327_11477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7974 VDD nmat.rowon_n[2] a_44174_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7975 VSS a_2149_45717# a_2093_46070# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7976 vcm a_18162_69222# a_30210_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7977 a_41254_14512# a_18546_14510# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7978 VDD a_6553_53047# a_6559_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7979 VSS _1194_.A2 a_83238_4175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X798 a_44570_18894# nmat.rowon_n[5] a_44174_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7980 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.sky130_fd_sc_hd__buf_4_1.X vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X7981 a_1757_27797# a_1591_27797# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7982 a_44174_62154# a_18162_62194# a_44266_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7983 VSS a_32072_38567# a_32035_38825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X7984 a_31165_29199# a_21365_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7985 a_1881_55357# a_1846_55123# a_1643_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7986 a_27106_72194# a_18162_72234# a_27198_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7987 a_14925_24847# a_14371_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X7988 VSS pmat.row_n[4] a_29510_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7989 VSS pmat.row_n[11] a_29510_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X799 VSS a_1643_74005# a_1591_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7990 a_6330_33053# a_5253_32687# a_6168_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7991 VDD a_82788_9991# nmat.col_n[19] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X7992 a_31214_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7993 VDD nmat.rowon_n[10] a_34134_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7994 a_19470_66210# pmat.rowon_n[10] a_19074_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7995 a_14466_28879# a_13479_26935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7996 a_16612_39655# a_15549_39867# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X7997 a_6637_69367# a_3339_70759# a_6800_69251# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7998 a_30210_12504# a_18546_12502# a_30118_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7999 VDD VDD a_21082_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 VSS a_32687_46607# a_34850_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X80 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u M=530
X800 a_16966_29423# a_17306_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=0p ps=0u w=650000u l=150000u M=4
X8000 inp_analog clk_ena ctopp VDD sky130_fd_pr__pfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7075e+12p ps=2.185e+07u w=1.9e+06u l=220000u M=4
X8001 VDD pmat.rowoff_n[4] a_47186_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8002 VDD config_2_in[10] a_1591_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X8003 a_2764_45577# a_1683_45205# a_2417_45173# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8004 vcm a_18162_68218# a_34226_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8005 a_45270_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8006 a_38546_69222# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8007 VDD a_5138_65479# a_4508_65845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8008 a_14734_64015# a_11067_64015# a_14648_64015# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8009 a_21174_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X801 a_12792_58633# a_11877_58261# a_12445_58229# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X8010 VSS a_38905_28853# a_38851_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8011 a_1846_67755# a_2124_67771# a_2080_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8012 VSS pmat.row_n[11] a_42562_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8013 a_6568_59887# a_5939_60137# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X8014 a_9395_27791# a_8951_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8015 VSS a_16800_47213# a_16911_52423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8016 a_2319_54965# a_2124_55107# a_2629_55357# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X8017 a_34226_61150# a_18546_61192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8018 VDD a_2199_13887# a_1687_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8019 a_34530_7850# VDD a_34134_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X802 a_7995_54281# a_7479_53909# a_7900_54269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X8020 a_50690_7452# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8021 a_51598_17890# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8022 a_8560_54281# a_7479_53909# a_8213_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8023 a_18162_15516# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8024 a_38242_61150# a_18546_61192# a_38150_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8025 VSS a_12345_36924# a_12764_37277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8026 VDD a_13327_70741# a_13909_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8027 a_32126_21946# a_18162_21540# a_32218_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8028 a_13988_55369# a_12907_54997# a_13641_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8029 VSS a_16657_42567# a_17867_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X803 VDD nmat.sample_n a_18162_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X8030 VDD pmat.rowon_n[7] a_42166_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8031 nmat.col[3] _1194_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8032 a_28110_11906# a_18162_11500# a_28202_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8033 a_6975_34538# a_7067_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X8034 VDD nmat.rowon_n[5] a_46182_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8035 VDD a_28049_50613# pmat.col_n[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8036 VSS a_6283_31591# a_38391_48469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8037 a_10045_19677# a_3688_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8038 a_13985_40229# a_11773_39087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X8039 a_2325_20149# a_2107_20553# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X804 a_17996_40743# a_16837_40955# a_17900_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X8040 a_9759_62607# a_9135_62613# a_9651_62985# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X8041 VSS pmat.row_n[2] a_36538_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8042 VSS a_24407_31375# a_29915_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X8043 a_12243_16733# a_11619_16367# a_12135_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8044 VSS config_2_in[7] a_1591_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8045 a_25494_9858# nmat.rowon_n[14] a_25098_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8046 a_13236_74941# a_6292_65479# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8047 VSS pmat.row_n[12] a_19470_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8048 VSS a_1643_69653# a_1591_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8049 a_39154_61150# pmat.row_n[5] a_39646_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X805 a_8581_56053# a_8363_56457# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8050 a_14335_16519# a_11067_16359# a_14569_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8051 a_10681_12879# a_10471_12791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8052 vcm a_18162_19532# a_29206_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8053 a_47186_69182# a_18162_69222# a_47278_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8054 VSS pmat.row_n[1] a_49590_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8055 a_51294_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8056 vcm a_18162_14512# a_30210_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8057 a_37238_67174# a_18546_67216# a_37146_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8058 a_36234_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8059 a_28969_27765# a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X806 a_14471_4943# a_10883_3303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X8060 a_13633_71855# a_8491_47911# a_13158_71285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8061 a_5603_32687# a_5087_32687# a_5508_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X8062 VDD pmat.rowon_n[13] a_41162_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8063 a_36631_52047# a_24867_53135# pmat.col[17] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8064 VDD a_25931_27221# nmat.col[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8065 a_24673_52271# _1224_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8066 a_30210_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8067 a_20570_71552# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8068 a_41254_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8069 a_33322_46607# a_32687_46607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X807 VSS pmat.row_n[1] a_21478_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8070 a_43533_29423# a_38851_28327# a_43451_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8071 VDD a_16324_36911# a_16430_36911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8072 VDD pmat.rowon_n[8] a_19074_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8073 a_24186_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8074 a_23604_42919# a_22541_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X8075 a_26498_57174# pmat.rowon_n[1] a_26102_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8076 VSS a_2648_29397# a_9913_16950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8077 a_23479_43447# a_22361_41479# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X8078 a_41558_66210# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8079 vcm a_18162_63198# a_38242_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X808 a_45270_57134# a_18546_57176# a_45178_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8080 a_34134_7890# a_18162_7484# a_34226_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8081 a_38150_67174# pmat.row_n[11] a_38642_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8082 VSS a_7085_15055# a_7717_14735# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X8083 a_34277_38550# a_33765_39141# a_34887_39095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8084 a_42658_65528# pmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8085 a_19873_44219# a_19417_43990# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X8086 a_11665_72943# a_3339_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X8087 a_22578_8456# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8088 a_20445_50345# a_10515_13967# a_20349_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8089 a_45270_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X809 VDD a_45282_32143# ANTENNA__1196__A2.DIODE VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u M=16
X8090 a_42166_55126# a_18162_55166# a_42258_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8091 VSS a_10873_40693# a_11292_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8092 VSS pmat.row_n[7] a_31518_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8093 a_34425_50639# a_30571_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8094 a_28202_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8095 a_38546_22910# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8096 VDD a_6787_47607# a_8231_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X8097 a_42166_14918# pmat.row_n[6] a_42658_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8098 a_45670_17492# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8099 VSS pmat.row_n[12] a_42562_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X81 a_34552_36391# a_33309_36039# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X810 a_18272_42693# a_17113_42405# a_18176_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X8100 a_45574_23914# pmat.rowoff_n[15] a_45178_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8101 a_32218_72194# a_18546_72236# a_32126_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8102 a_5508_18543# a_5257_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8103 a_25098_24958# VDD a_25590_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8104 VDD a_47592_35643# a_47591_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8105 a_5092_41935# a_4149_41941# a_4984_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X8106 VSS a_3571_13627# a_11711_12565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8107 a_26552_36165# a_25393_35877# a_26456_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8108 a_2464_61519# a_2250_61519# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8109 a_35534_15882# pmat.rowoff_n[7] a_35138_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X811 a_2250_67869# a_2124_67771# a_1846_67755# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X8110 a_36545_51727# a_34705_51959# pmat.col[17] VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8111 VDD a_6787_47607# a_7111_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8112 a_28110_56130# a_18162_56170# a_28202_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8113 VDD a_32305_51335# a_31631_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X8114 a_17996_41831# a_16837_42043# a_17900_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8115 VDD nmat.rowon_n[6] a_22086_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8116 vcm a_18162_24552# a_37238_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8117 VSS a_7663_27247# a_7840_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X8118 vcm a_18162_66210# a_36234_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8119 a_46182_13914# pmat.row_n[5] a_46674_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X812 a_42166_58138# pmat.row_n[2] a_42658_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8120 a_26779_47197# a_26155_46831# a_26671_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X8121 a_10853_75119# a_9581_73487# a_10781_75119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8122 a_20170_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8123 a_40250_64162# a_18546_64204# a_40158_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8124 a_50690_11468# nmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8125 a_49686_55488# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8126 a_29114_23954# pmat.row_n[15] a_29606_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8127 VSS a_7658_71543# a_13183_72405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8128 a_40650_68540# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8129 a_33130_72194# VDD a_33622_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X813 ANTENNA__1190__A1.DIODE a_47449_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X8130 a_29114_19938# a_18162_19532# a_29206_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8131 a_36634_58500# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8132 a_33622_21508# nmat.col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8133 a_3685_66237# a_3207_65845# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8134 a_33222_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8135 a_30118_14918# a_18162_14512# a_30210_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8136 a_10513_24135# a_10239_20291# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8137 a_18162_72234# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X8138 a_16863_29239# a_14691_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8139 VDD a_5935_46983# a_5621_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X814 a_13459_28111# a_30663_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X8140 a_39550_14878# nmat.rowon_n[9] a_39154_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8141 VSS pmat.row_n[3] a_36538_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8142 VSS a_42683_32375# a_40903_32375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8143 VDD a_20645_42044# a_20251_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8144 VSS a_16083_50069# a_18521_46837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8145 VSS pmat.row_n[0] a_25494_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8146 a_19689_41317# a_19233_41479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X8147 a_19074_15922# pmat.row_n[7] a_19566_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8148 vcm a_18162_8488# a_43262_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8149 VSS pmat.row_n[13] a_19470_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X815 a_18035_27791# a_7840_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8150 a_23582_13476# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8151 a_20078_10902# pmat.row_n[2] a_20570_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8152 VSS pmat.row_n[2] a_49590_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8153 a_40966_46653# a_40837_46261# a_40467_46261# VSS sky130_fd_pr__nfet_01v8 ad=1.155e+11p pd=1.39e+06u as=3.465e+11p ps=2.49e+06u w=420000u l=150000u
X8154 VSS a_22199_30287# a_43072_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8155 vcm a_18162_60186# a_41254_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8156 VDD VSS a_26102_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8157 VDD a_33839_46805# a_33797_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8158 a_41162_64162# pmat.row_n[8] a_41654_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8159 vcm a_18162_8488# a_19166_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X816 VSS a_7658_71543# a_12815_74581# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8160 a_27198_23548# a_18546_23546# a_27106_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8161 VSS a_12431_69367# a_11487_69653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X8162 VDD a_14340_19783# pmat.rowoff_n[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X8163 a_34134_13914# a_18162_13508# a_34226_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8164 VSS a_27794_28879# a_28442_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X8165 VSS a_30913_38779# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X8166 a_13739_51701# a_14174_51859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8167 a_12954_12559# a_11877_12565# a_12792_12937# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8168 a_5843_44905# a_4128_46983# a_5747_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8169 pmat.rowoff_n[11] a_14460_60137# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X817 VSS pmat.row_n[6] a_45574_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8170 a_10621_21583# a_10498_19631# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X8171 a_29206_8488# a_18546_8486# a_29114_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8172 VDD a_7999_31359# a_7986_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8173 a_26498_10862# nmat.rowon_n[13] a_26102_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8174 a_2858_59475# a_3136_59459# a_3092_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8175 a_2969_55785# a_2791_57703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8176 a_22281_49667# a_18547_51565# a_22199_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8177 a_4608_41909# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8178 vcm a_18162_71230# a_31214_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8179 a_35230_15516# a_18546_15514# a_35138_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X818 VSS a_19965_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X8180 VSS a_5589_14967# a_5547_14735# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X8181 a_49286_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8182 a_11255_35862# a_11225_35836# a_11183_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X8183 a_10591_42089# a_10651_42035# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X8184 vcm a_18162_61190# a_27198_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8185 nmat.col[3] a_10883_3303# a_13086_4175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X8186 a_2847_23743# a_2672_23817# a_3026_23805# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8187 VSS a_33617_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X8188 vcm.sky130_fd_sc_hd__nand2_1_1.A vcm.sky130_fd_sc_hd__buf_4_0.A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8189 a_31614_63520# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X819 a_42562_11866# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8190 VDD pmat.rowoff_n[12] a_36142_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8191 a_6316_8903# a_6412_8725# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8192 a_39246_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8193 a_45556_27247# ANTENNA__1395__A1.DIODE a_45253_27221# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X8194 a_5383_48783# a_5411_48695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X8195 a_2215_47375# a_1775_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8196 a_25494_58178# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8197 a_22963_35041# a_10873_38517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8198 a_39550_71230# pmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8199 vcm a_18162_11500# a_36234_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X82 a_13236_74941# a_6292_65479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X820 a_39154_10902# a_18162_10496# a_39246_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8200 VDD a_28116_38567# a_28020_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8201 a_12783_18377# a_12337_18005# a_12687_18377# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X8202 a_37146_24958# a_18162_24552# a_37238_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8203 a_6829_46607# a_6637_46348# a_5935_46983# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8204 a_14751_28341# a_14365_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8205 vcm a_18162_10496# a_49286_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8206 a_41254_22544# a_18546_22542# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8207 a_37238_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8208 a_3295_23060# a_3387_22869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8209 VSS a_25997_42902# a_26331_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X821 a_31518_9858# nmat.rowon_n[14] a_31122_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8210 a_46109_51727# _1224_.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8211 VSS a_7343_16042# a_6679_15492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8212 a_16025_29469# a_14691_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8213 result_out[9] a_1644_66933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8214 VSS a_10049_60663# a_12032_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8215 a_30118_59142# a_18162_59182# a_30210_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8216 vcm a_18162_22544# a_26194_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8217 a_30210_20536# a_18546_20534# a_30118_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8218 a_44570_24918# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8219 VDD a_5651_66975# a_12237_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X822 a_2834_34141# a_1757_33775# a_2672_33775# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8220 a_50594_17890# nmat.rowon_n[6] a_50198_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8221 a_26194_10496# a_18546_10494# a_26102_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8222 a_44811_36469# a_44647_36201# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8223 VSS a_29825_30557# a_29931_30517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X8224 a_12213_53359# a_11737_53359# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.34e+11p pd=2.02e+06u as=0p ps=0u w=650000u l=150000u
X8225 VSS a_11149_36924# a_11568_37277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8226 vcm a_18162_16520# a_48282_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8227 _1192_.A2 a_47591_35407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8228 a_9666_32275# a_9944_32259# a_9900_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8229 a_40741_46565# a_40105_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X823 a_5363_70543# a_10795_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X8230 a_51294_56130# a_18546_56172# a_51202_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8231 VDD a_2672_28169# a_2847_28095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8232 VSS pmat.row_n[1] a_48586_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8233 a_34134_58138# a_18162_58178# a_34226_58138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8234 VSS a_12559_51325# a_12520_51451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8235 nmat.col[8] a_27763_27221# a_27535_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X8236 a_47582_15882# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8237 a_21082_18934# pmat.row_n[10] a_21574_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8238 VSS VDD a_21478_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8239 a_18162_23548# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X824 a_4865_12533# a_5331_13951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8240 a_25681_28879# a_25327_28992# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8241 VSS pmat.row_n[5] a_51598_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8242 a_7619_34102# a_6559_33767# a_7160_33927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8243 VDD a_29797_51701# pmat.col_n[10] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8244 VDD pmat.rowon_n[15] a_42166_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8245 a_34134_17930# pmat.row_n[9] a_34626_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8246 VSS pmat.row_n[15] a_34530_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8247 VDD pmat.rowon_n[5] a_38150_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8248 a_30140_43781# a_28981_43493# a_30044_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8249 VDD a_11067_27239# a_41699_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X825 a_31518_56170# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8250 a_9271_15101# a_7644_16341# a_8908_14967# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X8251 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8252 a_18546_15514# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X8253 a_4432_42313# a_3983_41941# a_4337_41935# VSS sky130_fd_pr__nfet_01v8 ad=1.44e+11p pd=1.52e+06u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X8254 a_40040_50639# _1183_.A2 pmat.col_n[19] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X8255 VDD a_21032_44007# a_20936_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X8256 a_25190_71190# a_18546_71232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8257 a_27502_18894# nmat.rowon_n[5] a_27106_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8258 VSS pmat.row_n[7] a_24490_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8259 a_6999_15645# a_6375_15279# a_6891_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X826 VSS VDD a_28506_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8260 a_26767_34967# cgen.dlycontrol1_in[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8261 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8262 a_9234_31094# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X8263 a_14257_16189# a_12447_16143# a_14185_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8264 a_36142_11906# a_18162_11500# a_36234_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8265 VDD a_12345_39100# a_12289_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8266 a_2121_71855# a_1643_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8267 a_28202_57134# a_18546_57176# a_28110_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8268 a_12195_38870# a_12013_38870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X8269 a_40554_66210# pmat.rowon_n[10] a_40158_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X827 a_15669_48169# nmat.sw a_15574_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X8270 VSS a_2422_29575# a_2882_31965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X8271 a_25098_58138# pmat.row_n[2] a_25590_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8272 a_50290_17524# a_18546_17522# a_50198_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8273 a_45178_8894# pmat.row_n[0] a_45670_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8274 a_27995_30287# a_23021_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8275 VDD pmat.rowon_n[3] a_32126_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8276 VSS pmat.row_n[6] a_28506_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8277 a_25494_11866# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8278 a_8722_53903# a_7645_53909# a_8560_54281# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8279 a_4945_30511# a_4901_30753# a_4779_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X828 a_25494_21906# nmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8280 a_29493_31375# a_29455_31293# a_29243_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8281 a_47678_24520# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8282 VDD a_17842_27497# a_40967_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8283 VSS a_30571_50959# a_46934_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X8284 VDD VDD a_19074_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8285 a_37238_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8286 VDD nmat.rowon_n[1] a_51202_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8287 a_77528_39738# vcm.sky130_fd_sc_hd__dlymetal6s6s_1_4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8288 a_32072_42919# a_30913_43131# a_31976_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8289 a_11569_14191# a_11525_14433# a_11403_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X829 a_2369_50095# a_2325_50337# a_2203_50095# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X8290 a_37542_64202# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8291 a_36617_42043# a_34924_41605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X8292 a_44570_65206# pmat.rowon_n[9] a_44174_65166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8293 a_27502_8854# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8294 VDD a_10985_44220# a_10591_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X8295 a_14385_49257# nmat.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X8296 VDD a_7255_71829# a_6602_72007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8297 vcm a_18162_13508# a_51294_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8298 VDD nmat.rowon_n[9] a_41162_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8299 a_34552_41831# a_33489_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X83 a_29206_59142# a_18546_59184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X830 vcm a_18162_24552# a_20170_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8300 a_17786_47081# a_11067_64015# a_17690_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8301 a_2882_72221# a_2163_71997# a_2319_72092# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X8302 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8303 a_42166_63158# a_18162_63198# a_42258_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8304 a_48190_20942# pmat.row_n[12] a_48682_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8305 VSS a_2419_53351# a_5065_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X8306 a_48190_16926# a_18162_16520# a_48282_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8307 VSS a_1923_61759# a_3445_66237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8308 VDD a_7415_29397# a_33101_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X8309 a_34530_57174# pmat.rowon_n[1] a_34134_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X831 a_25794_49007# a_25850_48981# a_18823_50247# VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X8310 VSS a_2835_13077# a_13593_8573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8311 VSS a_34724_44527# a_34830_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8312 VDD a_22963_42657# a_22787_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X8313 a_3119_22729# a_2769_22357# a_3024_22717# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X8314 a_22186_30485# a_15753_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X8315 a_22265_48579# a_18823_50247# a_22193_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8316 a_14287_57711# a_12447_16143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X8317 a_32256_44869# a_31097_44581# a_32219_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8318 vcm a_18162_15516# a_24186_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8319 a_47582_56170# pmat.rowon_n[0] a_47186_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X832 a_3307_77129# a_2861_76757# a_3211_77129# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X8320 a_1846_31851# a_2124_31867# a_2080_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8321 VDD a_1823_76181# a_4319_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8322 a_38150_12910# pmat.row_n[4] a_38642_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8323 VDD nmat.rowon_n[10] a_45178_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8324 a_42658_10464# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8325 a_27995_30287# a_28715_28879# a_28774_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X8326 VDD pmat.rowoff_n[15] a_28110_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8327 vcm a_18162_19532# a_50290_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8328 VDD a_2659_35015# a_4307_35639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8329 a_28110_64162# a_18162_64202# a_28202_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X833 a_28110_57134# pmat.row_n[1] a_28602_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8330 a_12479_39958# a_12228_39605# a_12020_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8331 a_32218_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8332 VDD a_2787_55535# a_2882_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8333 a_10217_54223# a_6559_33767# a_9871_53903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X8334 a_30610_8456# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8335 a_40250_72194# a_18546_72236# a_40158_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8336 a_36234_62154# a_18546_62196# a_36142_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8337 a_2215_43023# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8338 VDD pmat.rowon_n[13] a_39154_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8339 a_36634_66532# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X834 a_37238_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8340 VDD a_4956_59317# a_3956_59317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8341 VDD a_2199_13887# a_8996_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8342 a_30118_22950# a_18162_22544# a_30210_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8343 VDD pmat.rowon_n[8] a_40158_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8344 a_14458_58799# a_10515_13967# a_14372_58799# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8345 a_29206_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8346 a_49286_61150# a_18546_61192# a_49194_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8347 VDD a_15660_31029# a_15259_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8348 a_36142_56130# a_18162_56170# a_36234_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8349 a_9237_17455# a_8305_20871# a_9155_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X835 VSS a_16981_37462# a_16045_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X8350 VSS a_15420_41831# a_15383_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8351 a_22482_61190# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8352 VDD nmat.en_bit_n[1] pmat.en_bit_n[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X8353 a_12449_22895# a_5899_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8354 a_19074_66170# a_18162_66210# a_19166_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8355 VSS a_1586_33927# a_1591_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8356 a_19566_11468# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8357 a_41162_72194# VDD a_41654_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8358 VDD a_22085_42902# a_23512_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8359 VDD a_5046_67655# a_3838_70455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X836 VSS a_29076_48695# a_30219_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X8360 VSS a_7072_26311# a_6664_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8361 VSS a_28325_27221# nmat.col_n[8] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8362 a_37146_62154# pmat.row_n[6] a_37638_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8363 a_12133_9001# a_11731_8751# a_11969_8751# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X8364 VSS a_2411_16101# a_3381_22717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8365 VDD a_7415_29397# a_33515_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=8
X8366 VDD a_1591_14735# a_1769_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8367 nmat.rowon_n[4] a_14460_11177# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X8368 VSS pmat.row_n[2] a_47582_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8369 a_41654_60508# pmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X837 VDD pmat.rowon_n[15] a_49194_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8370 a_33719_44527# a_33542_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8371 a_4719_30287# a_5423_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8372 a_26498_60186# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8373 a_26498_19898# nmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8374 VDD pmat.en_bit_n[1] a_34134_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8375 a_5510_9295# a_4865_8181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X8376 a_43267_28879# a_43659_28853# a_21739_29415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X8377 a_35230_23548# a_18546_23546# a_35138_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8378 a_38531_51348# a_38575_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8379 a_4031_20884# a_4123_20693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X838 a_32618_55488# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8380 VDD VDD a_21082_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8381 a_29685_34954# clk_ena VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8382 VDD a_32367_51946# pmat.col[12] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X8383 vcm a_18162_8488# a_51294_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8384 a_38546_71230# pmat.rowon_n[15] a_38150_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8385 VSS a_17012_47349# a_14379_6567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X8386 a_48282_22544# a_18546_22542# a_48190_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8387 a_31614_71552# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8388 a_1644_57685# a_1591_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8389 a_27598_61512# pmat.col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X839 a_42258_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8390 a_31122_61150# a_18162_61190# a_31214_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8391 a_34530_10862# nmat.rowon_n[13] a_34134_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8392 a_6173_6575# a_5558_9527# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X8393 VSS a_43965_27221# nmat.col_n[23] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8394 a_50198_23954# pmat.row_n[15] a_50690_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8395 a_50198_19938# a_18162_19532# a_50290_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8396 VDD a_2952_25045# a_5070_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=2
X8397 a_14578_51727# a_14491_51969# a_14174_51859# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8398 VSS a_6283_31591# a_38391_47381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8399 VDD a_31339_31787# a_31297_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 VSS a_14491_51969# a_14452_51843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X840 vcm a_18162_23548# a_33222_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8400 a_40591_39095# a_39469_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8401 a_3354_74575# a_3228_74691# a_2950_74707# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=360000u l=150000u
X8402 a_29159_39783# cgen.dlycontrol2_in[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8403 a_43662_18496# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8404 a_43566_24918# VSS a_43170_24958# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8405 a_40158_15922# pmat.row_n[7] a_40650_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8406 a_37238_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8407 a_32522_69222# pmat.rowon_n[13] a_32126_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8408 a_28715_28879# a_28442_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8409 a_12061_74895# a_10515_75895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X841 VSS a_7129_57685# a_7063_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8410 a_32367_51946# a_32319_50345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X8411 VSS a_1643_54965# a_1591_54991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8412 a_11403_14191# a_10957_14191# a_11307_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8413 a_11188_73309# a_10751_72917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8414 a_2325_63669# a_2107_64073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X8415 a_21124_42919# a_19965_43131# a_21028_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X8416 a_46578_57174# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8417 a_46578_15882# pmat.rowoff_n[7] a_46182_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8418 VDD nmat.rowon_n[5] a_20078_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8419 a_29510_67214# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X842 a_22186_30485# a_15753_28879# a_23352_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.345e+12p ps=1.269e+07u w=1e+06u l=150000u M=4
X8420 a_42258_7484# a_18546_7482# a_42166_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8421 a_41878_29673# a_38905_28853# a_41786_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X8422 VSS pmat.row_n[9] a_33526_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8423 cgen.dlycontrol4_in[1] a_1626_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8424 VDD a_14336_48071# a_13462_48071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8425 vcm a_18162_24552# a_48282_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8426 VDD nmat.rowon_n[6] a_33130_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8427 VSS a_24407_31375# a_41876_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8428 vcm a_18162_66210# a_47278_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8429 VSS a_20310_28029# a_22015_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X843 a_22482_14878# nmat.rowon_n[9] a_22086_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8430 a_31214_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8431 a_51294_64162# a_18546_64204# a_51202_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8432 a_3579_15113# a_3229_14741# a_3484_15101# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8433 VDD nmat.rowon_n[7] a_14460_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X8434 VDD a_31263_28309# a_33775_29111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.25e+11p ps=2.85e+06u w=1e+06u l=150000u
X8435 a_7805_76001# a_6795_76989# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8436 a_51694_68540# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8437 a_19470_59182# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8438 a_12337_18005# a_12171_18005# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8439 a_45719_36495# a_43533_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X844 a_2107_43401# a_1757_43029# a_2012_43389# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8440 a_21082_69182# a_18162_69222# a_21174_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8441 a_47678_58500# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8442 a_13962_22671# a_11159_23145# a_13643_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.6875e+11p ps=4.35e+06u w=650000u l=150000u
X8443 VSS a_3751_64757# a_3697_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8444 VSS pmat.row_n[1] a_23486_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8445 a_39634_47375# a_38557_47381# a_39472_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8446 vcm a_18162_9492# a_23182_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8447 VSS pmat.row_n[3] a_47582_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8448 VDD a_8693_11769# a_8723_11510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8449 a_45921_42167# a_44774_40821# a_46084_42051# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X845 a_46912_34319# a_29937_31055# a_35244_32411# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X8450 a_24186_66170# a_18546_66212# a_24094_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8451 a_34626_13476# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8452 a_31976_42919# a_30913_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8453 VDD nmat.rowon_n[4] a_24094_19938# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8454 a_30121_31599# a_30219_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8455 VDD a_30543_40721# a_30403_40747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8456 VSS ANTENNA__1395__A2.DIODE a_83092_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8457 a_10029_26819# a_2952_25045# a_9957_26819# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8458 VSS a_7527_30676# a_7047_31226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8459 a_4461_46805# a_4128_46983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X846 VSS a_13653_35516# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X8460 a_10591_44265# a_10985_44220# a_10651_44211# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X8461 a_6800_22869# a_6651_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8462 a_14457_15823# a_14103_15936# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8463 VDD config_1_in[10] a_1626_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8464 a_2411_33749# a_2511_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X8465 a_3337_22325# a_3119_22729# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X8466 a_14369_57533# a_11067_16359# a_14287_57280# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8467 a_42166_56130# pmat.row_n[0] a_42658_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8468 a_28202_65166# a_18546_65208# a_28110_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8469 vcm a_18162_62194# a_25190_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X847 a_18162_7484# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8470 a_28602_69544# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8471 a_25098_66170# pmat.row_n[10] a_25590_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8472 a_23815_48981# a_23971_49140# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X8473 a_14453_31599# a_14287_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8474 a_36538_64202# pmat.rowon_n[8] a_36142_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8475 VDD nmat.rowon_n[14] a_25098_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8476 VDD pmat.rowon_n[11] a_32126_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8477 a_46274_15516# a_18546_15514# a_46182_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8478 vcm a_18162_12504# a_43262_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8479 a_9011_6409# a_8565_6037# a_8915_6409# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X848 VDD VSS a_41162_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8480 VDD ANTENNA__1197__A.DIODE a_41791_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X8481 a_21063_48723# a_21279_48999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X8482 VSS a_4421_70741# a_4036_70741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8483 VDD a_3909_17209# a_3939_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8484 a_4025_6397# a_3981_6005# a_3859_6409# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X8485 a_37238_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8486 a_33205_32143# a_32771_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X8487 a_3859_56311# a_2879_57487# a_4033_56417# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8488 a_4767_21302# a_4516_21531# a_4308_21495# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8489 a_46182_55126# VDD a_46674_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X849 a_28506_12870# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8490 VDD a_13503_39069# a_13529_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X8491 a_37542_72234# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8492 VDD a_8213_53877# a_8103_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8493 a_17159_47919# pmat.rowon_n[7] pmat.rowoff_n[4] VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X8494 a_32522_22910# nmat.rowon_n[1] a_32126_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8495 VSS pmat.row_n[14] a_41558_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8496 a_19166_17524# a_18546_17522# a_19074_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8497 a_29114_65166# pmat.row_n[9] a_29606_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8498 vcm a_18162_21540# a_51294_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8499 a_7527_30676# a_7619_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X85 VSS pmat.row_n[9] a_20474_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X850 VSS a_4061_63303# a_2467_63125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8500 vcm a_18162_11500# a_47278_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8501 a_36345_42567# a_36617_43131# a_37739_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8502 a_30118_60146# pmat.row_n[4] a_30610_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8503 VSS a_20616_27791# a_27339_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8504 a_45428_49007# a_44774_48695# a_45328_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X8505 a_9301_69679# a_9135_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8506 a_5747_44655# a_6141_44629# a_5597_44807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.665e+11p ps=2.12e+06u w=650000u l=150000u
X8507 a_1823_64213# a_2847_63999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8508 a_48190_24958# a_18162_24552# a_48282_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8509 VSS a_1586_18231# a_1591_18005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X851 a_6657_27497# a_4516_21531# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X8510 a_46578_10862# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8511 a_19074_57134# pmat.row_n[1] a_19566_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8512 a_23582_55488# pmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8513 a_83178_14735# _1183_.A2 a_82787_14709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8514 a_29510_20902# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8515 VDD a_13896_74953# a_14071_74879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8516 vcm a_18162_23548# a_24186_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8517 VSS pmat.row_n[5] a_44570_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8518 a_23090_9898# a_18162_9492# a_23182_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8519 a_22199_49667# a_19584_52423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X852 a_46523_39733# a_44444_32233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X8520 a_6793_56417# a_6175_60039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8521 a_47582_8854# nmat.rowon_n[15] a_47186_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8522 VSS pmat.row_n[15] a_27502_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8523 VDD a_13091_28327# a_29829_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X8524 a_24186_11500# a_18546_11498# a_24094_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8525 a_18546_56172# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8526 VDD a_9335_51727# a_10299_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8527 a_9133_6005# a_8915_6409# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8528 a_19470_12870# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8529 VSS pmat.row_n[2] a_23486_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X853 a_34948_50069# a_10883_3303# a_35171_50095# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X8530 a_4043_33535# a_3868_33609# a_4222_33597# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8531 VSS a_33283_42333# a_33223_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8532 vcm a_18162_59182# a_45270_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8533 a_21478_61190# pmat.rowon_n[5] a_21082_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8534 a_46182_72194# a_18162_72234# a_46274_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8535 VSS pmat.row_n[4] a_48586_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8536 a_12585_40443# a_15549_39867# a_16671_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X8537 a_45574_16886# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8538 VSS pmat.row_n[11] a_48586_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8539 VSS a_12116_40871# a_23883_40693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X854 VSS pmat.row_n[2] a_32522_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8540 a_33765_41317# a_33309_41479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X8541 a_50290_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8542 a_11883_62063# a_12107_62037# a_11711_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8543 a_36234_70186# a_18546_70228# a_36142_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8544 a_6469_21813# a_2683_22089# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8545 a_23700_39655# a_22541_39867# a_23604_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8546 a_43170_10902# a_18162_10496# a_43262_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8547 VDD _1154_.A a_36175_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8548 VDD VDD a_40158_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8549 a_32126_18934# pmat.row_n[10] a_32618_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X855 a_82778_4399# ANTENNA__1187__B1.DIODE nmat.col[21] VSS sky130_fd_pr__nfet_01v8 ad=1.2675e+12p pd=1.3e+07u as=3.64e+11p ps=3.72e+06u w=650000u l=150000u M=4
X8550 VSS VDD a_32522_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8551 a_29206_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8552 a_39154_8894# a_18162_8488# a_39246_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8553 VDD pmat.rowon_n[6] a_36142_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8554 a_36142_64162# a_18162_64202# a_36234_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8555 a_9092_31287# a_9307_31068# a_9234_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X8556 VSS a_47211_50069# a_11067_27239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X8557 a_6772_62927# a_5081_53135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8558 a_40250_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8559 a_22178_59142# a_18546_59184# a_22086_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X856 a_37680_41831# a_36617_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X8560 VDD nmat.rowon_n[1] a_49194_22950# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8561 a_7578_60214# a_4075_50087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8562 vcm a_18162_58178# a_49286_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8563 a_11014_71855# a_10699_72943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X8564 VDD a_26276_39429# a_26180_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8565 a_5919_52521# a_5785_48463# a_5823_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8566 VSS a_25209_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X8567 a_47026_45519# a_43720_32143# a_46940_45519# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X8568 a_12629_68047# a_12597_68279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8569 a_23182_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X857 vcm a_18162_55166# a_19166_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8570 a_25494_60186# pmat.rowon_n[4] a_25098_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8571 a_49286_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8572 VSS pmat.row_n[8] a_22482_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8573 a_25494_19898# nmat.rowon_n[4] a_25098_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8574 a_29825_30557# a_29455_31293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8575 a_44666_7452# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8576 a_40554_7850# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8577 a_37146_70186# pmat.row_n[14] a_37638_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8578 VDD nmat.rowon_n[9] a_39154_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8579 a_9112_77129# a_8197_76757# a_8765_76725# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X858 a_34530_67214# pmat.rowon_n[11] a_34134_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8580 a_2012_41213# a_1895_41018# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8581 VSS a_11067_64015# a_25280_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8582 result_out[8] a_1644_65845# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8583 a_30210_68178# a_18546_68220# a_30118_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8584 a_23807_41959# a_10767_39087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8585 a_51202_21946# a_18162_21540# a_51294_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8586 a_12585_37179# a_17113_35877# a_18235_35831# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8587 a_7005_41935# a_4128_46983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X8588 a_26194_58138# a_18546_58180# a_26102_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8589 vcm a_18162_55166# a_23182_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X859 vcm a_18162_9492# a_36234_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8590 a_47186_11906# a_18162_11500# a_47278_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8591 a_23090_59142# pmat.row_n[3] a_23582_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8592 VDD a_23707_40693# a_12197_41570# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8593 VSS VDD a_26498_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8594 a_2250_61519# a_2163_61761# a_1846_61651# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8595 a_12703_31055# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8596 a_51598_66210# pmat.rowon_n[10] a_51202_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8597 a_11925_53609# a_10641_52815# a_11737_53359# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8598 VDD a_1674_57711# a_9135_62613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8599 VSS a_1899_35051# a_5271_35407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X86 a_46578_56170# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X860 a_19074_59142# pmat.row_n[3] a_19566_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8600 VSS pmat.row_n[12] a_38546_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8601 VSS _1224_.X a_39219_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X8602 a_8919_71615# a_8744_71689# a_9098_71677# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8603 a_24186_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8604 VSS a_1925_26935# a_1738_26677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8605 VDD a_7037_70521# a_7067_70262# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8606 VSS a_1586_50247# a_1591_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8607 VSS a_8841_60405# a_8599_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X8608 a_21028_42919# a_19965_43131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8609 VSS a_27509_44219# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X861 vcm a_18162_15516# a_41254_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8610 a_14825_50095# a_14287_50345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8611 a_48586_64202# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8612 VDD a_1717_13647# a_6879_10473# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8613 a_20572_40517# a_19413_40229# a_20476_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8614 a_2651_49334# a_1769_13103# a_2192_49159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8615 a_18568_51959# a_16083_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X8616 a_31518_23914# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8617 a_3123_69135# a_2727_58470# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8618 pmat.rowon_n[10] a_10515_61839# a_14553_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8619 a_16113_52271# a_15757_52535# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X862 a_47582_66210# pmat.rowon_n[10] a_47186_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8620 a_35630_61512# pmat.col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8621 a_38546_56170# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8622 vcm a_18162_16520# a_22178_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8623 a_25190_19532# a_18546_19530# a_25098_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8624 a_13514_31421# a_1858_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8625 a_43262_69182# a_18546_69224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8626 a_40158_66170# a_18162_66210# a_40250_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8627 a_45574_57174# pmat.rowon_n[1] a_45178_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8628 a_39646_16488# nmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8629 a_28110_7890# a_18162_7484# a_28202_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X863 a_20315_29098# a_13643_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X8630 a_14094_15055# a_10515_61839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X8631 pmat.rowoff_n[8] a_25743_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8632 a_13073_26159# a_8013_25615# a_12987_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X8633 a_28506_67214# pmat.rowon_n[11] a_28110_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8634 vcm a_18162_15516# a_35230_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8635 a_21478_15882# nmat.col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8636 a_31103_28585# a_19405_28853# a_31021_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.8e+11p pd=2.76e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8637 VSS a_40105_47375# a_40741_46565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X8638 VSS a_1586_63927# a_8031_64789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8639 a_2007_42644# a_2051_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X864 a_38150_22950# pmat.row_n[14] a_38642_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8640 VSS pmat.row_n[7] a_50594_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8641 VSS a_46522_34293# a_46130_34639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8642 a_5403_67655# a_7099_74313# a_7301_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8643 a_40509_31849# a_38913_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X8644 a_2215_36495# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8645 a_22276_46831# a_21797_47081# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X8646 a_30514_70226# pmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8647 a_29217_41570# a_30913_42043# a_31976_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8648 VDD a_7497_11769# a_7527_11510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8649 VDD a_7370_27791# a_7663_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X865 a_46274_9492# a_18546_9490# a_46182_9898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8650 VDD a_15753_28879# a_22216_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X8651 a_6615_37039# a_6099_37039# a_6520_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X8652 a_12437_28335# a_12155_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8653 a_51294_72194# a_18546_72236# a_51202_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8654 a_44174_24958# VDD a_44666_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8655 a_47278_62154# a_18546_62196# a_47186_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8656 VSS a_3983_43567# a_2315_44124# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X8657 a_47678_66532# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8658 a_20474_62194# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8659 VDD pmat.rowon_n[8] a_51202_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X866 VDD pmat.rowoff_n[15] a_45178_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8660 VSS VDD a_19470_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8661 a_47186_56130# a_18162_56170# a_47278_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8662 a_33526_61190# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8663 a_6559_44431# a_4399_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X8664 VDD a_33109_52245# pmat.col[13] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8665 a_17113_41317# a_13503_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X8666 VDD a_46027_44905# a_46667_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X8667 a_48682_9460# nmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8668 a_12449_40693# a_12116_40871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8669 VDD pmat.rowon_n[0] a_41162_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X867 a_42658_20504# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8670 a_21574_24520# nmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8671 a_50290_7484# a_18546_7482# a_50198_7890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8672 a_48190_62154# pmat.row_n[6] a_48682_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8673 VSS a_35084_31599# a_35312_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X8674 VDD a_4036_67477# a_3983_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8675 VSS a_21867_34709# a_14773_37218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8676 a_24186_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8677 a_7131_19407# a_4976_16091# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X8678 VSS a_36663_34191# a_36769_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8679 VSS a_7658_71543# a_7847_73493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X868 a_6619_42479# a_6173_42479# a_6523_42479# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X8680 VSS pmat.row_n[13] a_38546_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8681 a_10867_43447# a_11261_43421# a_10927_43421# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X8682 VDD a_5351_19913# a_14471_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8683 vcm a_18162_70226# a_25190_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8684 VDD VSS a_45178_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8685 vcm a_18162_9492# a_31214_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8686 a_13565_3087# ANTENNA__1196__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X8687 a_36538_72234# VDD a_36142_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8688 a_25590_23516# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8689 a_22086_20942# pmat.row_n[12] a_22578_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X869 a_42258_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8690 a_22086_16926# a_18162_16520# a_22178_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8691 a_25190_19532# a_18546_19530# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8692 vcm a_18162_20536# a_43262_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8693 a_46274_23548# a_18546_23546# a_46182_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8694 VSS a_43720_32143# a_45064_44807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X8695 nmat.col_n[22] a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X8696 VDD pmat.rowon_n[9] a_28110_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8697 a_50594_67214# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8698 VSS a_2621_48981# a_2555_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8699 pmat.rowon_n[4] a_10515_61839# a_14094_60751# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X87 VDD a_10409_53903# a_10815_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X870 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8700 a_28202_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8701 a_7370_27791# a_7023_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X8702 VDD a_1586_33927# a_1591_33775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8703 a_45574_10862# nmat.rowon_n[13] a_45178_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8704 a_22745_27247# ANTENNA__1395__A2.DIODE a_22527_27221# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8705 a_41227_29423# a_40954_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8706 a_28602_14480# nmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8707 a_28506_20902# pmat.rowoff_n[12] a_28110_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8708 a_40554_59182# pmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8709 a_26102_15922# a_18162_15516# a_26194_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X871 a_13855_24847# a_13563_24527# a_13769_24847# VSS sky130_fd_pr__nfet_01v8 ad=1.47e+11p pd=1.54e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8710 VDD pmat.rowoff_n[4] a_32126_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8711 vcm a_18162_61190# a_46274_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8712 pmat.rowon_n[4] a_11067_16359# a_14011_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X8713 a_30210_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8714 a_23486_69222# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8715 VSS a_2411_16101# a_3841_15101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8716 VSS a_3866_57399# a_3824_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8717 a_50690_63520# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8718 a_14864_34215# a_13801_34427# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X8719 a_20811_42359# a_19689_42405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X872 a_16890_36911# a_16713_36911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8720 a_10873_39605# a_30679_40513# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X8721 VSS a_1923_69823# a_1881_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8722 a_2882_59165# a_2124_59067# a_2319_59036# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8723 VSS nmat.sw a_14427_46519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8724 a_38150_71190# a_18162_71230# a_38242_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8725 a_14369_12265# a_10239_14183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=0p ps=0u w=1e+06u l=150000u
X8726 a_29114_10902# pmat.row_n[2] a_29606_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8727 VDD a_43132_48071# a_42292_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8728 a_44570_58178# pmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8729 a_23182_61150# a_18546_61192# a_23090_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X873 a_45178_64162# a_18162_64202# a_45270_64162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8730 a_35252_52271# a_11067_27239# a_34949_52245# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X8731 a_18546_64204# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8732 a_27502_68218# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8733 a_22178_8488# a_18546_8486# a_22086_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8734 a_18162_18528# nmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X8735 VDD a_14113_43132# a_13719_43177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8736 VDD nmat.rowon_n[5] a_31122_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8737 VSS a_11927_27399# a_12987_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8738 a_12052_71671# a_8491_47911# a_11980_71671# VSS sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8739 a_41297_27221# a_21739_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X874 a_30219_48783# a_28901_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8740 vcm a_18162_67214# a_45270_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8741 VDD a_45019_38645# a_44757_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=8
X8742 a_9135_60967# a_9231_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8743 VSS pmat.row_n[15] a_35534_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8744 a_9493_66415# a_9643_66389# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8745 VSS pmat.row_n[2] a_21478_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8746 VDD a_36854_44527# a_37731_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8747 a_24094_61150# pmat.row_n[5] a_24586_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8748 a_34611_44265# a_11113_39747# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X8749 a_32126_69182# a_18162_69222# a_32218_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X875 a_32218_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8750 VSS pmat.row_n[1] a_34530_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8751 VDD pmat.rowon_n[14] a_36142_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8752 a_28110_16926# pmat.row_n[8] a_28602_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8753 a_45270_10496# a_18546_10494# a_45178_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8754 a_6265_6825# a_5558_9527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X8755 VDD a_1781_9308# a_2193_9334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X8756 VDD a_2944_67752# a_2882_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8757 VDD a_5768_9527# a_5325_9269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8758 a_31122_9898# a_18162_9492# a_31214_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8759 a_22178_67174# a_18546_67216# a_22086_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X876 VDD pmat.rowoff_n[7] a_35138_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8760 a_49590_7850# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8761 a_36234_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8762 VDD a_25695_28111# a_34942_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8763 a_24033_28111# a_11067_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8764 a_23663_44535# a_23700_44869# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X8765 a_50198_65166# pmat.row_n[9] a_50690_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8766 a_11113_36483# a_19689_34789# a_20752_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8767 a_19166_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8768 VSS a_3688_17179# a_10239_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8769 a_13605_71017# a_12809_69679# a_13533_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X877 a_20075_43447# a_18953_43493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X8770 VSS VDD a_40554_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8771 a_40158_57134# pmat.row_n[1] a_40650_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8772 a_2080_74397# a_1643_74005# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8773 vcm a_18162_63198# a_23182_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8774 a_50594_20902# nmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8775 a_23090_67174# pmat.row_n[11] a_23582_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8776 VSS a_13335_31359# a_13269_31433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X8777 a_44266_16520# a_18546_16518# a_44174_16926# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8778 VDD a_1586_8439# a_1591_15829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8779 VSS a_25315_28335# a_24374_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X878 VDD a_28116_37479# a_28020_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X8780 VSS a_1923_61759# a_1881_61885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8781 a_39550_17890# nmat.col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8782 VDD a_14336_46983# a_13830_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8783 a_30210_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8784 VSS pmat.row_n[7] a_43566_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8785 a_40554_12870# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8786 VDD a_9135_60967# a_9195_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8787 nmat.col[18] _1183_.A2 a_82998_2473# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X8788 a_23486_22910# nmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8789 VSS a_10967_77532# a_10898_77661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X879 a_13620_50095# a_4991_69831# a_13140_50247# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8790 VDD a_11435_58791# a_14287_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8791 a_13549_8181# a_13331_8585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X8792 a_30610_17492# nmat.col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8793 a_30514_23914# pmat.rowoff_n[15] a_30118_23954# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8794 a_7896_11079# a_8111_11209# a_8038_11254# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X8795 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8796 VSS pmat.row_n[1] a_41558_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8797 a_48586_72234# pmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8798 a_7201_62313# a_5784_52423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8799 a_14342_55357# a_1957_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X88 a_45193_50639# a_17139_30503# pmat.col[26] VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X880 VDD nmat.rowon_n[9] a_48190_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8800 a_19470_61190# pmat.rowon_n[5] a_19074_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8801 a_44174_58138# pmat.row_n[2] a_44666_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8802 a_24833_34191# a_24667_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8803 a_20474_15882# pmat.rowoff_n[7] a_20078_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8804 a_9583_10121# a_14071_8511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8805 a_44570_11866# nmat.col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8806 a_51598_9858# nmat.rowon_n[14] a_51202_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8807 a_31976_41831# a_30913_42043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8808 a_6127_40516# a_5233_40553# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8809 a_27502_21906# nmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X881 a_36753_46805# a_30111_47911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8810 a_7109_15521# a_6891_15279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8811 vcm a_18162_24552# a_22178_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8812 vcm a_18162_66210# a_21174_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8813 VSS pmat.row_n[6] a_42562_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8814 a_31122_13914# pmat.row_n[5] a_31614_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8815 a_39246_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8816 a_27502_9858# nmat.rowon_n[14] a_27106_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8817 a_34626_55488# pmat.en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8818 VDD a_9112_77129# a_9287_77055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8819 vcm a_18162_23548# a_35230_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X882 a_46274_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8820 a_21574_58500# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8821 a_30765_40513# a_24833_40719# a_30679_40513# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8822 a_11255_36189# a_11001_35862# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8823 VSS _1224_.X a_82778_4399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8824 a_3615_71631# a_11071_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X8825 a_24490_14878# nmat.rowon_n[9] a_24094_14918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8826 VSS pmat.row_n[3] a_21478_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8827 a_18162_10496# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8828 a_38242_7484# a_18546_7482# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8829 VDD VSS a_43170_24958# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X883 a_43170_12910# a_18162_12504# a_43262_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8830 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8831 a_13683_24847# a_11337_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8832 VSS pmat.row_n[2] a_34530_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8833 VDD a_28247_34191# a_29391_36395# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8834 VSS a_7896_11079# a_7276_11739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8835 a_36637_28111# a_26891_28327# a_36419_28023# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8836 a_77882_39738# a_77978_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8837 VDD a_2163_74173# a_2124_74299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8838 a_43913_31849# a_41949_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8839 a_12651_35823# a_12474_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X884 VDD a_1959_10615# a_1959_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X8840 vcm.sky130_fd_sc_hd__buf_4_2.A vcm.sky130_fd_sc_hd__dlymetal6s6s_1_5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8841 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8842 VDD a_13503_37981# a_13529_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X8843 VDD a_3911_44431# a_4313_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X8844 a_47278_70186# a_18546_70228# a_47186_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8845 VSS a_6637_69367# a_5497_62839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8846 a_49590_66210# pmat.rowon_n[10] a_49194_66170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8847 a_45282_32143# a_44571_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X8848 VSS a_11565_39061# a_11597_39453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X8849 a_44666_20504# nmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X885 VDD a_28325_27221# nmat.col_n[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8850 VDD pmat.rowoff_n[15] a_47186_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8851 VDD a_26283_42325# a_14497_42658# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8852 VDD VDD a_51202_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8853 a_44266_16520# a_18546_16518# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8854 VSS pmat.row_n[7] a_19470_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8855 VSS a_2411_33749# a_2369_36861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8856 a_47186_64162# a_18162_64202# a_47278_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8857 a_20474_8854# nmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8858 a_24586_8456# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8859 a_51294_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X886 a_22178_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8860 a_13331_8585# a_12815_8213# a_13236_8573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X8861 a_10219_30877# a_9595_30511# a_10111_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X8862 a_7107_44905# a_2935_38279# a_7011_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X8863 a_17808_44869# a_16745_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8864 a_20170_15516# a_18546_15514# a_20078_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8865 a_34226_72194# a_18546_72236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8866 VDD pmat.rowoff_n[7] a_37146_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8867 a_8957_67325# a_8891_66964# a_8885_67325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8868 a_48190_70186# pmat.row_n[14] a_48682_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8869 VDD pmat.rowoff_n[12] a_21082_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X887 VSS a_6451_67655# a_6794_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X8870 a_5351_60663# a_4025_54965# a_5696_60751# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X8871 a_48282_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8872 a_45178_12910# a_18162_12504# a_45270_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8873 a_9309_20291# a_4613_19087# a_9227_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8874 a_24186_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8875 a_41558_61190# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8876 VDD a_15747_50069# a_9963_13967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X8877 a_14558_5263# ANTENNA__1190__A2.DIODE VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X8878 a_22357_39141# a_20848_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X8879 a_24490_71230# pmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X888 a_49194_63158# a_18162_63198# a_49286_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8880 vcm a_18162_11500# a_21174_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8881 a_38642_11468# nmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8882 a_23063_36885# a_23239_37217# a_23191_37277# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8883 a_22086_24958# a_18162_24552# a_22178_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8884 VDD a_1923_53055# a_3016_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8885 a_17842_27497# _0467_ a_17424_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X8886 a_5257_69679# a_4719_69929# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8887 VDD nmat.sample_n a_18162_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X8888 vcm a_18162_10496# a_34226_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8889 a_22178_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X889 VDD a_26479_32117# a_25688_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8890 a_40676_46653# a_40645_46519# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X8891 a_45187_38129# a_46815_37013# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X8892 a_28202_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8893 a_25098_60146# a_18162_60186# a_25190_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8894 a_46934_52047# ANTENNA__1197__A.DIODE a_46848_52047# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8895 VSS pmat.row_n[12] a_49590_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8896 a_36936_49257# a_33957_48437# a_36265_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.05e+11p pd=7.61e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8897 a_45567_47081# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8898 VDD a_3956_59317# a_3894_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8899 VSS a_11455_50237# a_11416_50363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X89 a_5277_37039# a_2563_34837# a_5205_37039# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X890 a_36142_66170# a_18162_66210# a_36234_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8900 a_30819_40191# cgen.dlycontrol4_in[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8901 VDD comp.adc_inverter_1.out comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=3.32e+06u w=500000u l=150000u M=4
X8902 VDD a_34948_50069# pmat.col[15] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8903 VDD a_27913_42333# a_27519_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8904 a_11541_46831# a_11506_47083# a_11071_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8905 vcm a_18162_8488# a_45270_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8906 a_26102_23954# a_18162_23548# a_26194_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8907 a_30085_30761# a_23021_29199# a_30013_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8908 a_25647_39783# a_25671_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8909 VDD nmat.rowon_n[13] a_28110_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X891 a_22482_71230# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8910 a_43566_58178# pmat.rowon_n[2] a_43170_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8911 a_20329_35431# a_20438_35431# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8912 a_9213_53903# a_8735_54207# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8913 a_50690_71552# pmat.col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8914 a_13726_22351# a_3305_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X8915 a_39469_39141# a_38972_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X8916 VSS a_12263_50959# a_19441_47491# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X8917 a_26498_68218# pmat.rowon_n[12] a_26102_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8918 VDD pmat.rowon_n[8] a_49194_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8919 a_16945_31375# nmat.en_bit_n[1] a_15660_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X892 VDD _1179_.X a_83178_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X8920 a_46674_61512# pmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8921 VSS a_33084_40743# a_33047_41001# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8922 VSS _1192_.B1 a_25776_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8923 vcm a_18162_16520# a_33222_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8924 VDD a_7631_55687# a_3345_62839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X8925 VSS cgen.dlycontrol1_in[1] a_25755_34343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X8926 a_37638_19500# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8927 VDD a_12155_20719# a_12167_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X8928 a_3395_19465# a_3045_19093# a_3300_19453# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8929 vcm a_18162_71230# a_19166_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X893 VSS a_21219_36885# a_21857_36950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8930 a_32522_15882# nmat.col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8931 a_8155_20969# a_7533_19087# a_7935_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8932 VDD pmat.rowon_n[0] a_39154_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8933 VSS a_7068_11703# a_6853_14967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8934 a_3262_59343# a_3136_59459# a_2858_59475# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=360000u l=150000u
X8935 a_12587_32182# a_9135_60967# a_12128_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8936 VDD a_82788_10357# nmat.col_n[24] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X8937 a_19566_63520# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8938 VDD a_21977_52245# pmat.col[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8939 VDD pmat.rowon_n[5] a_23090_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X894 a_36634_11468# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8940 VDD a_13459_28111# a_46765_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8941 cgen.dlycontrol1_in[3] a_1591_33231# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X8942 a_37892_32509# a_5179_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8943 a_9919_51959# a_9427_50095# a_10159_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X8944 a_45645_45895# a_7109_29423# a_45808_45993# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8945 a_5265_28335# a_4075_28335# a_5156_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X8946 a_33436_44527# a_33259_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8947 nmat.en_bit_n[0] pmat.en_bit_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8948 a_45178_57134# a_18162_57174# a_45270_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8949 VDD a_6787_47607# a_12437_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X895 VSS a_11149_36924# a_11093_36950# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8950 a_10979_43222# a_10949_43124# a_10907_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X8951 VSS a_21124_39655# a_21087_39913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8952 a_11793_56079# a_11444_55535# a_11711_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8953 a_21082_11906# a_18162_11500# a_21174_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8954 a_3184_74575# a_2747_74549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8955 a_28110_67174# a_18162_67214# a_28202_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8956 VDD pmat.rowon_n[4] a_27106_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8957 a_30210_8488# a_18546_8486# a_30118_8894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8958 VDD a_20711_34191# nmat.sample VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X8959 a_14747_2767# a_10883_3303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X896 a_9557_17705# a_8305_20871# a_9485_17705# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8960 a_50290_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8961 VDD a_2046_30184# a_6743_31061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8962 VDD pmat.sample_n a_18162_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X8963 a_32618_24520# nmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8964 a_23329_37462# a_22725_38053# a_23788_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8965 a_22178_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8966 a_3181_52093# a_2802_51727# a_3109_52093# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8967 VSS a_1923_31743# a_2369_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8968 a_4061_63303# a_4266_63303# a_4224_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8969 a_38546_17890# nmat.rowon_n[6] a_38150_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X897 VDD a_2621_48981# a_2651_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8970 VDD a_8583_29199# a_21341_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X8971 a_36142_16926# pmat.row_n[8] a_36634_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8972 a_11285_41046# a_11113_40835# a_11071_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8973 a_8257_54269# a_8213_53877# a_8091_54281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8974 VSS pmat.row_n[11] a_25494_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8975 a_22482_64202# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8976 a_49194_15922# pmat.row_n[7] a_49686_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8977 VSS pmat.row_n[13] a_49590_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8978 a_20078_21946# pmat.row_n[13] a_20570_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8979 a_20078_17930# a_18162_17524# a_20170_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X898 VSS a_4043_22869# a_2835_13077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X8980 a_44266_24552# a_18546_24550# a_44174_24958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8981 a_5704_11471# a_5173_9839# a_5602_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=150000u
X8982 a_19409_40719# a_19143_41085# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8983 a_43262_66170# a_18546_66212# a_43170_66170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8984 a_50198_10902# pmat.row_n[2] a_50690_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8985 a_26515_35831# a_25393_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X8986 a_39246_56130# a_18546_56172# a_39154_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8987 a_2563_34837# a_2847_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8988 a_5821_18785# a_5603_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8989 a_12461_29673# a_8583_29199# a_12651_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X899 a_20078_24958# a_18162_24552# a_20170_24552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8990 a_33130_20942# pmat.row_n[12] a_33622_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8991 a_9176_50345# a_7373_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8992 a_18180_38341# a_17021_38053# a_18143_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X8993 a_33130_16926# a_18162_16520# a_33222_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8994 VDD pmat.rowon_n[2] a_43170_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8995 VSS pmat.sample_n a_18162_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X8996 VSS pmat.row_n[5] a_39550_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8997 a_43566_11866# nmat.rowon_n[12] a_43170_11906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8998 a_25232_31375# a_24374_29941# a_25042_31055# VSS sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=2.86e+11p ps=2.18e+06u w=650000u l=150000u
X8999 a_7631_15253# a_7456_15279# a_7810_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9 vcm a_18162_19532# a_27198_19532# VSS sky130_fd_pr__nfet_01v8 ad=1.54997e+14p pd=1.73788e+09u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X90 VDD nmat.rowon_n[6] a_20078_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X900 a_12792_58633# a_11711_58261# a_12445_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X9000 a_36532_46805# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9001 a_24002_47741# a_2263_43719# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9002 a_32522_56170# pmat.rowon_n[0] a_32126_56130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9003 VDD nmat.rowon_n[5] a_29114_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9004 a_26594_15484# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9005 a_23090_12910# pmat.row_n[4] a_23582_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9006 a_26498_21906# nmat.rowon_n[2] a_26102_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9007 a_22895_47893# a_22459_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X9008 a_6608_70455# a_6292_65479# a_6750_70589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9009 VDD nmat.rowon_n[10] a_30118_13914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X901 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9010 vcm a_18162_62194# a_44266_62154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9011 a_44174_66170# pmat.row_n[10] a_44666_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9012 VDD a_13091_52047# a_17183_52251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9013 a_5185_51727# a_2389_45859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9014 a_34887_36919# a_33765_36965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9015 a_11597_39453# a_11327_39087# a_11507_39087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9016 a_46109_44905# a_44966_43255# a_46027_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9017 a_2193_9334# a_2021_9563# a_1979_9334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X9018 VDD start_conversion_in a_1591_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X9019 a_10873_36341# a_29391_36395# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X902 a_19566_21508# nmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9020 a_27106_11906# pmat.row_n[3] a_27598_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9021 a_10676_30511# a_9595_30511# a_10329_30753# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X9022 a_21174_62154# a_18546_62196# a_21082_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9023 VDD pmat.rowon_n[13] a_24094_69182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9024 a_38242_17524# a_18546_17522# a_38150_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9025 VSS a_3417_47919# a_3983_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9026 a_21574_66532# pmat.col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9027 a_34226_61150# a_18546_61192# a_34134_61150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9028 a_11842_59887# a_9135_60967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X9029 a_21082_56130# a_18162_56170# a_21174_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X903 a_22725_38053# a_20848_38341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X9030 vcm a_18162_68218# a_43262_68178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9031 a_8197_64789# a_8031_64789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9032 a_10195_30186# a_10287_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X9033 a_22753_50345# a_19584_52423# a_22657_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9034 a_47186_8894# pmat.row_n[0] a_47678_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9035 a_1644_77813# a_1823_77821# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9036 VDD a_2422_29575# a_2882_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X9037 a_16837_36603# a_13779_36595# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X9038 a_25590_65528# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9039 a_22086_62154# pmat.row_n[6] a_22578_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X904 vcm a_18162_10496# a_32218_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9040 a_12227_58633# a_11711_58261# a_12132_58621# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X9041 vcm a_18162_13508# a_39246_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9042 a_25931_27221# a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X9043 VSS pmat.row_n[2] a_32522_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9044 a_43262_11500# a_18546_11498# a_43170_11906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9045 VSS pmat.row_n[15] a_46578_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9046 a_37553_46607# a_33467_46261# a_36532_46805# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9047 a_35138_61150# pmat.row_n[5] a_35630_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9048 a_4243_54991# a_3970_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9049 a_29510_8854# nmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X905 a_19166_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9050 a_44266_24552# a_18546_24550# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9051 VDD a_19176_35279# a_19282_35279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9052 a_27411_46805# a_27236_46831# a_27590_46831# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9053 VDD a_5821_18785# a_5711_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9054 a_45246_41167# a_44382_40847# a_44444_32233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9055 a_2672_8585# a_1757_8213# a_2325_8181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X9056 a_4634_32182# a_4075_31591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9057 VSS a_1586_50247# a_6651_51733# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9058 a_10677_41831# a_10985_42044# a_10651_42035# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X9059 VSS pmat.row_n[12] a_25494_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X906 a_5351_60663# a_3866_57399# a_5518_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9060 a_47278_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9061 a_20170_23548# a_18546_23546# a_20078_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9062 a_40554_61190# pmat.rowon_n[5] a_40158_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9063 a_20811_41271# a_19689_41317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9064 a_28602_56492# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9065 a_8497_76457# a_2149_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9066 a_4349_62313# a_4509_62037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9067 a_23486_71230# pmat.rowon_n[15] a_23090_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9068 a_33222_22544# a_18546_22542# a_33130_22950# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9069 a_4699_28701# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X907 a_49686_10464# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9070 VDD nmat.rowon_n[15] a_34134_8894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9071 a_29206_12504# a_18546_12502# a_29114_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9072 a_51202_18934# pmat.row_n[10] a_51694_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9073 VSS VDD a_51598_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9074 vcm a_18162_19532# a_38242_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9075 a_45178_20942# a_18162_20536# a_45270_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9076 a_48282_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9077 a_19086_34343# a_19565_35279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9078 a_41254_59142# a_18546_59184# a_41162_59142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9079 a_5829_9615# a_5768_9527# a_5510_9615# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=4.7125e+11p ps=4.05e+06u w=650000u l=150000u
X908 a_23479_39095# a_22357_39141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9080 a_1959_10615# a_1979_11254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9081 a_11737_72943# a_11358_73309# a_11665_72943# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X9082 a_14471_27497# a_11337_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9083 a_40554_8854# nmat.rowon_n[15] a_40158_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9084 a_37542_18894# nmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9085 a_38759_31375# a_38851_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X9086 a_24270_49783# a_21371_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9087 VSS a_10864_68565# a_10740_68841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9088 a_44570_60186# pmat.rowon_n[4] a_44174_60146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9089 a_44570_19898# nmat.rowon_n[4] a_44174_19938# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X909 VDD a_40349_40726# a_40532_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9090 a_11322_72105# a_11019_71543# a_11014_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9091 VSS pmat.row_n[8] a_41558_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9092 a_27502_70226# pmat.rowon_n[14] a_27106_70186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9093 a_2847_41151# a_2411_33749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9094 a_7467_63303# a_7131_64822# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9095 VDD nmat.sample_n a_18162_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X9096 VDD a_4583_68021# a_4298_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9097 a_42065_50345# a_22199_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X9098 a_6872_8725# a_1586_8439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9099 a_22178_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X91 a_44174_13914# pmat.row_n[5] a_44666_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X910 a_26194_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9100 a_2203_41225# a_1757_40853# a_2107_41225# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X9101 a_45270_58138# a_18546_58180# a_45178_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9102 vcm a_18162_55166# a_42258_55126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9103 a_9234_31421# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9104 VDD a_5134_41909# a_5092_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9105 a_42166_59142# pmat.row_n[3] a_42658_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9106 a_43999_52521# a_16311_28327# a_43781_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9107 a_14365_22351# a_13798_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9108 a_4337_41935# a_4253_42729# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9109 a_4031_53034# a_4123_52789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X911 a_23090_60146# a_18162_60186# a_23182_60146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9110 a_22085_42902# a_22449_44219# a_23571_44265# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X9111 a_39387_41271# a_39781_41245# a_31793_41570# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X9112 a_5550_34319# a_4831_34561# a_4987_34293# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X9113 VSS pmat.row_n[9] a_27502_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9114 a_12132_58621# a_5535_57993# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9115 a_31518_57174# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9116 a_31518_15882# pmat.rowoff_n[7] a_31122_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9117 a_10388_51727# a_10245_51335# a_10045_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.15e+11p pd=2.83e+06u as=6.55e+11p ps=5.31e+06u w=1e+06u l=150000u
X9118 a_13896_8585# a_12815_8213# a_13549_8181# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9119 a_12061_26703# a_11713_26819# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X912 VSS pmat.row_n[12] a_47582_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9120 VDD a_14773_37218# a_13837_36893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X9121 a_37238_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9122 VSS a_6283_31591# a_22199_32149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9123 VDD VDD a_49194_72194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9124 a_42258_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9125 a_45648_31375# a_30663_50087# a_45345_31029# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X9126 vcm a_18162_24552# a_33222_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9127 VSS a_6651_44661# a_6800_44629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9128 vcm a_18162_66210# a_32218_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9129 a_43262_11500# a_18546_11498# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X913 a_40677_48437# a_33467_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9130 a_39666_30287# a_25575_31055# a_39497_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9131 vcm a_18162_56170# a_28202_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9132 a_9323_28879# a_4339_27804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9133 a_28704_29568# a_31399_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9134 a_22357_39141# a_20848_39429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X9135 a_3133_59709# a_2655_59317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9136 a_3026_16189# a_2411_16101# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9137 a_18162_8488# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X9138 VDD a_10927_43421# a_10985_44220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X9139 a_32618_58500# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X914 a_11203_62037# a_11713_64899# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X9140 a_28506_13874# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9141 a_24719_43957# a_11317_40188# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9142 VDD a_2021_11043# a_5746_11703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9143 VSS pmat.row_n[3] a_32522_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9144 a_34705_51959# a_41731_49525# a_41335_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9145 a_29206_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9146 a_19566_71552# pmat.col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9147 VDD pmat.rowoff_n[12] a_19074_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9148 a_34530_68218# pmat.rowon_n[12] a_34134_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9149 VSS a_9303_22351# a_10055_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X915 a_45921_42167# a_32405_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9150 vcm a_18162_16520# a_41254_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9151 VDD VDD a_23090_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9152 a_5232_72373# a_5257_69679# a_5361_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X9153 a_19074_61150# a_18162_61190# a_19166_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9154 VSS _1196_.B1 a_13354_2223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9155 a_38812_48829# a_38695_48634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9156 a_47582_67214# pmat.rowon_n[11] a_47186_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9157 VSS pmat.row_n[8] a_44570_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9158 a_5423_69367# a_2419_53351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9159 a_38150_23954# pmat.row_n[15] a_38642_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X916 a_26498_70226# pmat.col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9160 a_38150_19938# a_18162_19532# a_38242_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9161 a_2461_45565# a_2417_45173# a_2295_45577# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X9162 a_42658_21508# nmat.col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9163 a_10441_21263# a_10071_17999# a_10621_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9164 a_6412_8725# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9165 a_42258_17524# a_18546_17522# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9166 a_45178_65166# a_18162_65206# a_45270_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9167 a_10773_12559# comp_latch VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9168 VDD a_2149_45717# a_2093_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9169 a_37542_59182# pmat.rowon_n[3] a_37146_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X917 VDD a_10291_77269# a_10239_77295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9170 a_12709_19631# a_9528_20407# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9171 a_33869_31599# a_33331_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9172 VDD nmat.rowon_n[7] a_35138_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9173 a_7023_27907# a_7140_27805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9174 VDD a_10071_17999# a_10339_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X9175 vcm a_18162_17524# a_27198_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9176 a_21478_64202# pmat.rowon_n[8] a_21082_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9177 a_31165_28879# a_13641_23439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X9178 VSS a_23823_47679# a_23757_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X9179 a_31214_15516# a_18546_15514# a_31122_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X918 a_2648_29397# a_5547_14735# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X9180 VDD pmat.rowoff_n[7] a_48190_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9181 VSS a_13641_23439# a_31217_29429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9182 VDD a_29217_41570# a_28281_41245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X9183 VDD a_28969_27765# nmat.col[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9184 a_43170_13914# a_18162_13508# a_43262_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9185 pmat.col_n[31] a_11067_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9186 VSS a_45019_38645# a_44888_33205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9187 a_22178_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9188 a_22541_44581# a_21032_44007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X9189 a_36142_67174# a_18162_67214# a_36234_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X919 a_9493_66415# a_9405_66627# a_8891_66964# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9190 VSS VDD a_38546_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9191 a_31122_55126# VDD a_31614_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9192 a_22482_72234# pmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9193 a_14289_14441# a_10239_14183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9194 a_5741_38127# a_5687_38279# a_5659_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9195 a_24857_50959# a_15667_27239# pmat.col[5] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9196 a_49194_66170# a_18162_66210# a_49286_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9197 a_24847_43983# a_11317_40188# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9198 vcm a_18162_71230# a_40250_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9199 vcm a_18162_11500# a_32218_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X92 VDD a_10883_3303# a_13459_4943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.19e+12p ps=1.038e+07u w=1e+06u l=150000u M=2
X920 a_2769_22357# a_2603_22357# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9200 a_2215_8207# a_2199_13887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X9201 a_19166_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9202 a_35534_71230# pmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9203 a_49686_11468# nmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9204 a_39246_64162# a_18546_64204# a_39154_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9205 a_44266_7484# a_18546_7482# a_44174_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9206 a_40650_24520# nmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9207 VSS a_33423_47695# a_33519_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9208 VDD a_10883_3303# a_30558_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X9209 a_39646_68540# pmat.col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X921 a_31504_46831# a_29076_48695# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=0p ps=0u w=650000u l=150000u M=2
X9210 a_33130_24958# a_18162_24552# a_33222_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9211 VDD pmat.rowon_n[10] a_43170_66170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9212 a_9941_32509# a_9231_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9213 a_28639_47081# a_11067_49871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9214 a_31518_10862# nmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9215 VDD a_4955_40277# a_6733_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9216 a_5232_72373# a_5521_72373# a_5455_72719# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X9217 pmat.col_n[4] _1192_.A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9218 a_43262_56130# a_18546_56172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9219 a_37892_32509# a_5179_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X922 vcm a_18162_8488# a_25190_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9220 a_26194_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9221 vcm a_18162_9492# a_25190_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9222 vcm a_18162_70226# a_44266_70186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9223 VSS a_17996_36391# a_17959_36649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X9224 VDD nmat.rowon_n[12] a_26102_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9225 VDD a_2315_44124# a_4525_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9226 a_20051_30511# a_19605_30511# a_19955_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X9227 a_41162_20942# pmat.row_n[12] a_41654_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9228 a_36637_27497# a_34204_27765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X9229 a_41162_16926# a_18162_16520# a_41254_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X923 a_24094_23954# a_18162_23548# a_24186_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9230 VDD pmat.rowon_n[9] a_47186_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9231 a_44666_62516# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9232 vcm a_18162_59182# a_30210_59142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9233 a_29510_62194# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9234 a_41654_9460# nmat.col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9235 a_31122_72194# a_18162_72234# a_31214_72194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9236 VSS pmat.row_n[4] a_33526_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9237 a_34530_21906# nmat.rowon_n[2] a_34134_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9238 VSS a_4703_24527# a_7847_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9239 VSS pmat.row_n[11] a_33526_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X924 VDD a_43965_27221# nmat.col_n[23] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9240 a_30514_16886# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9241 a_21174_70186# a_18546_70228# a_21082_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9242 VDD pmat.rowon_n[1] a_37146_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9243 a_4601_35727# a_4307_35639# a_4517_35727# VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9244 a_18947_49811# a_19283_49783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X9245 a_9525_58255# a_9577_58229# a_5535_57993# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X9246 a_47582_20902# pmat.rowoff_n[12] a_47186_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9247 a_8289_46607# a_8079_46519# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9248 VDD nmat.rowon_n[14] a_51202_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9249 a_5721_8527# a_5558_9527# a_3663_9269# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X925 VDD pmat.rowon_n[9] a_34134_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9250 VDD pmat.rowon_n[6] a_21082_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9251 a_21082_64162# a_18162_64202# a_21174_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9252 a_42562_69222# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9253 VSS a_34553_42658# a_33617_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X9254 a_24869_49257# a_18823_50247# a_24773_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9255 vcm a_18162_58178# a_34226_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9256 VDD nmat.rowon_n[14] a_27106_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9257 a_37542_12870# pmat.rowoff_n[4] a_37146_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9258 VDD a_1761_4399# a_2025_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9259 a_2464_72221# a_2250_72221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X926 VDD a_2744_25223# a_2191_24501# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9260 VSS a_39505_38780# a_39197_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9261 a_22086_70186# pmat.row_n[14] a_22578_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9262 a_43170_58138# a_18162_58178# a_43262_58138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9263 VDD nmat.rowon_n[9] a_24094_14918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9264 vcm a_18162_21540# a_39246_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9265 a_2215_63695# a_1923_61759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9266 a_7645_17455# a_3305_15823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9267 a_32405_32463# a_9963_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9268 a_14369_21807# a_3305_15823# a_14005_22589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9269 a_5411_12167# a_5173_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X927 VDD nmat.rowon_n[13] a_26102_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9270 a_46578_68218# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9271 a_12267_38870# a_12237_38772# a_12195_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9272 a_43170_17930# pmat.row_n[9] a_43662_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9273 VDD a_10873_40693# a_11285_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9274 a_32126_11906# a_18162_11500# a_32218_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9275 a_18484_29967# a_12851_28853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X9276 VDD nmat.rowon_n[5] a_50198_18934# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9277 a_7477_31029# a_7259_31433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9278 ANTENNA_fanout52_A.DIODE pmat.sw VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X9279 VDD a_47207_35951# a_47035_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X928 a_41558_58178# pmat.rowon_n[2] a_41162_58138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9280 a_3175_72641# a_1674_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9281 a_8511_10422# comp_latch a_8511_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X9282 a_13913_65161# a_12723_64789# a_13804_65161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X9283 a_25590_10464# nmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9284 a_10071_17999# a_9820_18115# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9285 a_36538_18894# nmat.rowon_n[5] a_36142_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9286 VSS pmat.row_n[2] a_40554_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9287 VSS a_47915_46506# nmat.col[31] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9288 a_25327_28992# a_22307_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X9289 VSS pmat.row_n[12] a_23486_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X929 a_17619_43439# a_17442_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9290 a_49590_59182# pmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9291 a_11009_55785# a_10955_55687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9292 a_29206_20536# a_18546_20534# a_29114_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9293 a_20474_65206# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9294 a_2834_27791# a_1757_27797# a_2672_28169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9295 a_25098_9898# a_18162_9492# a_25190_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9296 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9297 a_51202_69182# a_18162_69222# a_51294_69182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9298 a_9510_10166# a_1717_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9299 a_14249_49525# a_6467_29415# a_14385_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X93 a_29510_66210# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X930 a_36142_9898# a_18162_9492# a_36234_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9300 vcm a_18162_69222# a_37238_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9301 a_11837_68591# a_11559_68619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X9302 a_47186_16926# pmat.row_n[8] a_47678_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9303 a_49590_8854# nmat.rowon_n[15] a_49194_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9304 a_41254_67174# a_18546_67216# a_41162_67174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9305 a_33986_47695# a_14887_46377# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X9306 a_33526_64202# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9307 a_17478_46805# a_16800_47213# a_17786_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9308 a_37238_57134# a_18546_57176# a_37146_57134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9309 VDD a_45529_51157# pmat.col_n[26] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X931 a_7461_19087# a_3688_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9310 VSS a_32957_30287# a_33607_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9311 VDD a_11883_62063# a_12079_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X9312 a_45705_33551# a_30663_50087# a_44888_33205# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9313 a_20221_40835# a_33765_40229# a_34828_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9314 a_38242_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9315 VDD pmat.rowon_n[3] a_41162_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9316 VSS pmat.row_n[6] a_37542_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9317 VSS a_2847_16127# a_2781_16201# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X9318 VSS pmat.row_n[3] a_26498_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9319 a_23486_56170# pmat.col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X932 a_13290_50095# a_11067_49871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9320 a_36380_34191# a_36203_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9321 a_20570_61512# pmat.col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9322 a_30514_57174# pmat.rowon_n[1] a_30118_57134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9323 a_24586_16488# nmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9324 VDD a_7079_40277# a_4955_40277# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X9325 a_7521_19631# a_6821_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9326 a_10873_38517# a_30771_39425# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X9327 VSS a_9963_13967# nmat.rowoff_n[9] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9328 vcm a_18162_63198# a_42258_63158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9329 a_27509_44219# a_26552_43781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X933 VDD pmat.rowon_n[8] a_47186_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9330 a_42166_67174# pmat.row_n[11] a_42658_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9331 a_1644_57685# a_1591_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9332 a_34883_52047# a_13091_28327# pmat.col[14] VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X9333 VSS a_35186_47375# a_43315_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9334 VDD a_25575_31055# a_38913_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9335 a_6087_67655# a_2879_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X9336 a_36142_7890# VDD a_36634_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9337 VSS a_1586_8439# a_2327_11477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9338 VSS a_4220_62037# a_2944_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X9339 a_36801_42405# a_36345_42567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X934 a_44666_61512# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9340 a_11193_43222# a_11021_43011# a_10979_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9341 result_out[7] a_1644_64213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9342 a_27502_55166# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9343 a_46674_7452# nmat.col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9344 a_42562_7850# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9345 VSS a_8851_63669# a_8782_63695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X9346 a_42562_22910# nmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9347 a_39154_21946# a_18162_21540# a_39246_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9348 a_36234_18528# a_18546_18526# a_36142_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9349 VSS a_18751_53034# pmat.rowoff_n[1] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X935 a_15048_36165# a_13985_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9350 vcm a_18162_64202# a_28202_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9351 a_28110_68178# pmat.row_n[12] a_28602_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9352 a_32218_62154# a_18546_62196# a_32126_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9353 a_6817_21807# a_6469_21813# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9354 a_32618_66532# pmat.col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9355 a_49286_17524# a_18546_17522# a_49194_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9356 VSS pmat.row_n[9] a_35534_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9357 pmat.col[29] a_47764_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9358 VSS VDD a_28506_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9359 a_32126_56130# a_18162_56170# a_32218_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X936 VSS pmat.row_n[4] a_20474_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9360 a_11501_10927# a_11167_11177# a_11417_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X9361 a_5510_9615# a_5654_9527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9362 a_46578_21906# nmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9363 a_4492_32375# a_4707_32156# a_4634_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9364 a_13259_35561# a_13653_35516# a_13319_35507# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X9365 vcm a_18162_24552# a_41254_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9366 a_12267_38543# a_12013_38870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9367 a_33526_9858# nmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9368 a_49194_57134# pmat.row_n[1] a_49686_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9369 vcm a_18162_14512# a_37238_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X937 a_34226_19532# a_18546_19530# a_34134_19938# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9370 a_9219_27497# a_4068_25615# a_9137_27253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9371 a_22459_48463# a_22015_48579# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9372 vcm a_18162_56170# a_36234_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9373 VSS a_38627_50613# a_38575_50639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9374 VSS VDD a_44570_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9375 VSS a_40949_48437# a_40707_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9376 VSS a_33467_46261# a_32827_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9377 a_40650_58500# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9378 a_37680_37479# a_36617_37691# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X9379 a_33130_62154# pmat.row_n[6] a_33622_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X938 VSS pmat.row_n[11] a_20474_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9380 a_36538_13874# nmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9381 VSS a_21037_43658# a_12228_40693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9382 a_34797_51727# a_34705_51959# pmat.col[14] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9383 a_18546_67216# pmat.sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X9384 a_50290_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9385 VSS a_12217_66389# a_12152_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.1125e+11p ps=1.95e+06u w=650000u l=150000u
X9386 VDD a_9919_51959# a_9827_53379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.85e+11p ps=2.57e+06u w=1e+06u l=150000u
X9387 a_2375_63316# a_2467_63125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X9388 VSS pmat.row_n[3] a_40554_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9389 a_19470_23914# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X939 a_46274_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9390 VSS a_13688_47893# a_14000_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9391 a_34887_35831# a_33765_35877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9392 a_49590_12870# nmat.col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9393 VSS pmat.row_n[13] a_23486_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9394 a_26594_57496# pmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9395 a_21478_72234# VDD a_21082_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9396 VDD VSS a_30118_55126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9397 a_28245_35877# a_27789_36039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X9398 a_31214_23548# a_18546_23546# a_31122_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9399 a_51598_61190# pmat.rowon_n[5] a_51202_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X94 VSS pmat.row_n[8] a_33526_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X940 a_29510_61190# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9400 a_25393_43493# a_24937_43655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X9401 a_27198_13508# a_18546_13506# a_27106_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9402 a_10609_28995# a_9741_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9403 VDD ANTENNA__1187__B1.DIODE a_14289_5737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9404 VSS a_79085_39738# a_78898_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9405 a_17012_47349# a_14653_53458# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X9406 a_45370_48169# a_30111_47911# a_45284_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X9407 VDD a_38711_37683# a_39505_38780# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=1.42e+06u
X9408 a_37837_29199# a_37795_29111# a_28812_29575# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X9409 pmat.en_bit_n[0] a_12461_29673# a_18484_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X941 VDD a_10991_68591# a_12629_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X9410 VDD a_40677_48437# a_11711_50959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X9411 a_11987_24847# a_10959_23983# a_12075_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9412 a_29510_15882# pmat.rowoff_n[7] a_29114_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9413 VSS pmat.row_n[4] a_26498_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9414 VSS pmat.row_n[7] a_38546_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9415 a_20474_9858# nmat.rowon_n[14] a_20078_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9416 a_19439_27497# a_6829_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X9417 a_30514_10862# nmat.rowon_n[13] a_30118_10902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9418 a_48586_18894# nmat.col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9419 VDD a_4339_27804# a_11251_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X942 a_34530_20902# pmat.rowoff_n[12] a_34134_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9420 a_4254_7351# a_3663_9269# a_4333_7913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9421 a_39246_72194# a_18546_72236# a_39154_72194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9422 vcm a_18162_61190# a_31214_61150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9423 VDD ANTENNA__1395__A2.DIODE a_47775_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9424 a_36634_22512# nmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9425 VSS a_9075_28023# a_10791_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9426 a_46753_41935# a_40837_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X9427 VSS a_11021_43011# a_20811_42359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X9428 a_31339_31787# a_37827_30793# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X9429 VDD pmat.rowoff_n[12] a_40158_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X943 a_31122_71190# a_18162_71230# a_31214_71190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9430 VSS a_2972_9991# a_4085_7663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9431 a_38812_48829# a_38695_48634# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9432 a_9301_69679# a_9135_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9433 a_43262_64162# a_18546_64204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9434 a_40158_61150# a_18162_61190# a_40250_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9435 a_6978_58799# a_5462_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9436 VSS a_6244_71829# a_5521_72373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X9437 a_12461_53903# a_12003_52815# a_11902_56775# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9438 a_23090_71190# a_18162_71230# a_23182_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9439 a_28506_62194# pmat.rowon_n[6] a_28110_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X944 a_30514_15882# nmat.col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9440 VSS a_5651_66975# a_8599_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9441 a_6520_37039# a_6403_37252# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9442 a_11711_60751# a_10878_58487# a_11797_60431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9443 VSS a_1923_31743# a_4853_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9444 VDD a_8765_64757# a_8655_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9445 a_41162_24958# a_18162_24552# a_41254_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9446 VSS a_2944_67752# a_2882_67869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X9447 VSS a_7808_61493# a_7563_63303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X9448 a_44666_70548# pmat.col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9449 a_37146_14918# a_18162_14512# a_37238_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X945 VSS pmat.row_n[10] a_33526_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9450 VSS a_33617_42333# a_33309_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9451 VDD a_14691_29575# a_14471_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9452 vcm a_18162_67214# a_30210_67174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9453 a_41254_12504# a_18546_12502# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9454 a_35230_9492# a_18546_9490# a_35138_9898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9455 VSS a_11067_30287# a_22083_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X9456 a_25315_28335# a_25325_29125# a_25143_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X9457 a_41558_69222# pmat.rowon_n[13] a_41162_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9458 a_44174_60146# a_18162_60186# a_44266_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9459 a_11547_48061# a_5363_33551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X946 VDD a_44763_34293# a_45107_34863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9460 a_30543_40721# cgen.dlycontrol4_in[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9461 a_27106_70186# a_18162_70226# a_27198_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9462 VSS pmat.row_n[15] a_20474_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9463 VSS a_12613_57141# a_12371_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9464 VDD nmat.rowon_n[12] a_34134_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9465 a_7140_27805# a_7888_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X9466 a_19470_64202# pmat.rowon_n[8] a_19074_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9467 vcm a_18162_12504# a_26194_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9468 a_27579_34967# a_24833_34191# a_27753_35073# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9469 a_3644_65871# a_3207_65845# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X947 VDD pmat.rowon_n[0] a_37146_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9470 VDD pmat.rowon_n[14] a_21082_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9471 a_30210_10496# a_18546_10494# a_30118_10902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9472 a_3325_26159# a_2847_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9473 VDD nmat.rowon_n[13] a_47186_10902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9474 a_38546_67214# pmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9475 a_14718_19631# a_10515_15055# a_14340_19783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9476 _1224_.X a_82863_64213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=8
X9477 a_21174_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9478 a_45574_68218# pmat.rowon_n[12] a_45178_68178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9479 VSS a_2467_35925# a_1895_36666# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X948 a_9161_12925# a_8782_12559# a_9089_12925# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9480 VSS pmat.row_n[9] a_42562_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9481 VDD a_13457_64757# a_13347_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9482 VDD clk_vcm vcm.sky130_fd_sc_hd__inv_1_4.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9483 a_45113_47375# a_33423_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9484 a_51598_15882# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9485 VSS a_37525_27221# nmat.col_n[17] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9486 VSS a_26041_36374# a_26331_36919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X9487 a_6316_8903# a_6412_8725# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9488 a_27249_31055# a_20616_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=0p ps=0u w=1e+06u l=150000u
X9489 a_18521_46837# a_18547_51565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X949 vcm a_18162_58178# a_21174_58138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9490 a_18162_13508# nmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X9491 VSS a_16083_50069# a_16219_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9492 a_38642_63520# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9493 a_8363_56457# a_8013_56085# a_8268_56445# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X9494 vcm a_18162_18528# a_25190_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9495 a_48586_59182# pmat.rowon_n[3] a_48190_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9496 VDD pmat.rowon_n[5] a_42166_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9497 VDD a_1858_25615# a_2511_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9498 a_3080_30333# a_2500_30345# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X9499 VDD nmat.rowon_n[7] a_46182_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X95 a_47678_55488# pmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X950 VDD a_9889_10681# a_9919_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9500 a_13645_59343# a_10239_14183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9501 a_24490_17890# nmat.col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9502 VDD a_1642_26935# a_1591_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9503 a_4037_69109# a_3508_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9504 VDD a_4737_21561# a_4767_21302# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9505 a_32957_30287# a_33011_29941# a_32969_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9506 VSS a_26891_28327# pmat.col_n[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.1125e+11p ps=1.95e+06u w=650000u l=150000u
X9507 VDD a_1739_47893# a_1941_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9508 a_50594_62194# pmat.col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9509 a_47186_67174# a_18162_67214# a_47278_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X951 VDD a_16890_36911# a_18999_35279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9510 VSS VDD a_49590_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9511 VSS a_29163_38545# a_29109_38571# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9512 a_13604_72765# a_6451_67655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9513 a_33526_72234# pmat.col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9514 a_18107_53034# a_18199_52789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X9515 a_14729_3311# a_10883_3303# nmat.col[12] VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X9516 a_37238_65166# a_18546_65208# a_37146_65166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9517 a_24186_8488# a_18546_8486# a_24094_8894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9518 a_37638_69544# pmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9519 VDD pmat.rowon_n[11] a_41162_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X952 a_18869_46831# a_18521_46837# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9520 a_35230_9492# a_18546_9490# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9521 VDD a_24719_43957# a_14773_43746# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9522 a_26102_10902# a_18162_10496# a_26194_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9523 a_12081_3855# a_9411_2215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9524 a_37146_59142# a_18162_59182# a_37238_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9525 a_51694_24520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9526 a_41254_57134# a_18546_57176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9527 a_32687_46607# a_9785_28879# a_33101_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9528 VDD pmat.rowon_n[6] a_19074_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9529 a_24186_67174# a_18546_67216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X953 VDD pmat.rowon_n[5] a_21082_61150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9530 a_26498_55166# VSS a_26102_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9531 a_37637_32149# a_37471_32149# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9532 a_41558_64202# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9533 a_41558_22910# nmat.rowon_n[1] a_41162_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9534 a_40041_27791# a_25879_31591# nmat.col_n[20] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9535 a_12153_74575# a_10697_75218# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9536 a_11041_36596# a_12267_36694# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9537 a_38150_65166# pmat.row_n[9] a_38642_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9538 cgen.dlycontrol1_in[3] a_1591_33231# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X9539 a_11145_17999# a_10975_17999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X954 a_25687_34743# a_24565_34789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9540 a_2629_69679# a_2250_70045# a_2557_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9541 a_2840_55509# a_3225_55509# a_2969_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X9542 VDD a_3960_19465# a_4135_19391# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9543 VDD a_10239_77295# a_10995_76207# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9544 a_27502_63198# pmat.col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9545 VDD a_11703_48156# a_11634_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9546 VSS a_20499_31274# a_9307_31068# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9547 VDD a_29051_39783# a_12345_39100# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X9548 a_22085_38550# a_22357_39141# a_23420_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9549 a_38546_20902# nmat.col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X955 a_23063_36885# a_14712_37429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9550 _1187_.A2 a_46947_39215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=8
X9551 a_45670_15484# nmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9552 a_42166_12910# pmat.row_n[4] a_42658_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9553 a_45574_21906# nmat.rowon_n[2] a_45178_21946# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9554 VSS a_10873_39605# a_10817_39958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9555 vcm a_18162_72234# a_28202_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9556 VDD pmat.rowon_n[1] a_48190_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9557 a_32218_70186# a_18546_70228# a_32126_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9558 a_25098_22950# pmat.row_n[14] a_25590_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9559 VDD a_2931_40277# a_1895_41018# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X956 a_48682_60508# pmat.col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9560 a_18162_58178# pmat.sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X9561 VDD pmat.rowoff_n[15] a_32126_23954# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9562 a_2464_65693# a_2250_65693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9563 a_41443_28879# a_41192_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X9564 a_32126_64162# a_18162_64202# a_32218_64162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9565 a_35534_13874# nmat.rowon_n[10] a_35138_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9566 a_27443_32463# a_27498_32117# a_27443_32143# VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9567 VSS a_39981_37462# a_39045_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X9568 VSS a_33341_38780# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X9569 VDD a_3576_17143# a_5271_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X957 a_10815_55785# a_10497_54697# a_11009_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9570 VDD pmat.rowoff_n[7] a_22086_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9571 a_48586_12870# pmat.rowoff_n[4] a_48190_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9572 VDD a_5331_28309# a_5318_28701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9573 a_46182_11906# pmat.row_n[3] a_46674_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9574 vcm a_18162_64202# a_36234_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9575 a_18660_47607# a_12263_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9576 a_36142_68178# pmat.row_n[12] a_36634_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9577 a_40250_62154# a_18546_62196# a_40158_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9578 a_29114_21946# pmat.row_n[13] a_29606_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9579 a_40650_66532# pmat.col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X958 a_28975_40871# cgen.dlycontrol3_in[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9580 a_29114_17930# a_18162_17524# a_29206_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9581 a_33130_70186# pmat.row_n[14] a_33622_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9582 VDD pmat.rowon_n[3] a_39154_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9583 a_32468_51433# a_28915_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9584 a_33765_38053# a_30431_37683# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
X9585 a_33222_15516# a_18546_15514# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9586 a_30118_12910# a_18162_12504# a_30210_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9587 VSS a_17996_35303# a_17959_35561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X9588 VDD a_2389_45859# a_5029_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9589 VSS pmat.row_n[1] a_43566_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X959 vcm a_18162_57174# a_34226_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9590 a_7847_20719# a_7048_23277# a_7935_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.665e+11p ps=2.12e+06u w=650000u l=150000u
X9591 a_18162_70226# pmat.sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X9592 VDD a_36946_34191# a_37823_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9593 a_9368_9991# a_9583_10121# a_9510_10166# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9594 a_10055_31591# a_18947_49811# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X9595 a_2163_53057# a_1586_50247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9596 a_12150_60137# a_10049_60663# a_11842_59887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9597 a_19074_13914# pmat.row_n[5] a_19566_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9598 a_23582_11468# nmat.col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9599 nmat.rowoff_n[13] a_12447_16143# a_14649_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X96 VSS a_10927_37981# a_10867_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X960 a_2203_50095# a_1757_50095# a_2107_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X9600 a_41162_62154# pmat.row_n[6] a_41654_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9601 a_27198_21540# a_18546_21538# a_27106_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9602 a_5101_76751# a_5047_76983# a_4123_76181# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X9603 VSS pmat.row_n[2] a_51598_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9604 a_29510_9858# nmat.rowon_n[14] a_29114_9898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9605 a_2629_61885# a_2250_61519# a_2557_61885# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9606 a_12255_44535# a_11133_44581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9607 a_7489_17455# a_4976_16091# a_7407_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9608 VSS pmat.row_n[12] a_34530_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9609 a_44963_45199# a_31675_47695# a_44855_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X961 VDD a_5967_5461# a_5558_9527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9610 vcm a_18162_69222# a_48282_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9611 a_10497_54697# a_10117_54697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X9612 a_45178_19938# pmat.row_n[11] a_45670_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9613 VSS a_30431_37683# a_30371_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X9614 a_35230_13508# a_18546_13506# a_35138_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9615 a_49286_70186# a_18546_70228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9616 VSS a_2375_18708# a_1895_18170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9617 VDD a_10781_42869# a_11193_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9618 a_8268_56445# a_4843_54826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9619 a_42562_71230# pmat.rowon_n[15] a_42166_71190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X962 a_14923_34473# a_13529_34951# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X9620 a_40158_8894# pmat.row_n[0] a_40650_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9621 a_27106_63158# pmat.row_n[7] a_27598_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9622 VDD a_3866_57399# a_5085_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X9623 VSS a_10223_26703# a_13073_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9624 a_31614_61512# pmat.col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9625 a_48282_12504# a_18546_12502# a_48190_12910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9626 a_4333_30511# a_4167_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9627 a_19283_49783# a_30189_48437# a_30219_48783# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u M=2
X9628 a_11117_8779# a_11051_8903# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9629 a_39246_62154# a_18546_62196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X963 a_34530_14878# nmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9630 VSS a_79085_40202# a_78898_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9631 a_22578_19500# nmat.col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9632 VDD pmat.rowon_n[0] a_24094_56130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9633 VDD a_34924_37253# a_34828_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9634 VDD a_24937_41479# a_25260_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9635 a_22482_8854# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9636 a_26594_8456# nmat.col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9637 a_40554_23914# nmat.col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9638 a_1757_38677# a_1591_38677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9639 a_37146_22950# a_18162_22544# a_37238_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X964 a_11444_55535# a_10815_55785# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9640 VSS a_14113_43132# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X9641 VDD a_11067_16359# a_14287_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9642 VSS a_13795_10687# a_13729_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X9643 a_41254_20536# a_18546_20534# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9644 a_8491_23555# a_2683_22089# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9645 a_29206_68178# a_18546_68220# a_29114_68178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9646 VSS pmat.row_n[0] a_32522_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9647 VSS a_4859_31274# a_4471_30724# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9648 VSS a_18277_37620# a_14712_37429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9649 a_47278_18528# a_18546_18526# a_47186_18934# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X965 a_16197_40517# a_16171_40157# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9650 VSS a_17740_31287# a_16635_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9651 a_19470_72234# VDD a_19074_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9652 vcm a_18162_20536# a_26194_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9653 a_36345_42567# a_36617_43131# a_37680_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9654 a_49590_61190# pmat.rowon_n[5] a_49194_61150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9655 a_30118_57134# a_18162_57174# a_30210_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9656 a_8399_18115# a_7809_17705# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X9657 a_10299_51433# a_9463_50877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9658 VDD a_40837_46261# a_44371_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X9659 a_31701_37462# a_30913_38053# a_32035_38007# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X966 a_25590_72556# pmat.col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9660 VSS pmat.row_n[9] a_46578_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9661 a_50594_15882# pmat.rowoff_n[7] a_50198_15922# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9662 nmat.col_n[10] a_14458_5487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9663 a_11476_36189# a_11225_35836# a_11255_35862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X9664 a_8765_76725# a_8547_77129# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X9665 a_8732_10749# a_8481_10396# a_8511_10422# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9666 a_15574_48169# a_6467_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9667 a_14287_50345# a_14249_49525# a_14369_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X9668 a_27198_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9669 a_2676_29941# a_1923_31743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X967 vcm a_18162_20536# a_39246_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9670 VSS a_6602_72007# a_6244_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X9671 a_7732_52105# a_6651_51733# a_7385_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9672 vcm a_18162_66210# a_51294_66170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9673 vcm a_18162_14512# a_48282_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9674 a_3339_70759# a_2389_45859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X9675 vcm a_18162_56170# a_47278_56130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9676 a_45471_27497# a_15667_27239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9677 VSS a_22725_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X9678 a_51694_58500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9679 a_23486_17890# nmat.rowon_n[6] a_23090_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X968 a_43170_57134# a_18162_57174# a_43262_57134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9680 a_47582_13874# nmat.col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9681 a_21082_16926# pmat.row_n[8] a_21574_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9682 nmat.col[5] a_10883_3303# a_23846_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X9683 VSS pmat.row_n[3] a_51598_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9684 a_48282_10496# a_18546_10494# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9685 a_38642_71552# pmat.col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9686 a_34134_15922# pmat.row_n[7] a_34626_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9687 vcm a_18162_8488# a_47278_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9688 VSS pmat.row_n[13] a_34530_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9689 a_11415_14557# a_10791_14191# a_11307_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X969 VSS a_4266_63303# a_4061_63303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9690 a_18546_13506# nmat.sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X9691 a_13211_26703# a_13145_26935# a_13103_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X9692 a_24186_56130# a_18546_56172# a_24094_56130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9693 a_21371_50087# a_45238_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9694 a_14646_19881# a_9963_13967# a_14340_19783# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9695 a_27502_16886# nmat.rowon_n[7] a_27106_16926# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9696 VSS pmat.row_n[5] a_24490_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9697 a_1644_68565# a_1823_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9698 a_5633_22057# nmat.sw a_5537_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9699 VSS pmat.row_n[7] a_49590_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 a_5325_9269# a_5654_9527# a_5612_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=4.2e+11p ps=2.84e+06u w=1e+06u l=150000u
X970 a_3951_77055# a_3776_77129# a_4130_77117# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9700 a_39550_69222# pmat.rowon_n[13] a_39154_69182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9701 VSS pmat.row_n[10] a_36538_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9702 vcm a_18162_17524# a_46274_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9703 a_40554_64202# pmat.rowon_n[8] a_40158_64162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9704 a_28202_55126# a_18546_55168# a_28110_55126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9705 a_8951_27907# a_4516_21531# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X9706 a_28602_59504# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9707 a_50290_15516# a_18546_15514# a_50198_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9708 a_11225_35836# a_11071_36694# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9709 a_11860_56873# a_6787_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X971 VSS a_2847_50069# a_2983_48071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9710 VSS a_11113_40835# a_37739_42089# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X9711 a_45866_38279# a_45625_36495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X9712 a_41254_65166# a_18546_65208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9713 a_47678_22512# nmat.col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9714 a_47084_37039# a_43533_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=0p ps=0u w=650000u l=150000u
X9715 a_2012_33775# a_1775_35113# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9716 a_37680_36391# a_36617_36603# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X9717 a_2250_72221# a_2163_71997# a_1846_72107# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X9718 VDD pmat.rowon_n[14] a_19074_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9719 a_38557_48469# a_38391_48469# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X972 VDD a_82818_69135# _1154_.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u M=16
X9720 a_37238_55126# a_18546_55168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9721 VDD pmat.rowoff_n[12] a_51202_20942# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9722 a_26498_63198# pmat.rowon_n[7] a_26102_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9723 a_41558_72234# pmat.col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9724 a_38927_42359# a_38737_41814# VSS VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X9725 a_44789_39215# a_45019_38645# ANTENNA__1395__A2.DIODE VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9726 a_23182_17524# a_18546_17522# a_23090_17930# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9727 a_10675_76029# a_10239_77295# a_10579_76029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9728 a_37638_14480# nmat.col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9729 a_4070_47375# a_2935_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X973 a_2319_65564# a_2124_65595# a_2629_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X9730 vcm a_18162_11500# a_51294_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9731 a_38242_18528# a_18546_18526# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9732 VDD pmat.rowoff_n[4] a_41162_12910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9733 a_5553_62607# a_5497_62839# a_5065_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9734 a_48190_14918# a_18162_14512# a_48282_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9735 a_20695_30485# a_1858_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9736 VDD a_2847_26133# a_2834_26525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9737 a_34530_55166# pmat.en_bit_n[1] a_34134_55126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9738 a_12687_18377# a_12337_18005# a_12592_18365# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X9739 VDD a_1586_33927# a_5823_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X974 VDD pmat.rowon_n[4] a_25098_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9740 a_4491_53511# a_4587_53505# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X9741 vcm a_18162_13508# a_24186_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9742 a_45270_66170# a_18546_66212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9743 a_38150_10902# pmat.row_n[2] a_38642_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9744 VSS pmat.row_n[15] a_31518_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9745 VDD nmat.rowon_n[12] a_45178_11906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9746 VDD a_40837_46261# a_42683_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9747 VDD pmat.rowon_n[12] a_35138_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9748 a_9099_47753# a_8583_47381# a_9004_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X9749 a_9685_74281# a_9831_74183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u
X975 a_5173_45743# a_4313_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9750 a_2325_8181# a_2107_8585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X9751 VDD a_17336_43439# a_17442_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9752 VDD nmat.rowon_n[2] a_28110_21946# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9753 a_83092_15055# ANTENNA__1183__B1.DIODE a_82787_14709# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X9754 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9755 a_3026_43389# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9756 a_28110_62154# a_18162_62194# a_28202_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9757 a_4181_37289# a_4127_37013# a_2467_35925# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9758 a_22015_28995# a_19405_28853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9759 VSS a_20848_41605# a_20811_41271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X976 a_46578_67214# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9760 a_4123_76181# a_4951_76983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9761 a_2215_23439# a_1591_23445# a_2107_23817# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X9762 a_32218_60146# a_18546_60188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9763 VSS a_13357_37429# a_24895_37429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9764 vcm a_18162_72234# a_36234_72194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9765 a_38812_47741# a_38569_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9766 a_17842_27497# a_7840_27247# a_16965_27247# VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X9767 VSS a_20572_40517# a_20645_42044# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.69e+06u
X9768 a_40250_70186# a_18546_70228# a_40158_70186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9769 a_10989_72943# a_10954_73195# a_10751_72917# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X977 a_8569_60405# a_8841_60405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9770 a_3697_65103# a_3609_65015# a_2944_65576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9771 a_36234_60146# a_18546_60188# a_36142_60146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9772 vcm a_18162_71230# a_49286_71190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9773 VDD pmat.rowon_n[11] a_39154_67174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9774 a_9820_18115# a_9557_17705# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9775 a_36634_64524# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9776 VSS a_6559_33767# a_7109_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X9777 a_30118_20942# a_18162_20536# a_30210_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9778 a_33222_23548# a_18546_23546# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9779 vcm a_18162_19532# a_23182_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X978 a_17323_28111# _0467_ VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0725e+12p pd=1.11e+07u as=0p ps=0u w=650000u l=150000u M=2
X9780 VDD pmat.rowon_n[6] a_40158_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9781 a_29206_13508# a_18546_13506# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9782 VSS a_23815_28023# nmat.col[4] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9783 a_33130_9898# pmat.row_n[1] a_33622_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9784 VDD a_2939_45503# a_2389_45859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X9785 a_49686_63520# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9786 VSS a_35099_34191# a_35205_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9787 VSS pmat.row_n[6] a_25494_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9788 VSS a_4308_21495# a_4123_20693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9789 a_22482_18894# nmat.col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X979 nmat.en_bit_n[1] a_12437_28879# a_17748_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X9790 VDD a_1957_43567# a_11071_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9791 a_11547_48061# a_5363_33551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9792 a_5227_13077# a_4895_12559# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9793 a_11877_12565# a_11711_12565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9794 a_30403_40747# a_24833_40719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9795 a_6639_63927# a_6568_59887# a_6984_64015# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X9796 a_39550_22910# nmat.rowon_n[1] a_39154_22950# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9797 a_35534_17890# nmat.col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9798 VSS a_7109_29423# a_47120_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9799 a_41162_70186# pmat.row_n[14] a_41654_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X98 a_27106_23954# pmat.row_n[15] a_27598_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X980 a_5248_30511# a_4333_30511# a_4901_30753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X9800 VSS a_22787_42325# a_15049_42902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9801 a_26194_71190# a_18546_71232# a_26102_71190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9802 VSS a_7048_23277# a_6800_22869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9803 a_37146_60146# pmat.row_n[4] a_37638_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9804 a_45178_68178# a_18162_68218# a_45270_68178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9805 a_27181_30511# a_20616_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X9806 a_30210_58138# a_18546_58180# a_30118_58138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9807 VDD pmat.rowon_n[7] a_26102_63158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9808 VDD a_5331_28309# a_3351_27249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9809 a_51202_11906# a_18162_11500# a_51294_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X981 a_4553_28089# a_2564_21959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9810 a_8291_23983# a_7847_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X9811 VSS a_5363_33551# a_14287_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9812 VDD a_17625_42902# a_18176_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9813 a_49194_8894# pmat.row_n[0] a_49686_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9814 VSS a_1674_57711# a_11711_58261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9815 a_35230_21540# a_18546_21538# a_35138_21946# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9816 a_27106_71190# pmat.row_n[15] a_27598_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9817 a_48190_59142# a_18162_59182# a_48282_59142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9818 a_22178_68178# a_18546_68220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9819 a_4737_23957# a_2564_21959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X982 VSS a_29404_44869# a_29367_44535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X9820 a_9217_49007# a_7373_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X9821 VDD nmat.rowon_n[14] a_20078_9898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9822 a_48282_20536# a_18546_20534# a_48190_20942# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9823 VSS a_11927_27399# a_14691_27399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9824 a_45469_53135# _1179_.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9825 VDD a_35224_50613# pmat.col[16] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9826 a_5156_28335# a_4241_28335# a_4809_28577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9827 VDD a_44791_43541# a_44739_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9828 VDD a_30571_50959# a_36175_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9829 a_28901_48437# a_30999_48071# a_32030_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3e+11p ps=5.26e+06u w=1e+06u l=150000u M=2
X983 VSS pmat.row_n[9] a_50594_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9830 a_13055_10761# a_12539_10389# a_12960_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X9831 a_50198_21946# pmat.row_n[13] a_50690_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9832 a_5749_30265# a_4075_31591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9833 VDD a_7658_71543# a_9135_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9834 a_50198_17930# a_18162_17524# a_50290_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9835 VSS pmat.row_n[3] a_45574_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9836 a_42562_56170# pmat.col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9837 a_39154_18934# pmat.row_n[10] a_39646_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9838 VSS VDD a_39550_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9839 a_43662_16488# nmat.col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X984 VDD nmat.rowon_n[6] a_50198_17930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9840 a_40158_13914# pmat.row_n[5] a_40650_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9841 VSS pmat.row_n[13] a_28506_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9842 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9843 a_25494_66210# pmat.col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9844 VSS a_21371_50087# a_22199_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9845 VSS a_3866_57399# a_5633_71631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9846 a_19891_36919# a_18769_36965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9847 a_32522_67214# pmat.rowon_n[11] a_32126_67174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9848 a_23090_23954# pmat.row_n[15] a_23582_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9849 VDD a_2791_57703# a_4319_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X985 a_15299_28879# a_14943_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X9850 conversion_finished_out a_1644_77813# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9851 a_23090_19938# a_18162_19532# a_23182_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9852 a_7737_17705# a_3305_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9853 a_30118_65166# a_18162_65206# a_30210_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9854 a_12954_58255# a_11877_58261# a_12792_58633# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9855 VSS a_2499_13077# a_2199_13887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9856 a_6752_24527# a_3305_27791# a_6646_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
X9857 a_29206_58138# a_18546_58180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9858 a_42562_8854# nmat.rowon_n[15] a_42166_8894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9859 a_22482_59182# pmat.rowon_n[3] a_22086_59142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X986 VSS a_20184_46983# nmat.rowon_n[12] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9860 a_46578_55166# pmat.col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9861 a_7179_44905# a_4128_46983# a_7107_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9862 VSS a_2163_56765# a_2124_56891# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9863 a_46578_13874# nmat.rowon_n[10] a_46182_13914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9864 VDD nmat.rowon_n[7] a_20078_16926# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9865 a_7779_22583# a_9227_20291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9866 a_29510_65206# pmat.col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9867 a_10478_25045# a_9528_20407# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9868 VSS a_1959_12791# a_1959_12559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9869 a_29606_17492# nmat.col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X987 a_36538_59182# pmat.col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9870 a_7079_40277# a_6904_40303# a_7258_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9871 VDD a_2672_39049# a_2847_38975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9872 VDD a_11067_30287# a_40979_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.344e+11p ps=1.7e+06u w=640000u l=150000u
X9873 a_38581_47081# a_1781_9308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9874 VDD pmat.rowoff_n[7] a_33130_15922# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9875 a_27106_18934# a_18162_18528# a_27198_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9876 VDD a_29076_48695# a_31053_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X9877 vcm a_18162_64202# a_47278_64162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9878 a_47186_68178# pmat.row_n[12] a_47678_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9879 a_51294_62154# a_18546_62196# a_51202_62154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X988 a_13091_52047# a_41663_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X9880 VSS a_1591_16367# a_1739_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X9881 a_2012_18365# a_1895_18170# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9882 a_51694_66532# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9883 a_20173_30753# a_19955_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9884 a_46487_49871# a_30663_50087# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=0p ps=0u w=650000u l=150000u M=4
X9885 a_19470_57174# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9886 a_11773_39087# a_11507_39087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9887 VDD a_33719_44527# a_33825_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9888 a_14477_22057# a_4523_21276# a_14005_22589# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9889 VSS a_3325_43023# a_3993_44431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X989 a_8292_27023# a_6664_26159# a_8031_26703# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X9890 VDD a_2149_45717# a_5553_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9891 a_21082_67174# a_18162_67214# a_21174_67174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9892 VSS VDD a_23486_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9893 a_5184_42301# a_3983_41941# a_4984_41935# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.47e+11p ps=1.54e+06u w=420000u l=150000u
X9894 a_7253_15055# a_3576_17143# a_7169_15055# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9895 cgen.dlycontrol1_in[0] a_1591_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X9896 a_51202_56130# a_18162_56170# a_51294_56130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9897 a_35230_21540# a_18546_21538# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9898 a_34134_66170# a_18162_66210# a_34226_66170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9899 a_26272_37253# a_25209_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X99 a_27106_19938# a_18162_19532# a_27198_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X990 VDD a_23239_37217# a_23063_36885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9900 VDD a_45908_33749# a_44533_33749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X9901 a_37776_37479# a_36617_37691# a_37739_37737# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9902 a_24186_64162# a_18546_64204# a_24094_64162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9903 a_34626_11468# nmat.col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9904 a_2215_50461# a_1591_50095# a_2107_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X9905 a_24586_68540# pmat.col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9906 a_8765_64757# a_8547_65161# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9907 VSS a_2879_60975# a_2727_58470# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9908 a_44266_8488# a_18546_8486# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9909 VDD a_20848_36165# a_20752_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X991 a_44984_48783# a_44870_48437# a_21279_48999# VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X9910 VSS a_9963_13967# nmat.rowoff_n[10] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9911 VDD a_8175_63669# a_1823_66941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9912 a_45670_57496# pmat.col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9913 a_17417_49667# a_16800_47213# a_17322_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X9914 a_28202_63158# a_18546_63200# a_28110_63158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9915 vcm a_18162_60186# a_25190_60146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9916 a_40554_72234# VDD a_40158_72194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9917 a_28602_67536# pmat.col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9918 a_25098_64162# pmat.row_n[8] a_25590_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9919 a_13798_22351# a_13768_22325# a_13726_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X992 a_36538_17890# nmat.rowon_n[6] a_36142_17930# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9920 a_50290_23548# a_18546_23546# a_50198_23954# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9921 VDD pmat.rowon_n[9] a_32126_65166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9922 a_46274_13508# a_18546_13506# a_46182_13914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9923 VDD VDD a_25098_7890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9924 VSS VDD a_21478_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9925 vcm a_18162_10496# a_43262_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9926 a_2021_11043# a_3583_11775# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9927 VSS _1192_.A2 nmat.col[5] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9928 a_37238_63158# a_18546_63200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9929 VDD a_3484_58229# a_2944_59048# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X993 VSS pmat.row_n[1] a_40554_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9930 VSS pmat.row_n[4] a_45574_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9931 a_13457_64757# a_13239_65161# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9932 a_31518_7850# VDD a_31122_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9933 VDD a_1923_53055# a_2464_59165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9934 a_2307_45199# a_2411_43301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9935 VDD pmat.rowon_n[1] a_22086_57134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9936 VDD a_1923_61759# a_4028_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X9937 VSS pmat.row_n[14] a_28506_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9938 VSS a_2847_43327# a_2781_43401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X9939 a_37542_70226# pmat.col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X994 a_29051_37607# a_29159_37607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9940 vcm a_18162_22544# a_20170_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9941 VDD a_12557_32441# a_12587_32182# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9942 a_32522_20902# pmat.rowoff_n[12] a_32126_20942# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9943 a_19166_15516# a_18546_15514# a_19074_15922# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9944 a_9455_31421# a_9307_31068# a_9092_31287# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X9945 VSS a_28704_29568# a_43548_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9946 VSS a_5271_35407# a_5550_34319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9947 VSS a_5331_53511# a_4081_61127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9948 VDD a_15093_39638# a_15048_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9949 a_12066_3087# a_9411_2215# a_11980_3087# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X995 a_19470_69222# pmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9950 a_48190_22950# a_18162_22544# a_48282_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9951 a_22482_12870# pmat.rowoff_n[4] a_22086_12910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9952 a_34530_63198# pmat.rowon_n[7] a_34134_63158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9953 a_19074_55126# VDD a_19566_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9954 nmat.col_n[25] a_16311_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9955 a_45475_35520# a_44763_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X9956 vcm a_18162_21540# a_24186_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9957 a_42166_71190# a_18162_71230# a_42258_71190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9958 a_47582_62194# pmat.rowon_n[6] a_47186_62154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9959 a_7074_49007# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X996 VDD a_16083_50069# a_18675_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9960 VSS pmat.row_n[10] a_44570_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9961 a_47764_51433# _1194_.A2 a_47673_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X9962 a_23090_7890# a_18162_7484# a_23182_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9963 a_47207_35951# a_46934_35951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9964 a_6179_65479# a_2879_57487# a_6524_65327# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X9965 vcm a_18162_7484# a_36234_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9966 VDD a_14264_72777# a_14439_72703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9967 VSS a_46449_46261# a_45112_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9968 a_31518_68218# pmat.col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9969 VSS a_9749_19061# a_7693_22365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X997 a_1644_72917# a_1591_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9970 result_out[12] a_1644_71285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9971 VSS a_24719_36341# a_15049_36374# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9972 a_2012_50095# a_1895_50308# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9973 a_19470_10862# nmat.col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9974 a_3118_45565# a_2411_43301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9975 a_46274_7484# a_18546_7482# a_46182_7890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9976 a_4699_13647# a_4075_13653# a_4591_14025# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X9977 vcm a_18162_57174# a_45270_57134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9978 VDD a_22307_27791# a_24861_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9979 a_46182_70186# a_18162_70226# a_46274_70186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X998 VSS pmat.row_n[11] a_23486_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9980 a_12895_53359# a_12213_53359# a_12723_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X9981 a_21478_18894# nmat.rowon_n[5] a_21082_18934# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9982 a_45574_14878# nmat.col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9983 a_7730_69109# a_2149_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X9984 a_34530_59182# pmat.col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9985 a_2557_74031# a_1923_69823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9986 a_36634_72556# pmat.col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9987 a_28506_24918# nmat.col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9988 VDD a_13432_62581# a_3923_68021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9989 vcm a_18162_9492# a_27198_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X999 a_20474_64202# pmat.col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9990 VDD pmat.rowon_n[14] a_40158_70186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9991 vcm a_18162_69222# a_22178_69182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9992 a_32126_16926# pmat.row_n[8] a_32618_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9993 VSS config_1_in[11] a_1626_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9994 VDD pmat.rowon_n[4] a_36142_60146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9995 a_11611_50332# a_11416_50363# a_11921_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X9996 a_34002_44527# a_33825_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9997 a_36142_62154# a_18162_62194# a_36234_62154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9998 VSS config_2_in[10] a_1591_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9999 a_49686_71552# pmat.col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
C0 _1192_.A2 _1183_.A2 4.98fF
C1 _1184_.A2 a_26891_28327# 2.00fF
C2 VDD a_1674_68047# 5.58fF
C3 m2_17932_71010# m3_18064_71142# 2.76fF
C4 a_12449_22895# nmat.col_n[1] 0.76fF
C5 VDD a_1923_53055# 2.81fF
C6 pmat.col_n[4] ctopp 2.02fF
C7 a_11071_36694# a_10873_36341# 0.30fF
C8 VDD a_37739_36649# 0.61fF
C9 a_35230_70186# vcm 0.62fF
C10 VDD a_30118_72194# 0.32fF
C11 a_22178_11500# vcm 0.65fF
C12 a_11067_64015# pmat.rowon_n[1] 0.68fF
C13 a_2835_13077# a_2411_16101# 2.09fF
C14 a_38851_28327# a_29937_31055# 0.39fF
C15 a_1586_18231# a_1591_27797# 0.33fF
C16 a_11339_39319# a_19505_38779# 0.33fF
C17 a_30663_50087# a_45450_48695# 0.66fF
C18 VDD a_18546_24550# 36.82fF
C19 ANTENNA__1184__B1.DIODE a_25879_31591# 0.94fF
C20 VDD config_2_in[14] 1.10fF
C21 nmat.sw m2_50060_24282# 0.32fF
C22 a_24186_19532# ctopn 3.58fF
C23 VDD a_38299_29673# 0.39fF
C24 VDD a_24186_21540# 0.52fF
C25 a_18546_59184# a_48190_59142# 0.35fF
C26 a_37238_65166# a_37238_64162# 1.00fF
C27 a_8695_63937# a_8656_63811# 0.72fF
C28 a_23182_10496# ctopn 3.58fF
C29 a_44266_57134# ctopp 3.57fF
C30 a_43262_71190# ctopp 3.40fF
C31 a_24833_34191# a_26767_34967# 0.59fF
C32 a_1899_35051# a_6283_31591# 0.43fF
C33 VDD a_2411_43301# 11.80fF
C34 a_30210_58138# ctopp 3.58fF
C35 a_26194_68178# vcm 0.62fF
C36 VDD a_1923_61759# 13.11fF
C37 VDD result_out[7] 0.65fF
C38 VDD a_39246_58138# 0.52fF
C39 a_2879_57487# a_5779_71285# 3.09fF
C40 a_46274_23548# a_47278_23548# 0.97fF
C41 a_16311_28327# a_35244_32411# 0.68fF
C42 a_2021_26677# cgen.start_conv_in 1.83fF
C43 a_26194_16520# a_26194_15516# 1.00fF
C44 pmat.row_n[2] ctopn 1.65fF
C45 a_48282_9492# a_49286_9492# 0.97fF
C46 a_18546_60188# a_24094_60146# 0.35fF
C47 cgen.dlycontrol4_in[1] a_3183_19258# 0.59fF
C48 a_6835_51183# a_4259_31375# 0.91fF
C49 m2_51064_18258# vcm 0.51fF
C50 a_15667_27239# a_38851_28327# 1.68fF
C51 a_11892_21959# a_7693_22365# 0.44fF
C52 pmat.rowoff_n[12] cgen.dlycontrol3_in[2] 0.67fF
C53 a_22628_30485# a_15101_29423# 0.86fF
C54 VDD a_44444_32233# 3.63fF
C55 a_1769_13103# config_1_in[14] 0.33fF
C56 a_4719_30287# a_2411_43301# 0.77fF
C57 a_17139_30503# nmat.col[13] 1.05fF
C58 a_31214_23548# vcm 0.65fF
C59 a_22178_69182# ctopp 3.58fF
C60 a_18546_19530# a_19074_19938# 0.35fF
C61 ANTENNA__1190__A1.DIODE nmat.col_n[23] 0.33fF
C62 a_33222_9492# vcm 0.65fF
C63 VDD a_31214_69182# 0.52fF
C64 a_18546_22542# a_50198_22950# 0.35fF
C65 nmat.col_n[4] ctopn 2.02fF
C66 a_49286_20536# vcm 0.65fF
C67 a_29159_39783# a_29159_37607# 0.77fF
C68 a_1769_47919# a_1823_58237# 0.44fF
C69 a_38242_65166# a_39246_65166# 0.97fF
C70 a_31214_59142# ctopp 3.58fF
C71 VDD nmat.col[23] 4.58fF
C72 m2_17932_67998# m3_18064_68130# 2.76fF
C73 a_25190_11500# ctopn 3.58fF
C74 a_1769_13103# config_2_in[6] 0.35fF
C75 VDD a_42307_31756# 0.39fF
C76 VDD a_40250_59142# 0.52fF
C77 _1184_.A2 a_9411_2215# 6.30fF
C78 a_45270_21540# a_46274_21540# 0.97fF
C79 VDD a_4265_71543# 1.07fF
C80 nmat.col_n[13] ctopn 2.02fF
C81 pmat.row_n[5] ctopp 1.65fF
C82 a_22199_30287# nmat.col[28] 0.76fF
C83 VDD m2_17932_13238# 1.00fF
C84 ANTENNA_fanout52_A.DIODE a_25879_31591# 0.49fF
C85 a_30641_44743# a_11149_40188# 0.38fF
C86 a_13459_28111# a_30663_50087# 3.07fF
C87 a_18546_16518# a_36142_16926# 0.35fF
C88 nmat.rowoff_n[6] ctopn 0.60fF
C89 m2_18936_24282# vcm 0.41fF
C90 a_12447_16143# a_10883_3303# 4.01fF
C91 m2_17932_23278# m2_18936_23278# 0.96fF
C92 a_18546_70228# a_18162_70226# 2.62fF
C93 a_46274_71190# a_46274_70186# 1.00fF
C94 VDD pmat.rowoff_n[13] 2.19fF
C95 a_3866_57399# a_5731_58951# 0.85fF
C96 VDD pmat.rowoff_n[9] 2.47fF
C97 a_13503_37981# a_12513_36924# 0.39fF
C98 a_10055_31591# a_10515_13967# 0.81fF
C99 a_19541_28879# a_10441_21263# 0.48fF
C100 a_29206_13508# vcm 0.65fF
C101 _1187_.A2 a_40837_46261# 0.86fF
C102 ANTENNA__1395__A1.DIODE _1192_.A2 1.76fF
C103 a_18546_62196# vcm 0.40fF
C104 m2_45040_7214# m2_46044_7214# 0.96fF
C105 a_29163_38545# a_23821_35279# 0.32fF
C106 a_17139_30503# nmat.col_n[27] 0.77fF
C107 a_27198_18528# vcm 0.65fF
C108 VDD a_1757_20181# 0.63fF
C109 a_7717_14735# clk_ena 0.56fF
C110 a_4075_50087# a_6559_57167# 0.34fF
C111 _1184_.A2 a_7939_31591# 0.30fF
C112 a_44266_13508# a_45270_13508# 0.97fF
C113 nmat.sw cgen.dlycontrol3_in[2] 1.63fF
C114 VDD m3_31116_72146# 0.40fF
C115 a_18162_21540# ctopn 1.49fF
C116 a_24591_28327# nmat.col[19] 1.11fF
C117 a_38242_15516# vcm 0.65fF
C118 VDD a_23182_17524# 0.52fF
C119 VDD a_32687_46607# 6.88fF
C120 a_18563_27791# a_12987_26159# 0.49fF
C121 a_42258_18528# a_43262_18528# 0.97fF
C122 VDD a_24186_8488# 0.55fF
C123 a_18546_21538# a_27106_21946# 0.35fF
C124 a_11067_64015# ANTENNA__1395__A1.DIODE 1.10fF
C125 a_29206_62154# a_29206_61150# 1.00fF
C126 ANTENNA__1184__B1.DIODE ndecision_finish 2.30fF
C127 a_34226_23548# ctopn 3.46fF
C128 a_2659_35015# a_4257_34319# 0.73fF
C129 VDD a_40250_19532# 0.52fF
C130 a_36234_9492# ctopn 3.57fF
C131 a_11927_27399# nmat.col[13] 0.41fF
C132 nmat.col_n[21] nmat.col[21] 0.87fF
C133 VDD a_9545_66567# 2.39fF
C134 a_34226_60146# vcm 0.62fF
C135 VDD a_39246_10496# 0.52fF
C136 VDD a_6311_42692# 0.67fF
C137 a_27913_42333# a_27947_41245# 0.46fF
C138 a_29206_15516# a_29206_14512# 1.00fF
C139 VDD a_2944_65576# 0.55fF
C140 a_2835_13077# a_9675_10396# 0.36fF
C141 m2_17932_64986# m3_18064_65118# 2.76fF
C142 a_18546_58180# a_46182_58138# 0.35fF
C143 a_31214_69182# a_31214_68178# 1.00fF
C144 nmat.rowon_n[7] a_3688_17179# 0.60fF
C145 pmat.row_n[4] a_2315_44124# 1.46fF
C146 a_18546_10494# a_46182_10902# 0.35fF
C147 a_39246_21540# a_39246_20536# 1.00fF
C148 VDD a_20711_34191# 0.35fF
C149 a_10239_14183# a_6927_30503# 0.42fF
C150 pmat.row_n[5] a_3746_58487# 2.00fF
C151 VDD a_18162_12504# 2.74fF
C152 a_46274_62154# ctopp 3.58fF
C153 a_40250_16520# vcm 0.65fF
C154 a_13779_43123# a_10949_43124# 0.75fF
C155 a_3339_70759# a_7563_63303# 0.77fF
C156 cgen.dlycontrol4_in[4] a_1586_18231# 0.86fF
C157 a_32218_13508# ctopn 3.58fF
C158 a_27198_57134# vcm 0.62fF
C159 a_26194_71190# vcm 0.60fF
C160 a_30210_18528# ctopn 3.58fF
C161 VDD a_10927_41245# 0.71fF
C162 a_8583_29199# a_15667_28111# 1.46fF
C163 pmat.row_n[15] a_10515_15055# 1.46fF
C164 nmat.col_n[30] nmat.col[28] 2.12fF
C165 inn_analog nmat.col[21] 0.38fF
C166 a_10873_38517# a_10927_37981# 0.30fF
C167 a_45270_70186# ctopp 3.57fF
C168 nmat.sw nmat.col[25] 0.61fF
C169 VDD a_77428_40594# 0.31fF
C170 VDD a_12907_54997# 0.51fF
C171 VDD a_7674_69135# 1.32fF
C172 a_41254_15516# ctopn 3.58fF
C173 VDD a_41254_11500# 0.52fF
C174 a_4383_7093# a_6448_5755# 0.46fF
C175 a_12513_39100# a_13597_37571# 0.38fF
C176 ANTENNA__1395__A2.DIODE _1192_.A2 3.59fF
C177 a_3339_70759# a_4396_69109# 0.58fF
C178 pmat.rowoff_n[8] pmat.row_n[8] 0.71fF
C179 a_50290_23548# a_50290_22544# 1.00fF
C180 a_6467_29415# a_1923_31743# 0.49fF
C181 VDD m2_31988_54946# 0.62fF
C182 a_40837_46261# a_46753_41935# 0.38fF
C183 a_49286_60146# a_50290_60146# 0.97fF
C184 nmat.rowon_n[13] nmat.rowon_n[6] 0.69fF
C185 a_2046_30184# a_2787_33237# 0.42fF
C186 a_18546_69224# a_41162_69182# 0.35fF
C187 VDD a_37471_32149# 0.30fF
C188 a_1923_61759# a_1823_60949# 0.70fF
C189 a_33222_11500# a_33222_10496# 1.00fF
C190 VDD a_19166_13508# 0.56fF
C191 a_10513_24135# a_8197_20871# 0.48fF
C192 a_24867_53135# a_11067_27239# 0.33fF
C193 ANTENNA__1184__B1.DIODE a_24591_28327# 1.59fF
C194 a_13091_52047# a_18823_50247# 0.35fF
C195 cgen.dlycontrol4_in[5] a_12197_43746# 5.25fF
C196 a_37820_30485# a_45187_38129# 0.30fF
C197 a_18546_8486# ctopn 1.30fF
C198 pmat.en_bit_n[2] ANTENNA__1197__A.DIODE 1.67fF
C199 a_1957_43567# a_1586_50247# 0.40fF
C200 cgen.dlycontrol3_in[2] a_12116_40871# 0.31fF
C201 a_12061_26703# nmat.col[3] 3.16fF
C202 a_38242_22544# vcm 0.65fF
C203 a_38242_61150# a_39246_61150# 0.97fF
C204 pmat.rowon_n[5] pmat.row_n[3] 0.46fF
C205 a_36234_68178# ctopp 3.58fF
C206 nmat.col_n[13] a_10498_19631# 0.33fF
C207 VDD a_45270_68178# 0.52fF
C208 pmat.col[27] m2_46044_54946# 0.39fF
C209 a_23182_12504# a_23182_11500# 1.00fF
C210 a_19166_22544# a_19166_21540# 1.00fF
C211 a_18162_65206# ctopp 1.49fF
C212 VDD a_21087_43177# 0.63fF
C213 a_4351_55527# a_5363_70543# 0.72fF
C214 pmat.row_n[6] a_18546_14510# 0.35fF
C215 ANTENNA__1190__A1.DIODE _1187_.A2 0.44fF
C216 pmat.sample_n a_32687_46607# 0.52fF
C217 m2_17932_61974# m3_18064_62106# 2.76fF
C218 a_7415_29397# a_7026_24527# 1.40fF
C219 VDD a_22216_30761# 0.70fF
C220 pmat.row_n[13] ctopp 1.65fF
C221 VDD pmat.rowoff_n[0] 1.88fF
C222 a_32218_20536# a_33222_20536# 0.97fF
C223 a_18546_20534# a_47186_20942# 0.35fF
C224 a_43262_16520# ctopn 3.58fF
C225 VDD a_4719_69929# 0.32fF
C226 VDD m2_23956_7214# 1.08fF
C227 a_20170_15516# vcm 0.65fF
C228 _1194_.B1 a_23933_32143# 0.55fF
C229 VDD a_6607_75895# 0.39fF
C230 a_18546_62196# a_32126_62154# 0.35fF
C231 nmat.col[30] vcm 8.25fF
C232 a_45270_67174# a_45270_66170# 1.00fF
C233 a_18546_66212# a_28110_66170# 0.35fF
C234 a_31214_9492# a_31214_8488# 1.00fF
C235 VDD a_50290_23548# 0.59fF
C236 VDD a_21174_66170# 0.52fF
C237 a_18546_11498# a_50198_11906# 0.35fF
C238 a_2199_13887# a_7939_7125# 0.33fF
C239 pmat.row_n[9] nmat.sample 0.34fF
C240 a_3339_70759# a_7467_63303# 0.63fF
C241 a_44266_17524# a_45270_17524# 0.97fF
C242 pmat.sw a_7717_14735# 0.89fF
C243 a_3923_68021# a_12993_66415# 0.45fF
C244 a_14641_57711# pmat.row_n[10] 0.30fF
C245 a_42258_57134# a_43262_57134# 0.97fF
C246 _1192_.A2 ANTENNA__1196__A2.DIODE 6.82fF
C247 ANTENNA__1195__A1.DIODE a_12263_50959# 0.50fF
C248 a_47278_20536# a_47278_19532# 1.00fF
C249 a_41254_71190# a_42258_71190# 0.97fF
C250 a_28202_58138# a_29206_58138# 0.97fF
C251 VDD a_14261_44219# 1.32fF
C252 a_46274_14512# vcm 0.65fF
C253 pmat.rowon_n[8] a_12263_50959# 0.34fF
C254 a_45270_64162# vcm 0.62fF
C255 a_27498_32117# a_27443_32143# 0.51fF
C256 VDD a_36539_47113# 0.36fF
C257 a_45270_8488# a_46274_8488# 0.97fF
C258 a_19166_65166# a_19166_64162# 1.00fF
C259 VDD a_20170_55126# 0.60fF
C260 VDD a_42701_31849# 0.51fF
C261 a_3339_59879# a_6175_60039# 0.42fF
C262 a_11921_37462# nmat.sample 0.44fF
C263 _1179_.X ANTENNA__1184__B1.DIODE 2.15fF
C264 a_21279_48999# a_28901_48437# 0.33fF
C265 a_33467_46261# a_33423_47695# 2.01fF
C266 VDD a_48282_13508# 0.52fF
C267 pmat.en_bit_n[0] _1192_.B1 1.91fF
C268 a_41254_22544# ctopn 3.57fF
C269 VDD a_46274_18528# 0.52fF
C270 a_20170_71190# m2_19940_72014# 1.00fF
C271 a_11067_64015# ANTENNA__1196__A2.DIODE 1.51fF
C272 a_28202_61150# a_28202_60146# 1.00fF
C273 pmat.row_n[11] ctopp 1.65fF
C274 a_18162_61190# ctopp 1.49fF
C275 a_36234_19532# a_36234_18528# 1.00fF
C276 a_18546_70228# a_30118_70186# 0.35fF
C277 nmat.col[9] nmat.col_n[8] 6.70fF
C278 a_1586_50247# cgen.enable_dlycontrol_in 0.97fF
C279 VDD a_38737_41814# 1.45fF
C280 a_18546_14510# a_48190_14918# 0.35fF
C281 a_29206_62154# vcm 0.62fF
C282 VDD a_1591_63701# 0.45fF
C283 a_18546_17522# a_25098_17930# 0.35fF
C284 pmat.rowon_n[7] pmat.row_n[5] 2.04fF
C285 a_18546_64204# a_46182_64162# 0.35fF
C286 m2_17932_58962# m3_18064_59094# 2.76fF
C287 a_11067_27239# a_38851_28327# 0.47fF
C288 _1192_.B1 a_32405_32463# 0.99fF
C289 a_19166_62154# pmat.col[0] 0.31fF
C290 a_18546_57176# a_21082_57134# 0.35fF
C291 pmat.rowoff_n[12] a_2263_43719# 1.89fF
C292 a_29206_59142# a_29206_58138# 1.00fF
C293 a_1923_69823# a_1823_76181# 0.54fF
C294 a_19541_28879# a_12604_47080# 0.43fF
C295 a_3746_58487# cgen.enable_dlycontrol_in 0.69fF
C296 VDD a_12815_26409# 0.45fF
C297 a_4075_50087# a_5784_52423# 1.59fF
C298 a_21174_15516# a_22178_15516# 0.97fF
C299 a_18546_15514# a_25098_15922# 0.35fF
C300 a_48282_65166# vcm 0.62fF
C301 VDD a_17927_47349# 0.34fF
C302 a_44266_60146# ctopp 3.58fF
C303 a_20170_69182# a_21174_69182# 0.97fF
C304 VDD a_3175_59585# 0.47fF
C305 a_28202_70186# vcm 0.62fF
C306 nmat.col[15] a_34226_24552# 0.40fF
C307 a_34226_17524# a_34226_16520# 1.00fF
C308 a_20170_22544# vcm 0.65fF
C309 VDD a_11897_21263# 0.73fF
C310 a_18546_68220# ctopp 1.59fF
C311 a_49286_14512# ctopn 3.57fF
C312 a_40250_12504# a_41254_12504# 0.97fF
C313 pmat.rowoff_n[15] a_9457_51163# 0.32fF
C314 a_4409_74183# a_5363_73807# 0.40fF
C315 ANTENNA_fanout52_A.DIODE _1179_.X 0.36fF
C316 a_29206_59142# a_30210_59142# 0.97fF
C317 a_18546_59184# a_41162_59142# 0.35fF
C318 a_13432_62581# a_13091_52047# 0.76fF
C319 a_37238_57134# ctopp 3.57fF
C320 VDD a_46339_31029# 0.98fF
C321 ANTENNA_fanout52_A.DIODE a_33423_47695# 0.32fF
C322 a_36234_71190# ctopp 3.40fF
C323 VDD a_46274_57134# 0.52fF
C324 _1154_.X nmat.col[30] 0.34fF
C325 a_23182_58138# ctopp 3.58fF
C326 VDD a_45270_71190# 0.55fF
C327 VDD a_32218_58138# 0.52fF
C328 pmat.row_n[11] a_5351_19913# 0.45fF
C329 VDD a_13183_72405# 0.47fF
C330 a_29206_62154# pmat.col[10] 0.31fF
C331 a_39246_71190# m2_39016_72014# 1.00fF
C332 pmat.col_n[11] pmat.col[11] 0.74fF
C333 VDD a_17927_48437# 0.36fF
C334 a_22153_37179# a_22537_36911# 0.33fF
C335 _1196_.B1 a_24867_53135# 0.68fF
C336 a_2163_53057# a_2124_52931# 0.75fF
C337 pmat.row_n[7] a_12263_50959# 0.58fF
C338 ANTENNA__1183__B1.DIODE nmat.col_n[30] 2.73fF
C339 pmat.rowon_n[7] a_1957_43567# 0.52fF
C340 a_10515_15055# pmat.rowon_n[3] 0.68fF
C341 VDD a_31793_41570# 3.84fF
C342 a_13459_28111# a_10883_3303# 1.08fF
C343 pmat.row_n[0] a_12079_9615# 1.83fF
C344 m2_26968_7214# m3_27100_7346# 2.79fF
C345 a_35230_55126# a_36234_55126# 0.97fF
C346 a_18546_24550# a_46182_24958# 0.35fF
C347 VDD a_12345_39100# 3.50fF
C348 m2_17932_55950# m3_18064_56082# 2.76fF
C349 a_25190_68178# a_25190_67174# 1.00fF
C350 a_9963_13967# a_14653_53458# 0.32fF
C351 a_24186_23548# vcm 0.65fF
C352 a_26194_9492# vcm 0.65fF
C353 VDD a_24186_69182# 0.52fF
C354 a_48282_61150# vcm 0.62fF
C355 VDD a_4627_50095# 0.48fF
C356 a_18546_22542# a_43170_22950# 0.35fF
C357 pmat.col_n[29] pmat.col[28] 0.39fF
C358 _1154_.X a_25695_28111# 0.87fF
C359 VDD m2_21948_24282# 0.62fF
C360 _1192_.B1 pmat.col[8] 0.35fF
C361 a_42258_20536# vcm 0.65fF
C362 a_11041_39860# a_22269_40391# 0.34fF
C363 a_24186_59142# ctopp 3.58fF
C364 VDD a_33222_59142# 0.52fF
C365 _1154_.X a_1781_9308# 0.35fF
C366 VDD a_2467_35015# 0.38fF
C367 cgen.dlycontrol4_in[3] a_11041_39860# 0.64fF
C368 a_13091_28327# a_25879_31591# 4.54fF
C369 a_23182_16520# a_24186_16520# 0.97fF
C370 a_18546_16518# a_29114_16926# 0.35fF
C371 _1192_.A2 a_12053_27497# 0.37fF
C372 VDD a_7803_67655# 0.44fF
C373 _1519_.A ctopp 2.16fF
C374 VDD a_8193_61493# 1.26fF
C375 a_4127_37013# a_4031_37191# 0.39fF
C376 a_22178_13508# vcm 0.65fF
C377 m2_38012_7214# m2_39016_7214# 0.96fF
C378 a_10767_39087# a_14589_40726# 0.46fF
C379 a_1923_69823# a_3175_72641# 0.32fF
C380 pmat.col_n[15] pmat.col[15] 0.94fF
C381 a_1899_35051# a_4128_46983# 0.31fF
C382 a_8305_20871# a_4383_7093# 0.57fF
C383 m2_51064_59966# m2_51064_58962# 0.99fF
C384 VDD pmat.rowon_n[14] 3.61fF
C385 pmat.row_n[8] ctopn 1.65fF
C386 a_31214_15516# vcm 0.65fF
C387 a_43720_32143# a_32405_32463# 1.71fF
C388 VDD a_11823_74895# 0.41fF
C389 VDD a_14528_48114# 0.30fF
C390 a_31214_63158# pmat.col[12] 0.31fF
C391 m2_18936_72014# m3_19068_72146# 2.79fF
C392 _1154_.A a_30571_50959# 0.60fF
C393 a_32218_70186# a_32218_69182# 1.00fF
C394 VDD a_6651_33239# 0.31fF
C395 a_25879_31591# a_27155_31599# 0.94fF
C396 VDD a_4003_7663# 0.36fF
C397 pmat.rowoff_n[15] ctopn 1.17fF
C398 a_50290_12504# vcm 0.65fF
C399 nmat.col_n[0] m2_18936_24282# 0.37fF
C400 ANTENNA__1197__A.DIODE nmat.col_n[18] 0.60fF
C401 a_21174_14512# a_21174_13508# 1.00fF
C402 nmat.col[5] ctopn 1.97fF
C403 nmat.col[16] vcm 5.76fF
C404 a_4167_30511# a_4333_30511# 0.69fF
C405 a_27198_23548# ctopn 3.40fF
C406 VDD a_33222_19532# 0.52fF
C407 cgen.enable_dlycontrol_in cgen.start_conv_in 1.14fF
C408 m2_44036_54946# m3_44168_55078# 2.79fF
C409 a_29206_9492# ctopn 3.57fF
C410 VDD m2_41024_72014# 0.98fF
C411 a_25190_57134# a_25190_56130# 1.00fF
C412 a_29206_19532# a_30210_19532# 0.97fF
C413 pmat.col_n[31] pmat.col[31] 1.14fF
C414 VDD a_1823_68565# 3.81fF
C415 a_27198_60146# vcm 0.62fF
C416 nmat.col_n[13] nmat.col[14] 6.69fF
C417 VDD a_32218_10496# 0.52fF
C418 a_3746_58487# a_2659_35015# 1.70fF
C419 pmat.rowon_n[3] cgen.dlycontrol4_in[3] 0.53fF
C420 a_3339_70759# a_5363_70543# 0.36fF
C421 VDD a_32072_38567# 1.34fF
C422 a_19541_28879# a_5535_29980# 2.38fF
C423 a_45270_20536# ctopn 3.58fF
C424 pmat.row_n[2] ctopp 1.67fF
C425 a_10883_3303# a_9528_20407# 0.49fF
C426 a_4843_54826# pmat.rowon_n[0] 0.77fF
C427 a_19166_57134# ctopp 3.24fF
C428 a_18546_58180# a_39154_58138# 0.35fF
C429 a_24591_28327# nmat.col_n[29] 0.31fF
C430 a_28202_10496# a_29206_10496# 0.97fF
C431 a_18546_10494# a_39154_10902# 0.35fF
C432 VDD a_1757_33775# 0.61fF
C433 a_28901_48437# a_29076_48695# 1.72fF
C434 a_11067_30287# a_14887_46377# 2.49fF
C435 a_39246_62154# ctopp 3.58fF
C436 VDD a_48282_62154# 0.52fF
C437 a_33222_16520# vcm 0.65fF
C438 a_11317_40188# cgen.dlycontrol4_in[1] 0.45fF
C439 a_17139_30503# a_25879_31591# 2.60fF
C440 a_3367_14906# a_3229_14741# 0.42fF
C441 a_39246_56130# a_40250_56130# 0.97fF
C442 VDD a_12247_20175# 0.55fF
C443 VDD a_12693_38543# 0.82fF
C444 VDD ANTENNA__1197__B.DIODE 19.70fF
C445 nmat.col[1] comp_latch 2.94fF
C446 a_25190_13508# ctopn 3.58fF
C447 VDD a_10378_7637# 0.97fF
C448 cgen.dlycontrol4_in[3] a_2648_29397# 0.40fF
C449 a_20170_57134# vcm 0.62fF
C450 VDD a_18180_38341# 1.36fF
C451 pmat.sw ANTENNA__1195__A1.DIODE 0.98fF
C452 a_23182_18528# ctopn 3.58fF
C453 a_19166_10496# m2_17932_10226# 0.96fF
C454 VDD a_27877_42043# 1.18fF
C455 VDD a_18546_14510# 32.63fF
C456 VDD pmat.row_n[6] 29.35fF
C457 a_28704_29568# a_37291_29397# 1.10fF
C458 nmat.col_n[28] nmat.col[26] 0.70fF
C459 ANTENNA__1196__A2.DIODE a_3571_13627# 1.29fF
C460 pmat.rowon_n[8] pmat.sw 2.66fF
C461 pmat.row_n[13] nmat.rowoff_n[1] 0.78fF
C462 cgen.enable_dlycontrol_in cgen.dlycontrol3_in[1] 1.62fF
C463 a_38242_70186# ctopp 3.57fF
C464 a_34226_15516# ctopn 3.58fF
C465 VDD a_47278_70186# 0.52fF
C466 VDD a_34226_11500# 0.52fF
C467 a_18546_72236# a_47186_72194# 0.35fF
C468 pmat.row_n[11] pmat.rowon_n[7] 0.39fF
C469 a_6787_47607# a_3746_58487# 0.40fF
C470 pmat.row_n[10] pmat.row_n[8] 14.75fF
C471 pmat.rowoff_n[12] a_10055_31591# 0.59fF
C472 a_21174_22544# a_22178_22544# 0.97fF
C473 pmat.col_n[21] ANTENNA__1195__A1.DIODE 0.38fF
C474 VDD a_43267_28879# 0.63fF
C475 a_44266_62154# a_45270_62154# 0.97fF
C476 VDD a_31675_47695# 9.66fF
C477 a_42258_66170# a_43262_66170# 0.97fF
C478 a_21739_29415# a_22199_30287# 7.94fF
C479 a_18546_69224# a_34134_69182# 0.35fF
C480 VDD a_24374_29941# 2.35fF
C481 VDD a_7299_58951# 0.35fF
C482 pmat.col_n[7] ctopp 2.02fF
C483 a_11041_36596# a_12069_36341# 1.42fF
C484 a_49286_56130# vcm 0.62fF
C485 VDD a_33130_72194# 0.32fF
C486 a_35230_63158# a_36234_63158# 0.97fF
C487 pmat.rowoff_n[12] a_1591_31599# 4.29fF
C488 a_31214_22544# vcm 0.65fF
C489 nmat.col_n[18] m2_37008_24282# 0.38fF
C490 a_29206_68178# ctopp 3.58fF
C491 VDD a_38242_68178# 0.52fF
C492 nmat.col_n[31] nmat.col_n[26] 0.82fF
C493 a_19166_12504# a_19166_11500# 1.00fF
C494 _1224_.X vcm 1.17fF
C495 a_30663_50087# a_32405_32463# 0.42fF
C496 a_45270_63158# vcm 0.62fF
C497 a_2407_49289# a_2879_57487# 0.44fF
C498 inp_analog ctopp 0.93fF
C499 a_44763_34293# nmat.col_n[26] 1.02fF
C500 a_18546_20534# a_40158_20942# 0.35fF
C501 a_11508_48187# a_11547_48061# 0.79fF
C502 a_36234_16520# ctopn 3.58fF
C503 ANTENNA_fanout52_A.DIODE nmat.sample_n 0.57fF
C504 a_4339_27804# a_9441_20189# 0.34fF
C505 VDD a_82787_54421# 0.59fF
C506 a_12237_38772# a_12228_40693# 0.35fF
C507 VDD a_9287_77055# 0.37fF
C508 a_18546_62196# a_25098_62154# 0.35fF
C509 a_18546_66212# a_21082_66170# 0.35fF
C510 a_22153_37179# a_12309_36483# 0.73fF
C511 _1154_.X nmat.col[16] 0.31fF
C512 nmat.rowon_n[2] vcm 0.56fF
C513 _1224_.X _1194_.B1 1.88fF
C514 VDD a_43262_23548# 0.55fF
C515 a_43262_70186# a_44266_70186# 0.97fF
C516 VDD a_45270_9492# 0.52fF
C517 a_2411_33749# a_9983_32385# 0.33fF
C518 a_30210_11500# a_31214_11500# 0.97fF
C519 a_18546_11498# a_43170_11906# 0.35fF
C520 a_10055_31591# nmat.sw 2.12fF
C521 a_10515_61839# pmat.rowon_n[3] 0.44fF
C522 a_40250_56130# m2_40020_54946# 0.99fF
C523 a_26891_28327# a_25879_31591# 0.75fF
C524 a_18563_27791# a_31263_28309# 1.09fF
C525 a_32218_64162# a_32218_63158# 1.00fF
C526 m2_51064_61974# vcm 0.50fF
C527 m2_18936_54946# m3_19068_55078# 2.79fF
C528 a_9307_31068# clk_ena 1.07fF
C529 a_35230_10496# a_35230_9492# 1.00fF
C530 a_20170_19532# a_21174_19532# 0.97fF
C531 a_50290_67174# vcm 0.62fF
C532 a_32218_58138# a_32218_57134# 1.00fF
C533 VDD a_3609_9295# 0.40fF
C534 a_39246_14512# vcm 0.65fF
C535 cgen.start_conv_in a_2411_33749# 0.47fF
C536 a_25997_42902# a_10873_40693# 0.31fF
C537 a_5363_33551# a_14379_6567# 1.52fF
C538 nmat.rowon_n[1] nmat.rowoff_n[1] 23.21fF
C539 a_38242_64162# vcm 0.62fF
C540 VDD m2_45040_24282# 0.62fF
C541 VDD a_35540_46983# 0.38fF
C542 nmat.col[18] ctopn 2.28fF
C543 a_36234_60146# a_36234_59142# 1.00fF
C544 a_1923_53055# a_2163_58941# 0.34fF
C545 a_41731_49525# nmat.col[28] 0.90fF
C546 a_24186_18528# a_24186_17524# 1.00fF
C547 VDD a_7663_27247# 0.31fF
C548 VDD vcm.sky130_fd_sc_hd__buf_4_0.A 0.44fF
C549 a_10515_15055# a_4068_25615# 0.49fF
C550 nmat.rowon_n[7] a_4516_21531# 1.01fF
C551 VDD a_14691_27399# 1.75fF
C552 a_11921_37462# cgen.dlycontrol1_in[3] 0.34fF
C553 a_18546_10494# a_21082_10902# 0.35fF
C554 nmat.en_bit_n[1] a_18243_28327# 0.67fF
C555 a_24591_28327# a_13091_28327# 0.91fF
C556 a_5991_23983# a_4703_24527# 1.00fF
C557 VDD a_41254_13508# 0.52fF
C558 a_4351_55527# a_4081_61127# 0.39fF
C559 a_34226_22544# ctopn 3.58fF
C560 a_14287_69455# pmat.col[0] 0.69fF
C561 a_2659_35015# cgen.start_conv_in 0.77fF
C562 a_35290_44527# a_11149_40188# 0.44fF
C563 a_13779_43123# cgen.dlycontrol4_in[2] 0.96fF
C564 VDD a_39246_18528# 0.52fF
C565 a_24186_63158# a_24186_62154# 1.00fF
C566 m2_26968_24282# vcm 0.42fF
C567 a_40250_67174# a_41254_67174# 0.97fF
C568 nmat.col[31] nmat.col_n[30] 7.24fF
C569 nmat.col_n[15] vcm 2.79fF
C570 a_24407_31375# nmat.col_n[31] 0.53fF
C571 a_18546_70228# a_23090_70186# 0.35fF
C572 a_15667_27239# a_20439_27247# 2.36fF
C573 a_6451_67655# a_4583_68021# 1.11fF
C574 pmat.col_n[4] pmat.col[4] 0.75fF
C575 a_37238_66170# a_37238_65166# 1.00fF
C576 a_30210_22544# a_30210_21540# 1.00fF
C577 VDD a_20811_42359# 0.59fF
C578 ANTENNA__1190__B1.DIODE _1192_.A2 6.85fF
C579 VDD a_50290_15516# 0.54fF
C580 a_18546_14510# a_41162_14918# 0.35fF
C581 a_29206_14512# a_30210_14512# 0.97fF
C582 a_22178_62154# vcm 0.62fF
C583 a_18546_24550# a_19074_24958# 0.35fF
C584 VDD a_9227_20291# 0.31fF
C585 a_28202_64162# a_29206_64162# 0.97fF
C586 a_18546_64204# a_39154_64162# 0.35fF
C587 a_34226_68178# a_35230_68178# 0.97fF
C588 VDD a_28812_29575# 1.96fF
C589 pmat.col_n[23] pmat.col[23] 0.83fF
C590 a_29206_8488# m2_28976_7214# 1.00fF
C591 a_23182_13508# a_23182_12504# 1.00fF
C592 a_41254_65166# vcm 0.62fF
C593 VDD a_6082_46831# 0.78fF
C594 a_48282_21540# vcm 0.65fF
C595 a_18546_8486# a_18162_8488# 2.61fF
C596 a_37238_60146# ctopp 3.58fF
C597 vcm comp_latch 1.24fF
C598 VDD a_46274_60146# 0.52fF
C599 a_21174_70186# vcm 0.62fF
C600 VDD a_12003_52815# 0.58fF
C601 a_10055_31591# a_1858_25615# 0.94fF
C602 pmat.row_n[15] pmat.rowoff_n[10] 1.32fF
C603 a_7415_29397# a_27001_30511# 0.52fF
C604 a_18546_17522# vcm 0.40fF
C605 _1154_.X _1224_.X 1.13fF
C606 a_25879_31591# a_9411_2215# 0.73fF
C607 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col[18] 0.41fF
C608 a_13641_23439# nmat.col[7] 0.75fF
C609 a_19166_8488# vcm 0.63fF
C610 a_42258_14512# ctopn 3.58fF
C611 pmat.col_n[21] pmat.col[21] 0.74fF
C612 VDD a_13443_43447# 0.61fF
C613 VDD a_11603_28335# 0.95fF
C614 _1179_.X a_13091_28327# 1.33fF
C615 a_18546_59184# a_34134_59142# 0.35fF
C616 a_30210_65166# a_30210_64162# 1.00fF
C617 pmat.row_n[15] a_4951_31029# 0.40fF
C618 a_30210_57134# ctopp 3.57fF
C619 a_10991_68591# a_11837_68591# 0.71fF
C620 VDD a_22459_28879# 1.67fF
C621 a_29206_71190# ctopp 3.40fF
C622 VDD a_39246_57134# 0.52fF
C623 a_1957_43567# a_4259_31375# 0.49fF
C624 VDD a_32162_34191# 0.40fF
C625 VDD a_38242_71190# 0.55fF
C626 VDD a_25190_58138# 0.52fF
C627 a_39246_23548# a_40250_23548# 0.97fF
C628 VDD vcm.sky130_fd_sc_hd__nand2_1_1.Y 0.48fF
C629 m2_51064_16250# m2_51064_15246# 0.99fF
C630 a_41254_9492# a_42258_9492# 0.97fF
C631 VDD a_46135_38127# 1.03fF
C632 a_48282_12504# a_48282_11500# 1.00fF
C633 pmat.row_n[7] a_12447_16143# 0.32fF
C634 pmat.rowon_n[7] pmat.row_n[2] 0.71fF
C635 a_2407_49289# a_2315_44124# 0.39fF
C636 a_4259_73807# a_4583_68021# 0.55fF
C637 a_6664_26159# nmat.col[2] 0.79fF
C638 a_18546_24550# a_39154_24958# 0.35fF
C639 a_12447_16143# a_7415_29397# 0.49fF
C640 a_18162_9492# vcm 6.95fF
C641 a_48282_8488# m2_48052_7214# 1.00fF
C642 a_41254_61150# vcm 0.62fF
C643 a_39246_23548# m2_39016_24282# 0.99fF
C644 pmat.rowoff_n[15] a_18546_71232# 4.09fF
C645 VDD m3_18064_21402# 0.31fF
C646 a_18546_22542# a_36142_22950# 0.35fF
C647 pmat.en_bit_n[2] ANTENNA__1184__B1.DIODE 1.94fF
C648 nmat.en_bit_n[1] a_12851_28853# 0.40fF
C649 a_11067_27239# nmat.en_bit_n[0] 1.18fF
C650 a_38851_28327# a_45019_38645# 0.46fF
C651 VDD m2_41024_54946# 0.62fF
C652 VDD a_4955_40277# 2.65fF
C653 a_35230_20536# vcm 0.65fF
C654 a_31214_65166# a_32218_65166# 0.97fF
C655 VDD a_50290_22544# 0.54fF
C656 a_3339_70759# a_5805_49007# 0.59fF
C657 VDD a_44571_32143# 0.47fF
C658 VDD a_20078_7890# 0.33fF
C659 VDD a_26194_59142# 0.52fF
C660 a_38242_21540# a_39246_21540# 0.97fF
C661 VDD a_25755_34343# 0.92fF
C662 a_47278_17524# vcm 0.65fF
C663 a_18546_16518# a_22086_16926# 0.35fF
C664 m2_22952_54946# vcm 0.42fF
C665 pmat.rowon_n[8] a_11435_58791# 0.85fF
C666 a_2263_43719# a_1769_47919# 0.72fF
C667 ANTENNA__1190__A1.DIODE a_25695_28111# 0.35fF
C668 a_39246_71190# a_39246_70186# 1.00fF
C669 a_48282_8488# vcm 0.64fF
C670 a_18563_27791# a_37795_29111# 0.32fF
C671 pmat.rowon_n[7] nmat.rowoff_n[6] 1.08fF
C672 VDD a_32072_42919# 1.15fF
C673 nmat.col_n[29] nmat.col[17] 0.31fF
C674 a_20170_14512# a_21174_14512# 0.97fF
C675 m2_30984_7214# m2_31988_7214# 0.96fF
C676 _1154_.A _1194_.A2 1.02fF
C677 a_19166_64162# a_20170_64162# 0.97fF
C678 _1179_.X a_17139_30503# 1.10fF
C679 pmat.col_n[15] pmat.en_bit_n[1] 0.31fF
C680 a_17139_30503# a_33423_47695# 1.12fF
C681 a_2835_13077# a_11619_16367# 0.72fF
C682 VDD a_9301_69679# 0.61fF
C683 a_37238_13508# a_38242_13508# 0.97fF
C684 a_24186_15516# vcm 0.65fF
C685 a_19166_60146# ctopp 3.43fF
C686 a_35230_18528# a_36234_18528# 0.97fF
C687 a_12309_38659# a_11681_35823# 1.58fF
C688 a_24591_28327# a_26891_28327# 0.72fF
C689 pmat.row_n[14] vcm 1.28fF
C690 a_22178_62154# a_22178_61150# 1.00fF
C691 a_43262_12504# vcm 0.65fF
C692 a_48282_64162# ctopp 3.58fF
C693 a_2648_29397# a_4339_27804# 0.81fF
C694 nmat.col[28] vcm 8.86fF
C695 nmat.rowon_n[12] a_18162_11500# 1.33fF
C696 a_1781_9308# a_1979_11254# 0.31fF
C697 VDD a_26194_19532# 0.52fF
C698 a_22178_9492# ctopn 3.57fF
C699 a_6927_30503# a_1586_50247# 1.14fF
C700 VDD m2_26968_72014# 1.34fF
C701 nmat.rowon_n[1] a_14457_15823# 0.36fF
C702 a_14917_23983# a_13145_26935# 0.50fF
C703 a_20170_60146# vcm 0.62fF
C704 VDD a_25190_10496# 0.52fF
C705 pmat.row_n[15] a_7373_49007# 0.42fF
C706 a_1591_31599# a_2051_44111# 0.63fF
C707 VDD a_14773_39394# 1.64fF
C708 cgen.start_conv_in a_14600_37607# 0.59fF
C709 pmat.row_n[9] pmat.row_n[3] 0.41fF
C710 a_38242_20536# ctopn 3.58fF
C711 a_10515_13967# a_16083_50069# 0.38fF
C712 a_46274_15516# a_47278_15516# 0.97fF
C713 a_22178_15516# a_22178_14512# 1.00fF
C714 pmat.col_n[12] m2_30984_54946# 0.37fF
C715 nmat.sw a_11057_35836# 0.69fF
C716 a_6927_30503# a_3746_58487# 2.67fF
C717 a_18546_58180# a_32126_58138# 0.35fF
C718 a_45270_69182# a_46274_69182# 0.97fF
C719 a_24186_69182# a_24186_68178# 1.00fF
C720 VDD a_4471_30724# 0.77fF
C721 _1194_.B1 nmat.col[28] 0.30fF
C722 VDD a_4719_30287# 6.73fF
C723 a_12345_36924# cgen.dlycontrol1_in[0] 2.60fF
C724 a_18546_10494# a_32126_10902# 0.35fF
C725 a_32218_21540# a_32218_20536# 1.00fF
C726 VDD a_19689_34789# 1.26fF
C727 a_24591_28327# _1184_.A2 4.95fF
C728 ANTENNA__1395__A2.DIODE a_16311_28327# 2.22fF
C729 a_24867_53135# pmat.col[12] 0.34fF
C730 a_50290_17524# ctopn 3.43fF
C731 a_30111_47911# a_29076_48695# 0.45fF
C732 a_32218_62154# ctopp 3.58fF
C733 VDD a_41254_62154# 0.52fF
C734 a_26194_16520# vcm 0.65fF
C735 a_11149_40188# a_11041_39860# 1.58fF
C736 a_14839_66103# _1194_.B1 0.37fF
C737 a_1781_9308# a_2021_26677# 1.60fF
C738 VDD a_2847_23743# 0.36fF
C739 VDD a_44515_38645# 0.52fF
C740 VDD nmat.rowoff_n[2] 2.83fF
C741 pmat.sample pmat.row_n[12] 0.45fF
C742 ANTENNA__1197__A.DIODE a_15667_27239# 2.79fF
C743 a_2315_44124# a_4399_51157# 0.70fF
C744 a_18546_55168# a_33130_55126# 0.35fF
C745 a_18546_24550# a_21082_24958# 0.35fF
C746 a_10049_60663# a_10190_60663# 0.37fF
C747 m2_17932_64986# vcm 0.44fF
C748 a_31214_70186# ctopp 3.57fF
C749 a_27198_15516# ctopn 3.58fF
C750 VDD a_40250_70186# 0.52fF
C751 VDD a_27198_11500# 0.52fF
C752 pmat.rowon_n[0] a_4075_31591# 0.57fF
C753 a_14641_57711# pmat.rowon_n[7] 0.31fF
C754 a_43262_23548# a_43262_22544# 1.00fF
C755 a_19541_28879# a_7717_14735# 2.38fF
C756 ANTENNA__1197__B.DIODE a_8583_29199# 0.71fF
C757 _1179_.X a_26891_28327# 0.34fF
C758 a_47278_63158# pmat.col[28] 0.31fF
C759 pmat.row_n[0] ctopn 1.37fF
C760 a_42258_60146# a_43262_60146# 0.97fF
C761 a_46274_12504# ctopn 3.58fF
C762 a_18546_69224# a_27106_69182# 0.35fF
C763 a_11149_36924# a_11057_35836# 0.58fF
C764 pmat.row_n[4] a_18546_12502# 0.35fF
C765 a_26194_11500# a_26194_10496# 1.00fF
C766 a_42258_56130# vcm 0.62fF
C767 VDD a_30913_36603# 1.44fF
C768 a_18546_11498# vcm 0.40fF
C769 a_24591_28327# a_9411_2215# 5.55fF
C770 a_15101_29423# a_10441_21263# 1.44fF
C771 a_19166_59142# a_19166_58138# 1.00fF
C772 a_18546_63200# a_46182_63158# 0.35fF
C773 m2_40020_24282# m3_40152_24414# 2.79fF
C774 nmat.col[12] nmat.col_n[11] 6.90fF
C775 a_50290_68178# a_50290_67174# 1.00fF
C776 a_1823_58237# a_3496_51701# 0.44fF
C777 a_14287_69455# pmat.rowoff_n[2] 1.60fF
C778 a_24186_22544# vcm 0.65fF
C779 a_31214_61150# a_32218_61150# 0.97fF
C780 a_22178_68178# ctopp 3.58fF
C781 a_24867_53135# a_22199_30287# 0.60fF
C782 a_2835_13077# a_2199_13887# 1.03fF
C783 a_45270_66170# vcm 0.62fF
C784 VDD a_31214_68178# 0.52fF
C785 nmat.col_n[18] nmat.col[19] 6.82fF
C786 a_10767_39087# a_12585_40443# 1.18fF
C787 ANTENNA__1395__A1.DIODE nmat.en_bit_n[2] 0.33fF
C788 a_19166_66170# a_19166_65166# 1.00fF
C789 pmat.col_n[2] vcm 2.80fF
C790 pmat.row_n[8] ctopp 1.65fF
C791 VDD a_39013_43655# 1.67fF
C792 a_1923_53055# a_2676_51843# 0.63fF
C793 a_2199_13887# a_4075_13653# 0.40fF
C794 a_38242_63158# vcm 0.62fF
C795 VDD a_12723_64789# 0.50fF
C796 _1179_.X _1184_.A2 7.87fF
C797 a_13459_28111# ANTENNA__1195__A1.DIODE 0.64fF
C798 ANTENNA__1196__A2.DIODE a_16311_28327# 1.17fF
C799 a_14641_57167# a_10515_13967# 0.75fF
C800 a_25190_20536# a_26194_20536# 0.97fF
C801 a_18546_20534# a_33130_20942# 0.35fF
C802 VDD comp.adc_inverter_1.out 0.59fF
C803 a_29206_16520# ctopn 3.58fF
C804 pmat.rowoff_n[15] ctopp 0.42fF
C805 VDD pmat.sample_n 34.70fF
C806 a_5651_66975# a_5462_62215# 0.45fF
C807 a_48282_16520# a_49286_16520# 0.97fF
C808 a_38242_67174# a_38242_66170# 1.00fF
C809 a_24186_9492# a_24186_8488# 1.00fF
C810 VDD a_36234_23548# 0.54fF
C811 a_12309_38659# a_15049_36374# 1.05fF
C812 VDD a_38242_9492# 0.52fF
C813 a_1899_35051# a_2283_39189# 0.33fF
C814 VDD a_12925_60431# 0.46fF
C815 a_18546_11498# a_36142_11906# 0.35fF
C816 VDD a_16045_37692# 1.16fF
C817 a_30663_50087# a_40951_31599# 0.45fF
C818 a_4068_25615# a_6634_26133# 0.60fF
C819 pmat.rowoff_n[4] a_2263_43719# 0.59fF
C820 nmat.col[31] a_18563_27791# 1.69fF
C821 nmat.sw a_25325_29125# 0.37fF
C822 m2_31988_7214# m3_32120_7346# 2.79fF
C823 pmat.en_bit_n[2] a_13641_23439# 1.08fF
C824 nmat.en_bit_n[0] a_9785_28879# 2.97fF
C825 a_10223_26703# a_9217_23983# 0.47fF
C826 a_37238_17524# a_38242_17524# 0.97fF
C827 a_35230_57134# a_36234_57134# 0.97fF
C828 a_18162_69222# ctopp 1.49fF
C829 a_40250_20536# a_40250_19532# 1.00fF
C830 a_34226_71190# a_35230_71190# 0.97fF
C831 a_18546_71232# a_51202_71190# 0.35fF
C832 a_43262_67174# vcm 0.62fF
C833 a_12263_50959# a_11067_30287# 0.99fF
C834 a_18546_12502# a_20078_12910# 0.35fF
C835 nmat.en_bit_n[1] a_15667_28111# 3.06fF
C836 a_21174_58138# a_22178_58138# 0.97fF
C837 a_20170_20536# ctopn 3.57fF
C838 VDD config_1_in[7] 0.89fF
C839 VDD a_21032_44007# 1.22fF
C840 a_32218_14512# vcm 0.65fF
C841 VDD a_6679_15492# 0.54fF
C842 a_11067_27239# a_6664_26159# 0.39fF
C843 a_31214_64162# vcm 0.62fF
C844 _1196_.B1 a_12175_27221# 0.72fF
C845 a_38242_8488# a_39246_8488# 0.97fF
C846 VDD nmat.col[20] 4.51fF
C847 nmat.col_n[13] a_4383_7093# 0.91fF
C848 VDD a_30219_29967# 0.41fF
C849 _1179_.X a_9411_2215# 1.05fF
C850 a_2419_69455# pmat.row_n[4] 1.62fF
C851 VDD pmat.rowoff_n[1] 2.18fF
C852 a_19584_52423# a_11948_49783# 1.16fF
C853 cgen.dlycontrol1_in[4] a_11681_35823# 0.75fF
C854 a_11067_49871# a_20475_49783# 0.32fF
C855 m2_17932_62978# m2_17932_61974# 0.99fF
C856 VDD a_34226_13508# 0.52fF
C857 a_46274_14512# a_46274_13508# 1.00fF
C858 a_27198_22544# ctopn 3.57fF
C859 VDD a_32218_18528# 0.52fF
C860 m2_17932_21270# m3_18064_21402# 2.76fF
C861 m2_46044_54946# vcm 0.42fF
C862 VDD m2_51064_66994# 1.02fF
C863 ANTENNA__1190__A2.DIODE a_3688_17179# 0.65fF
C864 a_50290_57134# a_50290_56130# 1.00fF
C865 a_21174_61150# a_21174_60146# 1.00fF
C866 a_6830_22895# a_11927_27399# 0.46fF
C867 _1184_.A2 a_4976_16091# 0.32fF
C868 a_29206_19532# a_29206_18528# 1.00fF
C869 VDD a_1823_60949# 2.00fF
C870 pmat.row_n[2] a_14457_15823# 0.62fF
C871 a_7109_29423# a_18597_31599# 11.90fF
C872 VDD a_4984_41935# 0.36fF
C873 VDD a_43262_15516# 0.52fF
C874 a_18546_14510# a_34134_14918# 0.35fF
C875 nmat.col[7] nmat.rowon_n[6] 0.40fF
C876 a_17139_30503# nmat.col[7] 0.72fF
C877 pmat.rowoff_n[15] a_5351_19913# 0.40fF
C878 a_18546_64204# a_32126_64162# 0.35fF
C879 a_10239_14183# a_13091_18535# 0.70fF
C880 cgen.dlycontrol4_in[3] a_2563_34837# 0.43fF
C881 a_22178_59142# a_22178_58138# 1.00fF
C882 a_11067_27239# a_27763_27221# 5.35fF
C883 a_19166_13508# a_19166_12504# 1.00fF
C884 VDD a_12449_22895# 2.26fF
C885 VDD m3_18064_72146# 0.33fF
C886 pmat.col_n[1] ANTENNA__1195__A1.DIODE 0.83fF
C887 a_34226_65166# vcm 0.62fF
C888 nmat.col[0] vcm 5.74fF
C889 a_41254_21540# vcm 0.65fF
C890 a_30210_60146# ctopp 3.58fF
C891 m2_23956_72014# m3_24088_72146# 2.79fF
C892 a_30210_62154# pmat.col[11] 0.31fF
C893 ANTENNA__1183__B1.DIODE vcm 3.51fF
C894 VDD a_39246_60146# 0.52fF
C895 a_2952_25045# a_4516_21531# 0.39fF
C896 a_4339_27804# a_4068_25615# 1.15fF
C897 VDD a_26331_36919# 0.63fF
C898 VDD a_11014_71855# 0.47fF
C899 nmat.col[25] vcm 5.76fF
C900 a_27198_17524# a_27198_16520# 1.00fF
C901 m2_49056_54946# m3_49188_55078# 2.79fF
C902 _1192_.A2 nmat.col[26] 2.29fF
C903 a_18546_19530# a_45178_19938# 0.35fF
C904 m2_31988_54946# m2_32992_54946# 0.96fF
C905 a_35230_14512# ctopn 3.58fF
C906 VDD a_13718_68591# 0.38fF
C907 a_33222_12504# a_34226_12504# 0.97fF
C908 a_18546_12502# a_49194_12910# 0.35fF
C909 pmat.rowon_n[8] pmat.row_n[9] 0.46fF
C910 cgen.dlycontrol4_in[5] cgen.dlycontrol1_in[1] 0.47fF
C911 a_46274_22544# a_47278_22544# 0.97fF
C912 VDD a_45270_16520# 0.52fF
C913 _1194_.B1 ANTENNA__1183__B1.DIODE 3.10fF
C914 VDD m2_17932_21270# 1.11fF
C915 a_11067_30287# clk_ena 2.82fF
C916 VDD a_19831_51316# 0.45fF
C917 pmat.rowon_n[3] pmat.rowoff_n[3] 20.32fF
C918 a_22178_59142# a_23182_59142# 0.97fF
C919 a_18546_59184# a_27106_59142# 0.35fF
C920 a_3339_70759# a_2935_38279# 0.42fF
C921 a_35244_32411# a_25575_31055# 0.55fF
C922 a_23182_57134# ctopp 3.57fF
C923 a_22178_71190# ctopp 3.40fF
C924 VDD a_32218_57134# 0.52fF
C925 _1154_.X a_22307_27791# 0.34fF
C926 a_48282_69182# vcm 0.62fF
C927 VDD a_31214_71190# 0.55fF
C928 VDD a_8013_73493# 0.71fF
C929 cgen.dlycontrol4_in[0] cgen.dlycontrol4_in[1] 4.33fF
C930 VDD vcm.sky130_fd_sc_hd__dlymetal6s6s_1_3.X 0.49fF
C931 a_3615_71631# a_13432_62581# 1.25fF
C932 VDD a_20170_9492# 0.52fF
C933 VDD a_28189_37981# 1.33fF
C934 VDD a_11113_40835# 8.16fF
C935 a_23182_56130# m2_22952_54946# 0.99fF
C936 a_34705_51959# pmat.col[16] 0.33fF
C937 a_7415_29397# a_6829_26703# 0.36fF
C938 a_18546_55168# a_43170_55126# 0.35fF
C939 a_18546_24550# a_32126_24958# 0.35fF
C940 a_12079_31061# a_5535_29980# 0.33fF
C941 a_20605_40719# a_21219_36885# 0.44fF
C942 inp_analog _1187_.A2 2.51fF
C943 nmat.sw nmat.col_n[19] 0.69fF
C944 a_41731_49525# nmat.col[31] 0.42fF
C945 a_34226_61150# vcm 0.62fF
C946 a_18546_72236# a_50198_72194# 0.35fF
C947 a_10223_26703# nmat.col[3] 0.58fF
C948 a_18546_22542# a_29114_22950# 0.35fF
C949 a_2411_33749# a_1591_38677# 0.34fF
C950 a_44266_21540# ctopn 3.58fF
C951 VDD a_4700_44655# 0.36fF
C952 cgen.start_conv_in a_10873_40693# 1.41fF
C953 VDD a_7840_27247# 1.98fF
C954 a_28202_20536# vcm 0.65fF
C955 VDD a_43262_22544# 0.52fF
C956 pmat.row_n[10] nmat.sample 0.35fF
C957 pmat.col_n[10] ctopp 2.02fF
C958 a_12069_36341# a_13779_36595# 0.72fF
C959 VDD a_13319_35507# 1.06fF
C960 VDD a_36142_72194# 0.32fF
C961 VDD a_4895_12559# 0.57fF
C962 a_48282_63158# ctopp 3.58fF
C963 pmat.col_n[2] pmat.col[2] 0.82fF
C964 a_40250_17524# vcm 0.65fF
C965 VDD a_12337_18005# 0.44fF
C966 a_4516_21531# a_2683_22089# 0.69fF
C967 a_11497_38543# a_12197_38306# 0.65fF
C968 pmat.rowoff_n[0] a_18546_56172# 4.09fF
C969 a_9135_60967# a_11007_58229# 0.99fF
C970 m2_28976_24282# m2_29980_24282# 0.96fF
C971 a_41254_8488# vcm 0.64fF
C972 nmat.col[14] m2_32992_24282# 0.39fF
C973 a_20438_35431# a_10873_36341# 0.49fF
C974 a_32687_46607# a_37291_29397# 0.36fF
C975 VDD a_12658_42895# 1.03fF
C976 m2_23956_7214# m2_24960_7214# 0.96fF
C977 ANTENNA__1197__A.DIODE a_11067_27239# 5.21fF
C978 _1194_.A2 nmat.en_bit_n[1] 0.59fF
C979 a_49286_18528# a_49286_17524# 1.00fF
C980 a_2149_45717# a_2983_48071# 1.38fF
C981 VDD a_41321_30511# 0.38fF
C982 VDD a_10595_53361# 0.91fF
C983 a_18546_13506# a_50198_13914# 0.35fF
C984 VDD a_1591_27797# 0.40fF
C985 pmat.row_n[12] a_18162_20536# 25.57fF
C986 VDD a_11023_76359# 0.56fF
C987 a_49286_63158# a_49286_62154# 1.00fF
C988 a_18546_18526# a_46182_18934# 0.35fF
C989 a_25190_70186# a_25190_69182# 1.00fF
C990 VDD a_4523_21276# 6.03fF
C991 a_12437_28879# a_17306_28879# 0.46fF
C992 a_21219_36885# a_22111_36950# 0.31fF
C993 VDD a_43533_30761# 3.31fF
C994 a_36234_12504# vcm 0.65fF
C995 a_41254_64162# ctopp 3.58fF
C996 a_24407_31375# a_34204_27765# 0.39fF
C997 VDD a_50290_64162# 0.56fF
C998 a_34226_24552# a_35230_24552# 0.97fF
C999 ANTENNA__1190__A1.DIODE comp_latch 0.31fF
C1000 pmat.col[30] vcm 5.88fF
C1001 a_10055_31591# pmat.rowoff_n[4] 1.43fF
C1002 pmat.sample a_18547_51565# 1.13fF
C1003 nmat.col_n[13] a_9075_28023# 0.74fF
C1004 a_22178_19532# a_23182_19532# 0.97fF
C1005 pmat.en_bit_n[2] a_13091_28327# 0.44fF
C1006 VDD a_22499_49783# 2.53fF
C1007 a_48282_13508# a_48282_12504# 1.00fF
C1008 cgen.start_conv_in a_13357_37429# 0.87fF
C1009 a_31214_20536# ctopn 3.58fF
C1010 pmat.col_n[8] m2_26968_54946# 0.37fF
C1011 VDD m2_18936_23278# 0.57fF
C1012 a_2007_25597# a_32771_31599# 0.37fF
C1013 pmat.rowon_n[3] a_18162_59182# 1.19fF
C1014 a_18546_58180# a_25098_58138# 0.35fF
C1015 VDD a_8583_29199# 8.24fF
C1016 _1224_.X pmat.col[6] 0.34fF
C1017 a_18546_10494# a_25098_10902# 0.35fF
C1018 a_21174_10496# a_22178_10496# 0.97fF
C1019 VDD a_12561_57167# 0.40fF
C1020 a_43262_17524# ctopn 3.58fF
C1021 a_25190_62154# ctopp 3.58fF
C1022 VDD a_34226_62154# 0.52fF
C1023 a_11067_64015# clk_ena 0.39fF
C1024 a_18162_16520# vcm 6.95fF
C1025 a_44266_8488# ctopn 3.40fF
C1026 a_32218_56130# a_33222_56130# 0.97fF
C1027 a_18546_56172# a_47186_56130# 0.35fF
C1028 VDD a_46182_24958# 0.44fF
C1029 VDD a_46897_40303# 0.54fF
C1030 pmat.rowon_n[15] vcm 0.59fF
C1031 a_44266_65166# ctopp 3.58fF
C1032 ANTENNA__1395__A1.DIODE a_24407_31375# 0.31fF
C1033 VDD a_10167_64239# 0.37fF
C1034 a_18546_55168# a_26102_55126# 0.35fF
C1035 a_21371_50087# a_33957_48437# 0.48fF
C1036 VDD a_14471_20175# 0.42fF
C1037 a_19166_17524# a_20170_17524# 0.97fF
C1038 ANTENNA__1395__B1.DIODE nmat.col[29] 0.87fF
C1039 a_9545_66567# a_9405_66627# 0.81fF
C1040 a_24186_70186# ctopp 3.57fF
C1041 VDD a_33222_70186# 0.52fF
C1042 a_22178_23548# m2_21948_24282# 0.99fF
C1043 a_13091_28327# a_5363_33551# 0.64fF
C1044 a_22178_63158# pmat.col[3] 0.31fF
C1045 a_44266_16520# a_44266_15516# 1.00fF
C1046 a_19166_15516# a_20170_15516# 0.97fF
C1047 a_37238_62154# a_38242_62154# 0.97fF
C1048 a_35230_66170# a_36234_66170# 0.97fF
C1049 a_39246_12504# ctopn 3.58fF
C1050 a_12237_36596# a_13779_36595# 0.77fF
C1051 a_35230_56130# vcm 0.62fF
C1052 pmat.rowon_n[0] cgen.dlycontrol2_in[4] 0.97fF
C1053 a_1586_63927# a_2215_47375# 0.54fF
C1054 VDD pmat.col_n[3] 6.18fF
C1055 pmat.rowoff_n[7] a_12447_16143# 2.21fF
C1056 a_18546_63200# a_39154_63158# 0.35fF
C1057 a_28202_63158# a_29206_63158# 0.97fF
C1058 VDD m2_17932_70006# 1.00fF
C1059 VDD a_1895_23610# 0.58fF
C1060 pmat.rowon_n[7] a_15899_47939# 1.57fF
C1061 a_38242_66170# vcm 0.62fF
C1062 VDD a_24186_68178# 0.52fF
C1063 pmat.en_bit_n[2] a_17139_30503# 0.51fF
C1064 m2_48052_72014# m2_49056_72014# 0.96fF
C1065 cgen.start_conv_in a_12934_35823# 0.36fF
C1066 a_31214_63158# vcm 0.62fF
C1067 VDD a_4128_64391# 7.99fF
C1068 a_1591_63701# a_1757_63701# 0.72fF
C1069 VDD a_45178_55126# 0.42fF
C1070 VDD a_24959_31055# 0.31fF
C1071 a_10873_36341# cgen.dlycontrol1_in[0] 0.36fF
C1072 a_18546_20534# a_26102_20942# 0.35fF
C1073 a_22178_16520# ctopn 3.58fF
C1074 VDD m2_17932_9222# 1.00fF
C1075 a_18243_28327# a_35244_32411# 0.46fF
C1076 a_2263_43719# a_33986_47375# 0.31fF
C1077 nmat.col[31] vcm 5.49fF
C1078 VDD a_5411_48695# 0.53fF
C1079 a_3727_66113# a_3688_65987# 0.72fF
C1080 VDD a_29206_23548# 0.55fF
C1081 a_44266_61150# ctopp 3.58fF
C1082 a_36234_70186# a_37238_70186# 0.97fF
C1083 ANTENNA__1187__B1.DIODE a_34705_51959# 0.48fF
C1084 a_24867_53135# a_34942_51701# 0.73fF
C1085 VDD a_31214_9492# 0.52fF
C1086 a_12513_36924# a_12585_37179# 0.78fF
C1087 a_18547_51565# a_18823_50247# 1.43fF
C1088 a_18546_11498# a_29114_11906# 0.35fF
C1089 a_23182_11500# a_24186_11500# 0.97fF
C1090 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top comp.adc_inverter_1.in 0.40fF
C1091 pmat.sample_n a_22499_49783# 1.74fF
C1092 VDD a_20811_41271# 0.60fF
C1093 nmat.col[13] nmat.col[7] 4.15fF
C1094 a_17842_27497# a_34204_27765# 0.37fF
C1095 nmat.col_n[18] nmat.col_n[29] 1.20fF
C1096 nmat.col_n[30] nmat.col_n[19] 3.92fF
C1097 a_45019_38645# a_46229_37583# 0.44fF
C1098 VDD a_47278_20536# 0.52fF
C1099 a_25190_64162# a_25190_63158# 1.00fF
C1100 VDD a_22541_39867# 1.39fF
C1101 pmat.row_n[14] ANTENNA__1190__A1.DIODE 0.48fF
C1102 a_28202_10496# a_28202_9492# 1.00fF
C1103 cgen.dlycontrol1_in[0] cgen.dlycontrol1_in[3] 2.08fF
C1104 a_18546_71232# a_44174_71190# 0.35fF
C1105 a_36234_67174# vcm 0.62fF
C1106 a_25190_58138# a_25190_57134# 1.00fF
C1107 _1196_.B1 ANTENNA__1197__A.DIODE 1.56fF
C1108 nmat.sample_n nmat.col[13] 6.21fF
C1109 _1194_.A2 a_19584_52423# 0.63fF
C1110 _1187_.A2 ANTENNA__1395__B1.DIODE 0.63fF
C1111 _1194_.B1 a_21739_29415# 0.64fF
C1112 a_5363_33551# a_17139_30503# 0.76fF
C1113 a_31675_47695# a_45277_32687# 0.37fF
C1114 VDD cgen.dlycontrol4_in[4] 6.18fF
C1115 a_25190_14512# vcm 0.65fF
C1116 a_4719_30287# a_5411_48695# 0.64fF
C1117 a_12447_16143# a_11067_30287# 1.40fF
C1118 ANTENNA__1187__B1.DIODE nmat.col[10] 2.95fF
C1119 a_24186_64162# vcm 0.62fF
C1120 a_29206_60146# a_29206_59142# 1.00fF
C1121 a_18546_65208# a_49194_65166# 0.35fF
C1122 a_4075_68583# a_4243_54991# 0.90fF
C1123 a_35244_32411# a_28704_29568# 0.32fF
C1124 m2_51064_70006# m3_51196_70138# 2.76fF
C1125 a_14773_37218# cgen.dlycontrol1_in[1] 1.04fF
C1126 a_6927_30503# a_4259_31375# 1.04fF
C1127 a_47278_62154# a_47278_61150# 1.00fF
C1128 VDD a_27198_13508# 0.52fF
C1129 _1154_.A ANTENNA__1197__B.DIODE 0.52fF
C1130 VDD a_25190_18528# 0.52fF
C1131 a_33222_67174# a_34226_67174# 0.97fF
C1132 a_18546_67216# a_49194_67174# 0.35fF
C1133 a_2648_29397# a_2191_25045# 0.35fF
C1134 VDD a_2124_67771# 0.65fF
C1135 VDD nmat.col_n[2] 5.34fF
C1136 VDD a_2124_61635# 0.56fF
C1137 a_23182_22544# a_23182_21540# 1.00fF
C1138 a_30210_66170# a_30210_65166# 1.00fF
C1139 a_18823_50247# a_11948_49783# 0.83fF
C1140 a_18546_13506# vcm 0.40fF
C1141 VDD a_36234_15516# 0.52fF
C1142 a_47278_15516# a_47278_14512# 1.00fF
C1143 a_22178_14512# a_23182_14512# 0.97fF
C1144 a_18546_14510# a_27106_14918# 0.35fF
C1145 m2_51064_16250# vcm 0.51fF
C1146 a_18546_7482# a_49194_7890# 0.35fF
C1147 a_21174_64162# a_22178_64162# 0.97fF
C1148 a_18546_64204# a_25098_64162# 0.35fF
C1149 pmat.row_n[0] a_18162_8488# 25.57fF
C1150 pmat.row_n[0] ctopp 1.39fF
C1151 a_49286_69182# a_49286_68178# 1.00fF
C1152 a_27198_68178# a_28202_68178# 0.97fF
C1153 a_3339_59879# a_11271_73085# 0.32fF
C1154 a_2046_30184# a_1923_31743# 0.86fF
C1155 pmat.row_n[15] pmat.rowon_n[0] 1.49fF
C1156 a_7663_71317# a_7829_71317# 0.70fF
C1157 a_12449_22895# a_4523_21276# 0.45fF
C1158 _1194_.B1 a_40105_47375# 0.62fF
C1159 VDD m2_39016_7214# 1.31fF
C1160 pmat.col[14] ctopp 1.98fF
C1161 a_27198_65166# vcm 0.62fF
C1162 VDD a_41663_47893# 0.43fF
C1163 a_34226_21540# vcm 0.65fF
C1164 VDD a_3305_15823# 4.72fF
C1165 a_23182_60146# ctopp 3.58fF
C1166 nmat.rowon_n[7] nmat.rowon_n[12] 1.23fF
C1167 VDD a_2787_33237# 0.44fF
C1168 VDD a_32218_60146# 0.52fF
C1169 a_31263_28309# a_21365_27247# 0.39fF
C1170 a_49286_58138# vcm 0.62fF
C1171 a_19166_63158# a_20170_63158# 0.97fF
C1172 a_14653_53458# ANTENNA__1395__A1.DIODE 0.46fF
C1173 a_18546_19530# a_38150_19938# 0.35fF
C1174 m2_24960_54946# m2_25964_54946# 0.96fF
C1175 a_38851_28327# a_47207_35951# 0.35fF
C1176 a_28202_14512# ctopn 3.58fF
C1177 pmat.en_bit_n[2] _1184_.A2 0.75fF
C1178 a_2879_57487# a_3967_56311# 0.40fF
C1179 a_1586_50247# cgen.dlycontrol3_in[4] 0.51fF
C1180 a_18546_12502# a_42166_12910# 0.35fF
C1181 a_27198_63158# pmat.col[8] 0.31fF
C1182 VDD a_28631_44265# 0.64fF
C1183 VDD a_38242_16520# 0.52fF
C1184 pmat.rowon_n[0] a_6283_31591# 1.22fF
C1185 a_23182_65166# a_23182_64162# 1.00fF
C1186 m2_51064_66994# m3_51196_67126# 2.76fF
C1187 nmat.sw a_7165_13353# 0.42fF
C1188 VDD a_28110_55126# 0.42fF
C1189 VDD a_48190_7890# 0.33fF
C1190 VDD a_9305_58229# 0.60fF
C1191 _1154_.X nmat.col[31] 1.33fF
C1192 VDD a_25190_57134# 0.52fF
C1193 _1154_.X a_21739_29415# 0.68fF
C1194 a_41254_69182# vcm 0.62fF
C1195 VDD a_24186_71190# 0.55fF
C1196 ANTENNA__1184__B1.DIODE a_15667_27239# 0.32fF
C1197 nmat.col[0] nmat.col_n[0] 0.75fF
C1198 a_32218_23548# a_33222_23548# 0.97fF
C1199 a_18546_23546# a_47186_23954# 0.35fF
C1200 cgen.dlycontrol4_in[4] a_39013_43655# 0.45fF
C1201 a_25190_71190# m2_24960_72014# 1.00fF
C1202 a_34226_9492# a_35230_9492# 0.97fF
C1203 a_18546_9490# a_51202_9898# 0.35fF
C1204 VDD a_3325_36495# 1.32fF
C1205 a_50290_59142# vcm 0.62fF
C1206 a_2389_45859# nmat.rowon_n[14] 0.65fF
C1207 VDD a_26460_40517# 1.19fF
C1208 a_9463_50877# a_9427_50095# 0.59fF
C1209 a_41254_12504# a_41254_11500# 1.00fF
C1210 a_18546_55168# a_36142_55126# 0.39fF
C1211 a_18546_24550# a_25098_24958# 0.35fF
C1212 a_45270_56130# ctopp 3.40fF
C1213 ANTENNA_fanout52_A.DIODE a_29937_31055# 0.35fF
C1214 VDD a_10955_55687# 0.42fF
C1215 a_26891_28327# a_28336_29967# 1.55fF
C1216 a_6200_70919# a_6051_74183# 0.39fF
C1217 a_27198_61150# vcm 0.62fF
C1218 a_2419_69455# a_4025_54965# 0.72fF
C1219 a_18546_22542# a_22086_22950# 0.35fF
C1220 a_37238_21540# ctopn 3.58fF
C1221 pmat.col_n[25] pmat.col[25] 1.02fF
C1222 a_2407_49289# a_2419_53351# 0.46fF
C1223 VDD a_28639_47081# 0.59fF
C1224 a_21174_20536# vcm 0.65fF
C1225 a_49286_9492# a_49286_8488# 1.00fF
C1226 VDD a_5725_76207# 0.69fF
C1227 a_24186_65166# a_25190_65166# 0.97fF
C1228 VDD a_36234_22544# 0.52fF
C1229 a_48282_66170# ctopp 3.58fF
C1230 a_2835_13077# a_11711_12565# 0.34fF
C1231 VDD a_18241_31698# 5.66fF
C1232 VDD a_2163_58941# 0.52fF
C1233 a_31214_21540# a_32218_21540# 0.97fF
C1234 _1184_.A2 a_10513_24135# 0.43fF
C1235 a_11067_64015# a_12447_16143# 0.88fF
C1236 a_41254_63158# ctopp 3.58fF
C1237 a_30571_50959# a_35244_32411# 1.02fF
C1238 VDD a_50290_63158# 0.54fF
C1239 a_33222_17524# vcm 0.65fF
C1240 a_1586_8439# config_1_in[8] 0.48fF
C1241 m2_45040_24282# m3_45172_24414# 2.79fF
C1242 a_25695_28111# a_40903_32375# 0.96fF
C1243 a_18546_61192# a_49194_61150# 0.35fF
C1244 VDD a_19074_24958# 0.44fF
C1245 a_24591_28327# a_25879_31591# 0.57fF
C1246 ANTENNA__1187__B1.DIODE _1183_.A2 0.85fF
C1247 VDD config_2_in[11] 1.15fF
C1248 nmat.sw a_10781_42869# 0.64fF
C1249 m2_21948_24282# m2_22952_24282# 0.96fF
C1250 a_32218_71190# a_32218_70186# 1.00fF
C1251 a_34226_8488# vcm 0.64fF
C1252 pmat.col_n[5] vcm 2.80fF
C1253 a_46274_58138# a_47278_58138# 0.97fF
C1254 a_2648_29397# a_8243_7290# 0.32fF
C1255 a_50290_19532# vcm 0.65fF
C1256 m2_51064_63982# m3_51196_64114# 2.76fF
C1257 a_18546_68220# a_19074_68178# 0.35fF
C1258 pmat.rowon_n[12] a_18162_68218# 1.19fF
C1259 a_49286_10496# vcm 0.65fF
C1260 VDD result_out[5] 0.58fF
C1261 a_30210_13508# a_31214_13508# 0.97fF
C1262 a_18546_13506# a_43170_13914# 0.35fF
C1263 a_10781_42869# a_15049_42902# 0.56fF
C1264 pmat.sw a_24747_29967# 1.00fF
C1265 a_44266_71190# m2_44036_72014# 1.00fF
C1266 VDD a_40949_48437# 0.86fF
C1267 a_46274_61150# a_46274_60146# 1.00fF
C1268 a_46274_67174# ctopp 3.58fF
C1269 a_28202_18528# a_29206_18528# 0.97fF
C1270 a_18546_18526# a_39154_18934# 0.35fF
C1271 m2_17932_17254# vcm 0.44fF
C1272 a_10190_60663# a_9135_60967# 0.33fF
C1273 pmat.col_n[15] pmat.col[16] 6.25fF
C1274 a_29206_12504# vcm 0.65fF
C1275 a_34226_64162# ctopp 3.58fF
C1276 VDD a_44266_14512# 0.52fF
C1277 m2_37008_7214# m3_37140_7346# 2.79fF
C1278 nmat.sw a_20439_27247# 0.65fF
C1279 VDD a_43262_64162# 0.52fF
C1280 pmat.rowoff_n[12] a_1739_47893# 0.50fF
C1281 a_47278_59142# a_47278_58138# 1.00fF
C1282 a_33423_47695# a_36532_46805# 0.51fF
C1283 ANTENNA__1184__B1.DIODE a_14943_26703# 0.57fF
C1284 a_24186_20536# ctopn 3.58fF
C1285 VDD a_31097_44581# 1.35fF
C1286 VDD a_20170_16520# 0.52fF
C1287 a_39246_15516# a_40250_15516# 0.97fF
C1288 pmat.col_n[4] m2_22952_54946# 0.37fF
C1289 _1196_.B1 a_45112_47607# 0.47fF
C1290 VDD a_41949_30761# 0.82fF
C1291 a_38242_69182# a_39246_69182# 0.97fF
C1292 a_25190_21540# a_25190_20536# 1.00fF
C1293 a_36234_17524# ctopn 3.58fF
C1294 pmat.row_n[15] a_4075_31591# 0.92fF
C1295 VDD a_27198_62154# 0.52fF
C1296 _1179_.X a_25879_31591# 0.32fF
C1297 cgen.dlycontrol4_in[3] cgen.dlycontrol4_in[1] 2.15fF
C1298 a_14839_20871# a_13768_22325# 0.67fF
C1299 a_17139_30503# a_44774_40821# 0.45fF
C1300 a_37238_8488# ctopn 3.40fF
C1301 nmat.rowon_n[7] ANTENNA__1196__A2.DIODE 0.39fF
C1302 pmat.rowoff_n[8] pmat.rowon_n[8] 21.01fF
C1303 a_18546_56172# a_40158_56130# 0.35fF
C1304 VDD a_39154_24958# 0.44fF
C1305 pmat.sample _1194_.A2 0.54fF
C1306 a_10515_15055# a_10515_13967# 0.61fF
C1307 a_10515_61839# a_10878_58487# 0.36fF
C1308 a_37238_65166# ctopp 3.58fF
C1309 a_2407_49289# a_2419_69455# 1.89fF
C1310 a_18162_62194# vcm 6.95fF
C1311 VDD a_46274_65166# 0.52fF
C1312 a_18546_55168# a_19074_55126# 0.35fF
C1313 a_38851_28327# a_41731_49525# 3.15fF
C1314 a_47278_59142# a_48282_59142# 0.97fF
C1315 m2_51064_60970# m3_51196_61102# 2.76fF
C1316 a_37238_62154# pmat.col[18] 0.31fF
C1317 a_18546_68220# a_48190_68178# 0.35fF
C1318 cgen.dlycontrol3_in[3] cgen.dlycontrol4_in[5] 0.35fF
C1319 a_1923_69823# a_2695_76757# 0.58fF
C1320 VDD a_26194_70186# 0.52fF
C1321 a_36234_23548# a_36234_22544# 1.00fF
C1322 a_10239_14183# a_10839_11989# 0.32fF
C1323 a_19166_21540# ctopn 3.42fF
C1324 a_24591_28327# nmat.col_n[9] 0.35fF
C1325 a_11435_58791# _1192_.A2 0.34fF
C1326 a_10781_42869# a_12116_40871# 0.82fF
C1327 a_11113_39747# cgen.dlycontrol2_in[3] 7.24fF
C1328 a_4351_55527# a_3866_57399# 0.72fF
C1329 VDD pmat.col[7] 4.82fF
C1330 a_4259_31375# a_6979_51157# 0.74fF
C1331 a_35230_60146# a_36234_60146# 0.97fF
C1332 m2_28976_72014# m3_29108_72146# 2.79fF
C1333 a_4075_31591# a_6283_31591# 0.70fF
C1334 a_32218_12504# ctopn 3.58fF
C1335 VDD a_45277_32687# 0.76fF
C1336 _1183_.A2 nmat.rowon_n[5] 1.08fF
C1337 _1192_.B1 nmat.col[29] 0.63fF
C1338 a_28202_56130# vcm 0.62fF
C1339 VDD a_8231_72105# 0.38fF
C1340 VDD a_8735_54207# 0.37fF
C1341 a_12309_38659# ndecision_finish 2.58fF
C1342 a_18563_27791# a_37827_30793# 1.52fF
C1343 pmat.row_n[13] nmat.rowon_n[2] 20.77fF
C1344 a_18546_63200# a_32126_63158# 0.35fF
C1345 pmat.rowon_n[0] a_2648_29397# 0.47fF
C1346 pmat.row_n[3] ctopn 1.65fF
C1347 a_43262_68178# a_43262_67174# 1.00fF
C1348 a_24186_61150# a_25190_61150# 0.97fF
C1349 a_31214_66170# vcm 0.62fF
C1350 a_15667_27239# a_13641_23439# 0.70fF
C1351 m2_41024_72014# m2_42028_72014# 0.96fF
C1352 a_11067_64015# a_11435_58791# 0.86fF
C1353 VDD a_13503_43421# 1.43fF
C1354 a_24186_63158# vcm 0.62fF
C1355 a_26891_28327# nmat.col_n[18] 1.25fF
C1356 VDD a_38150_55126# 0.42fF
C1357 VDD m2_51064_19262# 1.03fF
C1358 pmat.rowoff_n[12] cgen.dlycontrol4_in[0] 0.66fF
C1359 VDD a_19166_12504# 0.56fF
C1360 VDD a_1591_71855# 1.25fF
C1361 a_6829_26703# a_8831_24501# 0.46fF
C1362 a_41254_16520# a_42258_16520# 0.97fF
C1363 VDD nmat.col[15] 11.97fF
C1364 a_31214_67174# a_31214_66170# 1.00fF
C1365 VDD _1154_.A 17.74fF
C1366 VDD a_22178_23548# 0.55fF
C1367 VDD a_33341_38780# 1.16fF
C1368 a_37238_61150# ctopp 3.58fF
C1369 a_18546_18526# a_21082_18934# 0.35fF
C1370 VDD a_24186_9492# 0.52fF
C1371 VDD a_46274_61150# 0.52fF
C1372 a_18546_11498# a_22086_11906# 0.35fF
C1373 VDD a_36341_38053# 1.20fF
C1374 VDD a_40250_20536# 0.52fF
C1375 a_30210_17524# a_31214_17524# 0.97fF
C1376 m2_51064_57958# m3_51196_58090# 2.76fF
C1377 pmat.rowon_n[0] pmat.rowoff_n[2] 0.72fF
C1378 a_28202_57134# a_29206_57134# 0.97fF
C1379 a_24861_29673# clk_ena 0.79fF
C1380 a_33222_20536# a_33222_19532# 1.00fF
C1381 m2_51064_57958# m2_51064_56954# 0.99fF
C1382 a_27198_71190# a_28202_71190# 0.97fF
C1383 a_18546_71232# a_37146_71190# 0.35fF
C1384 a_29206_67174# vcm 0.62fF
C1385 a_44444_32233# a_46523_39733# 0.41fF
C1386 pmat.row_n[14] pmat.row_n[5] 5.34fF
C1387 pmat.rowoff_n[8] pmat.row_n[7] 1.23fF
C1388 a_37820_30485# a_25575_31055# 0.98fF
C1389 pmat.col_n[23] pmat.col[24] 5.99fF
C1390 VDD a_19439_28585# 0.39fF
C1391 a_1739_47893# a_1858_25615# 1.23fF
C1392 VDD m2_32992_54946# 0.61fF
C1393 a_22199_30287# a_16478_29423# 0.92fF
C1394 a_31214_8488# a_32218_8488# 0.97fF
C1395 a_18546_8486# a_45178_8894# 0.35fF
C1396 a_18546_65208# a_42166_65166# 0.35fF
C1397 a_50290_70186# a_50290_69182# 1.00fF
C1398 VDD a_3551_6202# 0.82fF
C1399 a_3325_26159# a_3325_23439# 0.69fF
C1400 pmat.col_n[13] ctopp 2.02fF
C1401 a_7644_16341# a_4976_16091# 0.38fF
C1402 VDD a_20811_35831# 0.60fF
C1403 pmat.rowon_n[8] a_10239_14183# 1.54fF
C1404 VDD a_39154_72194# 0.33fF
C1405 a_39246_14512# a_39246_13508# 1.00fF
C1406 VDD a_11711_50959# 9.01fF
C1407 VDD a_12429_62607# 0.80fF
C1408 a_12693_38543# a_10927_37981# 0.37fF
C1409 ANTENNA__1197__B.DIODE nmat.en_bit_n[1] 0.68fF
C1410 ANTENNA__1187__B1.DIODE ANTENNA__1395__A2.DIODE 0.45fF
C1411 ANTENNA__1184__B1.DIODE a_11067_27239# 1.39fF
C1412 _1187_.A2 _1192_.B1 1.29fF
C1413 a_18546_67216# a_42166_67174# 0.35fF
C1414 a_43262_57134# a_43262_56130# 1.00fF
C1415 pmat.row_n[10] pmat.row_n[3] 0.58fF
C1416 VDD a_21082_24958# 0.44fF
C1417 a_13091_18535# a_5351_19913# 0.44fF
C1418 a_47278_19532# a_48282_19532# 0.97fF
C1419 a_22178_19532# a_22178_18528# 1.00fF
C1420 a_40105_47375# a_40837_46261# 0.39fF
C1421 pmat.row_n[6] nmat.en_bit_n[1] 0.51fF
C1422 nmat.col_n[12] nmat.col[13] 6.94fF
C1423 VDD a_9463_53511# 1.12fF
C1424 a_2839_38101# a_2743_38279# 0.37fF
C1425 a_19166_65166# ctopp 3.43fF
C1426 VDD a_23700_42919# 1.22fF
C1427 VDD a_29206_15516# 0.52fF
C1428 nmat.col[21] nmat.col_n[24] 4.77fF
C1429 a_1823_74557# a_2163_69821# 0.40fF
C1430 a_18546_14510# a_19074_14918# 0.35fF
C1431 a_7717_14735# a_15101_29423# 0.62fF
C1432 a_18546_7482# a_42166_7890# 0.35fF
C1433 a_23395_53135# _1187_.A2 1.39fF
C1434 a_46274_10496# a_47278_10496# 0.97fF
C1435 VDD a_18546_56172# 32.67fF
C1436 a_1586_33927# config_2_in[8] 0.34fF
C1437 VDD a_5497_62839# 1.90fF
C1438 VDD a_48282_12504# 0.52fF
C1439 VDD m2_24960_7214# 0.91fF
C1440 a_11149_40188# a_11389_40443# 0.71fF
C1441 a_22199_30287# a_27763_27221# 0.30fF
C1442 a_20170_65166# vcm 0.62fF
C1443 pmat.row_n[1] ctopn 1.65fF
C1444 a_27198_21540# vcm 0.65fF
C1445 a_3615_71631# a_11007_58229# 0.82fF
C1446 VDD a_25190_60146# 0.52fF
C1447 VDD a_1591_36501# 0.42fF
C1448 a_4985_51433# a_5785_48463# 0.46fF
C1449 a_42258_58138# vcm 0.62fF
C1450 a_45270_56130# m2_45040_54946# 0.99fF
C1451 VDD a_7563_63303# 0.48fF
C1452 a_18546_9490# ctopn 1.57fF
C1453 ANTENNA__1395__A1.DIODE pmat.col[3] 0.52fF
C1454 _1192_.A2 a_13459_28111# 1.24fF
C1455 a_3663_9269# a_4003_7663# 0.38fF
C1456 a_18546_19530# a_31122_19938# 0.35fF
C1457 a_21174_14512# ctopn 3.58fF
C1458 a_18546_12502# a_35138_12910# 0.35fF
C1459 a_26194_12504# a_27198_12504# 0.97fF
C1460 a_39246_22544# a_40250_22544# 0.97fF
C1461 VDD a_15383_44265# 0.64fF
C1462 VDD a_31214_16520# 0.52fF
C1463 VDD a_2676_51843# 0.62fF
C1464 pmat.rowon_n[8] cgen.dlycontrol1_in[0] 0.43fF
C1465 VDD a_21082_55126# 0.42fF
C1466 VDD a_41162_7890# 0.33fF
C1467 ANTENNA__1187__B1.DIODE ANTENNA__1196__A2.DIODE 17.85fF
C1468 ANTENNA__1395__A1.DIODE a_16800_47213# 0.58fF
C1469 a_34226_69182# vcm 0.62fF
C1470 VDD a_4396_69109# 0.82fF
C1471 a_30111_47911# a_13275_48783# 0.38fF
C1472 pmat.col_n[2] pmat.row_n[5] 0.45fF
C1473 a_18546_23546# a_40158_23954# 0.35fF
C1474 a_18547_51565# a_21371_50087# 0.54fF
C1475 a_1899_35051# a_6369_39465# 0.46fF
C1476 VDD a_37471_49551# 0.42fF
C1477 a_18546_9490# a_44174_9898# 0.35fF
C1478 a_19166_61150# ctopp 3.43fF
C1479 m2_51064_18258# m3_51196_18390# 2.76fF
C1480 a_43262_59142# vcm 0.62fF
C1481 _1224_.X _1519_.A 3.10fF
C1482 _1192_.A2 a_6829_26703# 0.43fF
C1483 a_1586_50247# a_5785_48463# 0.35fF
C1484 _1154_.X a_24867_53135# 0.42fF
C1485 a_10515_61839# a_10515_13967# 0.67fF
C1486 VDD a_38627_50613# 0.34fF
C1487 ANTENNA__1190__A1.DIODE a_21739_29415# 1.34fF
C1488 a_20170_56130# m2_18936_55950# 0.96fF
C1489 VDD a_1757_63701# 0.56fF
C1490 VDD a_13283_2767# 0.39fF
C1491 a_38242_56130# ctopp 3.40fF
C1492 a_19166_57134# a_20170_57134# 0.97fF
C1493 pmat.col[9] vcm 5.88fF
C1494 a_1586_18231# a_1591_18005# 0.71fF
C1495 VDD a_47278_56130# 0.55fF
C1496 _1194_.A2 a_35244_32411# 0.59fF
C1497 a_18975_40871# a_19409_40719# 0.89fF
C1498 a_10239_14183# a_7415_29397# 0.38fF
C1499 a_18546_71232# a_18162_71230# 2.62fF
C1500 VDD pmat.col[31] 6.57fF
C1501 a_34226_8488# m2_33996_7214# 1.00fF
C1502 a_20170_61150# vcm 0.62fF
C1503 VDD m3_18064_59094# 0.32fF
C1504 ANTENNA__1195__A1.DIODE a_40951_31599# 0.37fF
C1505 a_30210_21540# ctopn 3.58fF
C1506 pmat.col_n[11] pmat.col[12] 5.95fF
C1507 VDD a_29206_22544# 0.52fF
C1508 a_41254_66170# ctopp 3.58fF
C1509 VDD a_50290_66170# 0.54fF
C1510 nmat.col[21] ctopn 2.00fF
C1511 a_48282_11500# a_49286_11500# 0.97fF
C1512 VDD pmat.col_n[6] 5.50fF
C1513 a_34226_63158# ctopp 3.58fF
C1514 a_10883_3303# a_5351_19913# 0.46fF
C1515 VDD a_43262_63158# 0.52fF
C1516 a_26194_17524# vcm 0.65fF
C1517 a_50290_64162# a_50290_63158# 1.00fF
C1518 pmat.rowon_n[8] ctopn 0.60fF
C1519 m2_51064_57958# vcm 0.62fF
C1520 a_21371_50087# a_11948_49783# 1.37fF
C1521 a_18546_61192# a_42166_61150# 0.35fF
C1522 VDD a_11892_21959# 0.93fF
C1523 a_18162_68218# ctopp 1.49fF
C1524 VDD comp.adc_comp_circuit_0.adc_comp_buffer_0.in 0.57fF
C1525 m2_48052_54946# m2_49056_54946# 0.96fF
C1526 pmat.row_n[13] pmat.row_n[14] 3.46fF
C1527 a_27198_8488# vcm 0.64fF
C1528 a_50290_58138# a_50290_57134# 1.00fF
C1529 a_10515_15055# a_2835_13077# 0.94fF
C1530 a_10873_38517# a_12069_36341# 0.34fF
C1531 a_6927_30503# a_1781_9308# 1.16fF
C1532 a_2411_43301# a_2935_38279# 0.31fF
C1533 VDD a_7467_63303# 0.52fF
C1534 a_4075_50087# a_4399_51157# 0.93fF
C1535 a_43262_19532# vcm 0.65fF
C1536 a_42258_18528# a_42258_17524# 1.00fF
C1537 VDD a_37291_29397# 4.47fF
C1538 a_40951_31599# a_45829_35407# 0.90fF
C1539 a_11067_30287# a_19541_28879# 0.78fF
C1540 ANTENNA__1197__A.DIODE a_22199_30287# 0.67fF
C1541 a_42258_10496# vcm 0.65fF
C1542 a_18546_13506# a_36142_13914# 0.35fF
C1543 a_42258_63158# a_42258_62154# 1.00fF
C1544 a_39246_67174# ctopp 3.58fF
C1545 a_18546_18526# a_32126_18934# 0.35fF
C1546 _1196_.B1 ANTENNA__1184__B1.DIODE 2.29fF
C1547 a_12309_38659# cgen.dlycontrol1_in[4] 2.76fF
C1548 VDD a_48282_67174# 0.52fF
C1549 a_10441_21263# a_9075_28023# 0.35fF
C1550 a_48282_22544# a_48282_21540# 1.00fF
C1551 a_7457_62037# a_8193_61493# 0.62fF
C1552 a_22178_12504# vcm 0.65fF
C1553 a_27198_64162# ctopp 3.58fF
C1554 VDD a_37238_14512# 0.52fF
C1555 a_47278_14512# a_48282_14512# 0.97fF
C1556 VDD a_36234_64162# 0.52fF
C1557 nmat.en_bit_n[0] a_18563_27791# 0.36fF
C1558 a_44444_32233# a_35244_32411# 0.30fF
C1559 VDD a_24667_40719# 0.38fF
C1560 a_46274_64162# a_47278_64162# 0.97fF
C1561 VDD a_23821_35279# 3.03fF
C1562 a_18546_57176# a_50198_57134# 0.35fF
C1563 a_17139_30503# a_29937_31055# 2.12fF
C1564 VDD a_10703_50069# 0.57fF
C1565 a_41254_13508# a_41254_12504# 1.00fF
C1566 a_44266_23548# m2_44036_24282# 0.99fF
C1567 a_24591_28327# pmat.col[0] 0.78fF
C1568 VDD m3_20072_7346# 0.30fF
C1569 VDD config_1_in[14] 0.88fF
C1570 VDD a_13805_43990# 1.12fF
C1571 VDD m2_22952_24282# 0.62fF
C1572 a_14287_70543# pmat.rowon_n[11] 0.91fF
C1573 a_18243_28327# a_37820_30485# 0.48fF
C1574 a_3609_9295# a_3663_9269# 0.44fF
C1575 a_29206_17524# ctopn 3.58fF
C1576 a_44266_11500# vcm 0.65fF
C1577 VDD a_20170_62154# 0.52fF
C1578 a_2659_35015# cgen.dlycontrol4_in[2] 0.52fF
C1579 a_44966_43255# a_44733_44431# 0.51fF
C1580 VDD config_2_in[6] 0.71fF
C1581 a_30210_8488# ctopn 3.40fF
C1582 pmat.row_n[11] a_14839_66103# 0.64fF
C1583 a_18546_56172# a_33130_56130# 0.35fF
C1584 a_25190_56130# a_26194_56130# 0.97fF
C1585 pmat.row_n[15] a_13768_22325# 0.58fF
C1586 VDD a_32126_24958# 0.44fF
C1587 nmat.col_n[13] nmat.rowon_n[2] 3.99fF
C1588 m2_45040_24282# m2_46044_24282# 0.96fF
C1589 a_18162_7484# vcm 7.34fF
C1590 VDD a_9405_66627# 1.80fF
C1591 a_13643_29415# nmat.col_n[3] 1.53fF
C1592 a_46274_19532# ctopn 3.58fF
C1593 a_30210_65166# ctopp 3.58fF
C1594 ANTENNA__1196__A2.DIODE pmat.col[3] 0.35fF
C1595 a_10515_13967# a_6821_18543# 0.38fF
C1596 VDD a_39246_65166# 0.52fF
C1597 VDD a_46274_21540# 0.52fF
C1598 pmat.row_n[14] nmat.rowon_n[1] 20.34fF
C1599 a_48282_65166# a_48282_64162# 1.00fF
C1600 a_11041_39860# ndecision_finish 0.50fF
C1601 _1224_.X inp_analog 10.41fF
C1602 a_45270_10496# ctopn 3.58fF
C1603 a_15667_27239# a_17139_30503# 2.10fF
C1604 a_18546_68220# a_41162_68178# 0.35fF
C1605 VDD a_3052_29967# 0.47fF
C1606 a_48282_68178# vcm 0.62fF
C1607 pmat.row_n[7] ctopn 1.65fF
C1608 VDD a_2879_26703# 0.46fF
C1609 ANTENNA_fanout52_A.DIODE _1196_.B1 2.15fF
C1610 VDD a_6292_65479# 2.68fF
C1611 a_30210_62154# a_31214_62154# 0.97fF
C1612 a_37238_16520# a_37238_15516# 1.00fF
C1613 m2_51064_14242# m2_51064_13238# 0.99fF
C1614 a_28202_66170# a_29206_66170# 0.97fF
C1615 a_18546_60188# a_46182_60146# 0.35fF
C1616 a_25190_12504# ctopn 3.58fF
C1617 VDD a_44888_33205# 0.32fF
C1618 _1187_.A2 a_30663_50087# 0.40fF
C1619 a_21174_56130# vcm 0.62fF
C1620 a_18546_21538# a_20078_21946# 0.35fF
C1621 a_18162_21540# nmat.rowon_n[2] 1.33fF
C1622 _1194_.A2 nmat.col_n[31] 0.68fF
C1623 nmat.col_n[19] vcm 4.78fF
C1624 a_7415_29397# a_10147_29415# 0.51fF
C1625 nmat.rowon_n[14] a_2129_10383# 0.40fF
C1626 pmat.col[28] vcm 5.88fF
C1627 a_21174_63158# a_22178_63158# 0.97fF
C1628 a_18546_63200# a_25098_63158# 0.35fF
C1629 VDD m2_42028_72014# 1.00fF
C1630 a_5991_23983# a_9075_28023# 0.49fF
C1631 a_6283_31591# cgen.dlycontrol2_in[4] 0.81fF
C1632 a_44266_69182# ctopp 3.58fF
C1633 a_13091_28327# a_14943_26703# 0.40fF
C1634 a_24186_66170# vcm 0.62fF
C1635 a_14379_6567# a_13091_7655# 3.81fF
C1636 ANTENNA_fanout52_A.DIODE a_9785_28879# 0.50fF
C1637 m2_33996_72014# m2_35000_72014# 0.96fF
C1638 VDD a_34277_38550# 1.03fF
C1639 VDD conversion_finished_out 0.69fF
C1640 a_49286_65166# a_50290_65166# 0.97fF
C1641 a_26891_28327# a_29937_31055# 3.64fF
C1642 a_47278_11500# ctopn 3.58fF
C1643 a_11067_27239# nmat.col_n[29] 0.51fF
C1644 a_18162_71230# ctopp 1.30fF
C1645 pmat.rowoff_n[4] pmat.rowoff_n[6] 0.69fF
C1646 a_5363_33551# a_4075_31591# 3.38fF
C1647 pmat.rowon_n[7] a_10883_3303# 0.40fF
C1648 a_1769_47919# a_1739_47893# 0.40fF
C1649 a_11149_40188# cgen.dlycontrol4_in[1] 2.24fF
C1650 a_10781_42869# a_12237_38772# 0.84fF
C1651 VDD a_38793_49007# 0.32fF
C1652 a_11202_55687# a_13073_54997# 0.35fF
C1653 VDD a_3305_17999# 2.61fF
C1654 VDD a_10927_37981# 1.25fF
C1655 VDD nmat.en_bit_n[1] 11.98fF
C1656 a_30210_61150# ctopp 3.58fF
C1657 a_11067_64015# a_19541_28879# 1.15fF
C1658 a_29206_70186# a_30210_70186# 0.97fF
C1659 VDD a_12133_9001# 0.31fF
C1660 VDD a_39246_61150# 0.52fF
C1661 VDD a_39781_40157# 1.52fF
C1662 VDD a_19233_38215# 0.93fF
C1663 VDD a_27421_41814# 1.29fF
C1664 nmat.col_n[21] nmat.col_n[26] 0.67fF
C1665 nmat.col_n[28] nmat.col_n[24] 3.23fF
C1666 a_49286_18528# vcm 0.65fF
C1667 VDD a_33222_20536# 0.52fF
C1668 a_21174_10496# a_21174_9492# 1.00fF
C1669 a_18546_71232# a_30118_71190# 0.35fF
C1670 a_22178_67174# vcm 0.62fF
C1671 nmat.rowoff_n[6] a_18546_17522# 4.09fF
C1672 m3_19068_56082# ctopp 0.46fF
C1673 ANTENNA__1395__A1.DIODE a_18243_28327# 0.32fF
C1674 a_14641_57167# pmat.rowoff_n[4] 1.27fF
C1675 pmat.rowoff_n[12] a_10515_15055# 0.93fF
C1676 VDD m3_51196_55078# 0.30fF
C1677 a_12116_39783# a_22085_38550# 0.30fF
C1678 VDD a_45270_17524# 0.52fF
C1679 m2_18936_55950# ctopp 0.36fF
C1680 VDD a_4075_28335# 0.41fF
C1681 VDD a_31105_46805# 0.86fF
C1682 a_18546_8486# a_38150_8894# 0.35fF
C1683 pmat.row_n[3] a_18199_52789# 0.42fF
C1684 a_22178_60146# a_22178_59142# 1.00fF
C1685 a_18546_65208# a_35138_65166# 0.35fF
C1686 a_35230_55126# pmat.col[16] 0.38fF
C1687 VDD a_46274_8488# 0.55fF
C1688 a_11041_36596# a_12309_36483# 2.27fF
C1689 pmat.row_n[15] cgen.dlycontrol1_in[4] 0.69fF
C1690 a_18546_21538# a_49194_21946# 0.35fF
C1691 a_40250_62154# a_40250_61150# 1.00fF
C1692 VDD a_14125_13647# 0.34fF
C1693 ANTENNA__1183__B1.DIODE nmat.col[12] 0.36fF
C1694 VDD a_5357_62779# 0.69fF
C1695 a_13091_52047# a_12263_50959# 1.71fF
C1696 m2_50060_24282# m3_50192_24414# 0.85fF
C1697 a_18546_67216# a_35138_67174# 0.35fF
C1698 a_26194_67174# a_27198_67174# 0.97fF
C1699 a_5535_57993# a_5682_56311# 0.86fF
C1700 a_10223_26703# a_11091_26311# 0.68fF
C1701 a_23182_66170# a_23182_65166# 1.00fF
C1702 pmat.col_n[8] vcm 2.80fF
C1703 cgen.start_conv_in a_10873_36341# 0.89fF
C1704 VDD a_4253_42729# 0.32fF
C1705 VDD a_22178_15516# 0.52fF
C1706 a_40250_15516# a_40250_14512# 1.00fF
C1707 a_31152_48071# clk_ena 0.43fF
C1708 a_18546_7482# a_35138_7890# 0.35fF
C1709 _1184_.A2 a_15667_27239# 0.55fF
C1710 a_20170_68178# a_21174_68178# 0.97fF
C1711 a_42258_69182# a_42258_68178# 1.00fF
C1712 a_13091_18535# a_4383_7093# 0.68fF
C1713 a_50290_21540# a_50290_20536# 1.00fF
C1714 VDD a_5363_70543# 11.47fF
C1715 a_9411_2215# a_29937_31055# 1.06fF
C1716 VDD a_41254_12504# 0.52fF
C1717 cgen.dlycontrol4_in[2] a_24833_40719# 0.84fF
C1718 nmat.rowon_n[7] cgen.dlycontrol4_in[5] 2.55fF
C1719 VDD a_43315_48437# 0.97fF
C1720 a_19166_66170# a_20170_66170# 0.97fF
C1721 pmat.row_n[3] ctopp 1.65fF
C1722 a_10515_15055# nmat.sw 1.37fF
C1723 a_49286_57134# vcm 0.62fF
C1724 a_4075_50087# pmat.rowoff_n[12] 0.61fF
C1725 VDD a_33007_37683# 1.02fF
C1726 a_48282_71190# vcm 0.60fF
C1727 a_35230_58138# vcm 0.62fF
C1728 m2_42028_7214# m3_42160_7346# 2.79fF
C1729 a_30571_50959# _1183_.A2 0.31fF
C1730 a_18563_27791# a_6664_26159# 1.93fF
C1731 VDD a_5257_19087# 0.53fF
C1732 nmat.col_n[23] m2_42028_24282# 0.37fF
C1733 m2_17932_60970# vcm 0.44fF
C1734 nmat.col_n[26] nmat.col[26] 5.95fF
C1735 a_18546_19530# a_24094_19938# 0.35fF
C1736 a_28455_47381# a_28621_47381# 0.45fF
C1737 VDD a_3663_9269# 1.62fF
C1738 a_18546_12502# a_28110_12910# 0.35fF
C1739 a_5547_77295# a_5713_77295# 0.72fF
C1740 VDD a_24186_16520# 0.52fF
C1741 a_11497_40719# a_10927_41245# 0.46fF
C1742 VDD m2_46044_24282# 0.62fF
C1743 nmat.col[9] ctopn 1.97fF
C1744 a_6467_29415# clk_ena 0.61fF
C1745 VDD a_11235_26159# 0.84fF
C1746 VDD a_34134_7890# 0.33fF
C1747 pmat.col_n[5] pmat.col[6] 6.14fF
C1748 a_12309_36483# cgen.dlycontrol1_in[1] 1.93fF
C1749 a_19166_10496# a_20170_10496# 0.97fF
C1750 a_44266_11500# a_44266_10496# 1.00fF
C1751 VDD a_8477_57141# 0.60fF
C1752 ANTENNA__1395__A2.DIODE a_18243_28327# 1.71fF
C1753 a_11067_27239# a_13091_28327# 2.36fF
C1754 a_27198_69182# vcm 0.62fF
C1755 nmat.col_n[28] ctopn 2.03fF
C1756 nmat.col[30] nmat.col[18] 1.83fF
C1757 a_25190_23548# a_26194_23548# 0.97fF
C1758 a_18546_23546# a_33130_23954# 0.35fF
C1759 a_38851_28327# a_40837_46261# 0.83fF
C1760 pmat.sample pmat.row_n[6] 0.43fF
C1761 m2_27972_24282# vcm 0.42fF
C1762 cgen.dlycontrol3_in[2] a_2411_33749# 0.44fF
C1763 pmat.rowon_n[0] a_10497_54697# 0.34fF
C1764 a_27198_9492# a_28202_9492# 0.97fF
C1765 a_18546_9490# a_37146_9898# 0.35fF
C1766 a_49286_61150# a_50290_61150# 0.97fF
C1767 nmat.col_n[16] vcm 2.79fF
C1768 VDD a_8891_66964# 1.00fF
C1769 a_36234_59142# vcm 0.62fF
C1770 a_34226_12504# a_34226_11500# 1.00fF
C1771 VDD a_24197_42405# 1.26fF
C1772 a_18546_24550# a_20078_24958# 0.39fF
C1773 VDD a_3688_17179# 2.52fF
C1774 nmat.rowon_n[13] nmat.rowoff_n[10] 0.52fF
C1775 a_5682_56311# a_6559_33767# 0.34fF
C1776 a_31214_56130# ctopp 3.40fF
C1777 VDD a_30603_29575# 0.60fF
C1778 a_4831_34561# a_4792_34435# 0.42fF
C1779 VDD a_40250_56130# 0.55fF
C1780 a_43262_20536# a_44266_20536# 0.97fF
C1781 a_6283_31591# a_6830_44655# 0.38fF
C1782 pmat.row_n[15] nmat.col[7] 0.60fF
C1783 VDD a_7072_26311# 0.46fF
C1784 VDD m3_48184_72146# 0.32fF
C1785 a_23182_21540# ctopn 3.58fF
C1786 _1224_.X ANTENNA__1395__B1.DIODE 4.70fF
C1787 ANTENNA__1190__A1.DIODE a_24867_53135# 0.99fF
C1788 a_18546_66212# a_50198_66170# 0.35fF
C1789 a_42258_9492# a_42258_8488# 1.00fF
C1790 a_2263_43719# a_1957_43567# 0.76fF
C1791 pmat.col_n[31] ANTENNA__1395__A2.DIODE 0.30fF
C1792 VDD a_22178_22544# 0.52fF
C1793 a_34226_66170# ctopp 3.58fF
C1794 a_25695_28111# nmat.col[18] 0.61fF
C1795 m2_33996_72014# m3_34128_72146# 2.79fF
C1796 a_10515_61839# a_13091_7655# 1.45fF
C1797 a_25879_31591# nmat.col_n[12] 0.46fF
C1798 VDD a_43262_66170# 0.52fF
C1799 a_24186_21540# a_25190_21540# 0.97fF
C1800 VDD a_18162_72234# 29.28fF
C1801 a_27198_63158# ctopp 3.58fF
C1802 VDD a_19584_52423# 4.22fF
C1803 VDD a_36234_63158# 0.52fF
C1804 a_35230_62154# pmat.col[16] 0.31fF
C1805 a_18546_61192# a_35138_61150# 0.35fF
C1806 VDD a_2191_24501# 0.37fF
C1807 nmat.sw cgen.dlycontrol4_in[3] 0.35fF
C1808 m2_41024_54946# m2_42028_54946# 0.96fF
C1809 a_25190_71190# a_25190_70186# 1.00fF
C1810 nmat.col[24] nmat.col_n[25] 0.42fF
C1811 a_39246_58138# a_40250_58138# 0.97fF
C1812 VDD a_6541_15279# 0.61fF
C1813 VDD nmat.col[8] 4.83fF
C1814 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[28] 0.60fF
C1815 VDD a_14691_29575# 0.91fF
C1816 ANTENNA__1190__B1.DIODE a_26479_32117# 0.39fF
C1817 a_36234_19532# vcm 0.65fF
C1818 a_18243_28327# ANTENNA__1196__A2.DIODE 0.80fF
C1819 pmat.row_n[1] ctopp 1.64fF
C1820 a_1923_61759# a_1591_65327# 0.51fF
C1821 a_2046_30184# a_5823_34863# 0.34fF
C1822 a_17139_30503# a_44870_48437# 0.36fF
C1823 m2_17932_60970# m2_17932_59966# 0.99fF
C1824 a_14887_46377# a_33839_46805# 0.35fF
C1825 a_18546_16518# ctopn 1.59fF
C1826 a_11067_27239# a_17139_30503# 0.38fF
C1827 ANTENNA__1395__A1.DIODE a_30571_50959# 0.50fF
C1828 a_35230_10496# vcm 0.65fF
C1829 a_23182_13508# a_24186_13508# 0.97fF
C1830 a_18546_13506# a_29114_13914# 0.35fF
C1831 _1194_.B1 a_13643_29415# 0.70fF
C1832 pmat.row_n[5] a_18546_13506# 0.35fF
C1833 nmat.col_n[20] ctopn 2.02fF
C1834 VDD m2_51064_62978# 1.03fF
C1835 VDD a_38695_48634# 0.40fF
C1836 a_11041_38772# a_11113_36483# 0.36fF
C1837 a_2407_49289# a_5065_63669# 0.57fF
C1838 a_39246_61150# a_39246_60146# 1.00fF
C1839 VDD a_45866_38279# 0.63fF
C1840 a_32218_67174# ctopp 3.58fF
C1841 a_18546_18526# a_25098_18934# 0.35fF
C1842 a_21174_18528# a_22178_18528# 0.97fF
C1843 a_47278_19532# a_47278_18528# 1.00fF
C1844 VDD a_41254_67174# 0.52fF
C1845 VDD a_10985_37692# 1.19fF
C1846 a_20170_64162# ctopp 3.57fF
C1847 VDD a_30210_14512# 0.52fF
C1848 a_28202_56130# m2_27972_54946# 0.99fF
C1849 VDD a_29206_64162# 0.52fF
C1850 a_17842_27497# nmat.col_n[21] 0.77fF
C1851 a_18546_17522# a_47186_17930# 0.35fF
C1852 nmat.rowon_n[12] ANTENNA__1190__A2.DIODE 0.72fF
C1853 a_18546_57176# a_43170_57134# 0.35fF
C1854 _1183_.A2 nmat.col_n[1] 0.31fF
C1855 a_40250_59142# a_40250_58138# 1.00fF
C1856 nmat.col_n[31] a_50290_23548# 0.33fF
C1857 a_1923_69823# a_1899_35051# 0.53fF
C1858 a_19166_9492# vcm 0.65fF
C1859 VDD a_8456_69135# 0.47fF
C1860 VDD a_6651_44661# 0.37fF
C1861 VDD a_46863_28585# 0.41fF
C1862 a_32218_15516# a_33222_15516# 0.97fF
C1863 a_18546_15514# a_47186_15922# 0.35fF
C1864 VDD m2_42028_54946# 0.62fF
C1865 a_5179_31591# a_2007_25597# 0.77fF
C1866 VDD a_11071_46805# 0.52fF
C1867 _1192_.A2 a_32405_32463# 1.83fF
C1868 a_8243_7290# a_7939_7125# 0.31fF
C1869 pmat.row_n[4] pmat.rowon_n[0] 4.61fF
C1870 a_31214_69182# a_32218_69182# 0.97fF
C1871 pmat.col_n[16] ctopp 2.04fF
C1872 cgen.dlycontrol1_in[4] a_29404_36165# 0.33fF
C1873 VDD a_29367_35831# 0.63fF
C1874 a_50290_70186# vcm 0.62fF
C1875 a_22178_17524# ctopn 3.58fF
C1876 VDD a_42166_72194# 0.32fF
C1877 a_37238_11500# vcm 0.65fF
C1878 pmat.col[19] ctopp 1.97fF
C1879 VDD a_7457_62037# 1.24fF
C1880 a_45270_17524# a_45270_16520# 1.00fF
C1881 m2_23956_54946# vcm 0.42fF
C1882 m2_51064_23278# m3_51196_23410# 2.76fF
C1883 a_23182_8488# ctopn 3.40fF
C1884 ANTENNA__1197__A.DIODE a_18563_27791# 0.78fF
C1885 a_18546_56172# a_26102_56130# 0.35fF
C1886 VDD a_25098_24958# 0.44fF
C1887 ANTENNA__1190__A1.DIODE a_38851_28327# 0.45fF
C1888 _1187_.A2 a_10883_3303# 0.40fF
C1889 m2_38012_24282# m2_39016_24282# 0.96fF
C1890 pmat.rowoff_n[6] vcm 0.32fF
C1891 pmat.rowon_n[7] a_7717_14735# 0.55fF
C1892 a_7109_29423# a_26479_32117# 4.23fF
C1893 a_39246_19532# ctopn 3.58fF
C1894 a_23182_65166# ctopp 3.58fF
C1895 VDD a_32035_43177# 0.66fF
C1896 a_29217_41570# a_30523_41245# 0.62fF
C1897 VDD a_32218_65166# 0.52fF
C1898 a_9963_28111# a_13479_26935# 0.74fF
C1899 ANTENNA__1190__B1.DIODE nmat.rowon_n[5] 0.45fF
C1900 VDD a_39246_21540# 0.52fF
C1901 a_40250_59142# a_41254_59142# 0.97fF
C1902 _1184_.A2 a_10423_16055# 0.39fF
C1903 a_38242_10496# ctopn 3.58fF
C1904 a_18546_68220# a_34134_68178# 0.35fF
C1905 a_45270_58138# ctopp 3.58fF
C1906 a_41254_68178# vcm 0.62fF
C1907 a_1899_35051# a_1586_63927# 1.93fF
C1908 a_29206_23548# a_29206_22544# 1.00fF
C1909 a_6283_31591# a_22199_32149# 0.40fF
C1910 nmat.sw a_5899_21807# 0.42fF
C1911 a_28525_43655# a_28981_43493# 0.31fF
C1912 a_5654_9527# a_5935_6575# 0.34fF
C1913 a_28202_60146# a_29206_60146# 0.97fF
C1914 a_18546_60188# a_39154_60146# 0.35fF
C1915 pmat.rowon_n[8] ctopp 1.57fF
C1916 a_22199_30287# nmat.col[19] 0.58fF
C1917 a_2419_53351# a_1586_63927# 0.43fF
C1918 VDD a_46130_34319# 1.33fF
C1919 a_11067_27239# a_26891_28327# 0.34fF
C1920 a_11067_49871# a_13643_29415# 0.93fF
C1921 pmat.rowoff_n[7] a_10239_14183# 1.05fF
C1922 VDD m2_27972_72014# 1.13fF
C1923 a_36234_68178# a_36234_67174# 1.00fF
C1924 a_46274_23548# vcm 0.65fF
C1925 a_37238_69182# ctopp 3.58fF
C1926 a_48282_9492# vcm 0.65fF
C1927 VDD a_46274_69182# 0.52fF
C1928 a_4259_31375# a_10883_3303# 3.19fF
C1929 m2_26968_72014# m2_27972_72014# 0.96fF
C1930 a_1591_65327# a_2944_65576# 0.34fF
C1931 VDD a_18272_39429# 1.14fF
C1932 VDD a_7907_52031# 0.45fF
C1933 a_46274_59142# ctopp 3.58fF
C1934 a_40250_11500# ctopn 3.58fF
C1935 VDD a_7047_31226# 0.51fF
C1936 a_11067_27239# _1184_.A2 0.76fF
C1937 a_21279_48999# a_38557_48469# 0.60fF
C1938 VDD a_1959_12791# 0.79fF
C1939 a_2199_13887# a_2327_11477# 0.45fF
C1940 a_11149_40188# a_10873_39605# 0.34fF
C1941 a_34226_16520# a_35230_16520# 0.97fF
C1942 a_6679_15492# a_6541_15279# 0.56fF
C1943 a_18546_16518# a_51202_16926# 0.35fF
C1944 a_4523_21276# a_3305_17999# 0.42fF
C1945 m2_51064_20266# m3_51196_20398# 2.76fF
C1946 pmat.col[20] vcm 5.88fF
C1947 a_24186_67174# a_24186_66170# 1.00fF
C1948 VDD a_3859_23699# 0.48fF
C1949 a_23182_61150# ctopp 3.58fF
C1950 nmat.col[7] nmat.col_n[6] 6.77fF
C1951 VDD a_32218_61150# 0.52fF
C1952 a_13597_37571# a_14719_37737# 0.48fF
C1953 a_15049_42902# a_11297_36091# 1.01fF
C1954 a_44266_13508# vcm 0.65fF
C1955 VDD a_15420_41831# 1.08fF
C1956 VDD a_2129_12559# 1.24fF
C1957 VDD a_6639_63927# 0.57fF
C1958 a_31339_31787# a_25575_31055# 0.40fF
C1959 a_42258_18528# vcm 0.65fF
C1960 VDD a_26194_20536# 0.52fF
C1961 a_23182_17524# a_24186_17524# 0.97fF
C1962 a_21174_57134# a_22178_57134# 0.97fF
C1963 a_26194_20536# a_26194_19532# 1.00fF
C1964 a_18546_71232# a_23090_71190# 0.35fF
C1965 a_20170_71190# a_21174_71190# 0.97fF
C1966 a_27198_23548# m2_26968_24282# 0.99fF
C1967 a_12513_39100# a_14773_38306# 1.06fF
C1968 VDD a_38242_17524# 0.52fF
C1969 a_10949_43124# a_16355_43123# 0.73fF
C1970 nmat.en_bit_n[1] a_8583_29199# 0.58fF
C1971 a_31675_47695# a_35244_32411# 2.18fF
C1972 _1196_.B1 a_17139_30503# 0.59fF
C1973 a_24186_8488# a_25190_8488# 0.97fF
C1974 a_18546_8486# a_31122_8894# 0.35fF
C1975 a_18546_65208# a_28110_65166# 0.35fF
C1976 a_43262_70186# a_43262_69182# 1.00fF
C1977 VDD a_39246_8488# 0.55fF
C1978 VDD a_9963_13967# 11.16fF
C1979 a_18546_21538# a_42166_21946# 0.35fF
C1980 VDD pmat.col_n[9] 5.66fF
C1981 a_11067_27239# a_9411_2215# 1.47fF
C1982 a_32218_14512# a_32218_13508# 1.00fF
C1983 a_14653_53458# a_12263_50959# 0.40fF
C1984 a_49286_23548# ctopn 3.39fF
C1985 cgen.dlycontrol4_in[4] a_13805_43990# 0.73fF
C1986 pmat.row_n[9] a_18162_17524# 25.57fF
C1987 a_18546_67216# a_28110_67174# 0.35fF
C1988 a_36234_57134# a_36234_56130# 1.00fF
C1989 pmat.rowon_n[0] a_18162_56170# 1.19fF
C1990 a_12447_16143# a_13091_52047# 0.53fF
C1991 VDD a_9063_24527# 0.31fF
C1992 ANTENNA__1184__B1.DIODE a_22199_30287# 2.15fF
C1993 a_5363_70543# a_10595_53361# 0.61fF
C1994 a_40250_19532# a_41254_19532# 0.97fF
C1995 a_49286_60146# vcm 0.62fF
C1996 nmat.col_n[30] nmat.col[19] 6.23fF
C1997 pmat.rowon_n[0] a_3305_27791# 1.40fF
C1998 nmat.col_n[5] ctopn 2.02fF
C1999 a_7109_29423# a_5179_31591# 0.51fF
C2000 pmat.row_n[7] ctopp 1.65fF
C2001 VDD a_40349_40726# 1.85fF
C2002 a_2199_13887# a_4241_13653# 0.63fF
C2003 pmat.col_n[29] m2_48052_54946# 0.43fF
C2004 pmat.col_n[17] pmat.col[18] 6.11fF
C2005 a_18546_7482# a_28110_7890# 0.35fF
C2006 a_5363_33551# a_14917_23983# 0.47fF
C2007 a_13459_28111# a_16311_28327# 1.84fF
C2008 pmat.rowon_n[0] nmat.rowon_n[15] 20.52fF
C2009 a_30571_50959# a_41926_46983# 0.40fF
C2010 a_20170_10496# ctopn 3.57fF
C2011 a_2419_69455# a_1586_63927# 0.30fF
C2012 a_39246_10496# a_40250_10496# 0.97fF
C2013 _1194_.A2 _1183_.A2 0.64fF
C2014 VDD a_34226_12504# 0.52fF
C2015 pmat.col[9] m2_27972_54946# 0.40fF
C2016 VDD pmat.sample 8.53fF
C2017 VDD a_3951_77055# 0.40fF
C2018 cgen.dlycontrol3_in[1] cgen.dlycontrol2_in[3] 1.80fF
C2019 a_19166_60146# a_20170_60146# 0.97fF
C2020 a_47278_13508# ctopn 3.58fF
C2021 VDD a_1644_59861# 0.33fF
C2022 a_42258_57134# vcm 0.62fF
C2023 VDD a_15651_37737# 0.59fF
C2024 a_2411_16101# a_2467_18517# 0.58fF
C2025 a_41254_71190# vcm 0.60fF
C2026 a_12116_40871# a_11297_36091# 0.58fF
C2027 pmat.rowon_n[7] pmat.row_n[1] 0.46fF
C2028 a_45270_18528# ctopn 3.58fF
C2029 a_17842_27497# nmat.col_n[10] 0.35fF
C2030 a_28202_58138# vcm 0.62fF
C2031 ANTENNA__1395__A2.DIODE nmat.col_n[1] 0.54fF
C2032 VDD a_31925_40955# 1.59fF
C2033 clk_vcm nmat.col[29] 1.00fF
C2034 VDD a_46523_39733# 0.94fF
C2035 a_1858_25615# a_19439_30511# 0.33fF
C2036 a_19166_69182# ctopp 3.43fF
C2037 pmat.col[21] ctopp 1.97fF
C2038 ANTENNA__1190__A1.DIODE nmat.col_n[19] 0.37fF
C2039 pmat.rowoff_n[7] ctopn 1.40fF
C2040 a_7717_14735# nmat.col[29] 1.07fF
C2041 a_50290_63158# pmat.col[31] 0.31fF
C2042 cgen.dlycontrol4_in[1] a_2467_35925# 0.51fF
C2043 VDD m3_35132_7346# 0.37fF
C2044 a_32218_22544# a_33222_22544# 0.97fF
C2045 VDD a_23700_44869# 1.00fF
C2046 ANTENNA__1187__B1.DIODE nmat.col_n[21] 0.38fF
C2047 _1196_.B1 a_11927_27399# 0.61fF
C2048 nmat.rowon_n[7] nmat.col_n[10] 1.20fF
C2049 a_14287_69455# pmat.rowoff_n[12] 0.33fF
C2050 VDD a_30527_31573# 0.33fF
C2051 VDD a_27106_7890# 0.34fF
C2052 a_14773_37218# a_11921_35286# 0.52fF
C2053 a_20170_69182# vcm 0.62fF
C2054 a_5363_70543# a_10167_64239# 0.38fF
C2055 a_18546_23546# a_26102_23954# 0.35fF
C2056 a_10515_13967# a_9411_2215# 1.08fF
C2057 a_46274_63158# a_47278_63158# 0.97fF
C2058 m2_47048_54946# vcm 0.42fF
C2059 VDD m2_17932_65990# 1.00fF
C2060 a_18546_9490# a_30118_9898# 0.35fF
C2061 VDD a_35230_24552# 0.58fF
C2062 VDD a_4396_66933# 0.44fF
C2063 a_29206_59142# vcm 0.62fF
C2064 VDD a_4081_61127# 0.85fF
C2065 a_37820_30485# a_44444_32233# 0.39fF
C2066 a_8472_11739# a_8479_11484# 0.62fF
C2067 pmat.row_n[15] a_4068_25615# 0.74fF
C2068 a_50290_16520# m2_51064_16250# 0.96fF
C2069 a_24186_56130# ctopp 3.40fF
C2070 VDD a_7939_29967# 0.58fF
C2071 VDD a_33222_56130# 0.55fF
C2072 a_11067_27239# nmat.col[13] 1.62fF
C2073 a_24591_28327# nmat.col_n[18] 0.96fF
C2074 a_30663_50087# a_25695_28111# 1.35fF
C2075 a_1717_13647# a_8511_10422# 0.30fF
C2076 VDD m3_20072_72146# 0.34fF
C2077 VDD a_20170_17524# 0.52fF
C2078 VDD a_38575_50639# 0.31fF
C2079 a_18546_62196# a_47186_62154# 0.35fF
C2080 _1196_.B1 _1184_.A2 12.42fF
C2081 VDD a_43267_47081# 0.40fF
C2082 a_18546_66212# a_43170_66170# 0.35fF
C2083 a_9135_60967# a_12447_16143# 3.83fF
C2084 a_27198_66170# ctopp 3.58fF
C2085 a_11711_50959# nmat.col[15] 0.50fF
C2086 VDD a_36234_66170# 0.52fF
C2087 pmat.row_n[15] nmat.col[3] 0.39fF
C2088 a_11317_36924# a_11113_36483# 0.32fF
C2089 a_41254_11500# a_42258_11500# 0.97fF
C2090 VDD a_30155_36893# 1.52fF
C2091 ANTENNA__1196__A2.DIODE nmat.col_n[1] 1.34fF
C2092 a_25743_49783# a_25839_49783# 0.32fF
C2093 a_20170_63158# ctopp 3.57fF
C2094 a_21739_29415# a_23021_29199# 0.34fF
C2095 nmat.col[27] vcm 5.76fF
C2096 pmat.row_n[14] pmat.row_n[8] 2.37fF
C2097 VDD a_29206_63158# 0.52fF
C2098 a_11435_58791# a_6467_29415# 5.83fF
C2099 a_43262_64162# a_43262_63158# 1.00fF
C2100 a_11067_64015# a_10239_14183# 3.17fF
C2101 _1224_.X _1192_.B1 4.71fF
C2102 ANTENNA__1197__A.DIODE a_16113_52271# 0.47fF
C2103 _1194_.A2 ANTENNA__1395__A1.DIODE 1.03fF
C2104 a_46274_10496# a_46274_9492# 1.00fF
C2105 a_18546_61192# a_28110_61150# 0.35fF
C2106 a_43262_58138# a_43262_57134# 1.00fF
C2107 _1184_.A2 a_9785_28879# 0.57fF
C2108 pmat.rowoff_n[15] pmat.row_n[14] 1.75fF
C2109 a_6451_67655# a_14287_70543# 0.58fF
C2110 pmat.rowon_n[8] pmat.rowon_n[7] 0.99fF
C2111 pmat.rowon_n[11] nmat.rowon_n[7] 0.53fF
C2112 a_19584_52423# a_22499_49783# 0.34fF
C2113 a_29937_31055# a_37637_32149# 0.54fF
C2114 VDD a_2847_43327# 0.35fF
C2115 pmat.sample_n pmat.sample 9.18fF
C2116 VDD a_18823_50247# 6.01fF
C2117 a_29206_19532# vcm 0.65fF
C2118 a_47278_60146# a_47278_59142# 1.00fF
C2119 a_35230_18528# a_35230_17524# 1.00fF
C2120 VDD a_35138_55126# 0.38fF
C2121 VDD a_5528_57685# 0.38fF
C2122 a_4075_50087# a_1586_63927# 0.41fF
C2123 VDD a_1923_31743# 9.36fF
C2124 a_4075_50087# a_1769_47919# 0.63fF
C2125 a_37820_30485# a_32687_46607# 0.36fF
C2126 a_28202_10496# vcm 0.65fF
C2127 a_18546_13506# a_22086_13914# 0.35fF
C2128 a_3305_17999# a_3305_15823# 1.11fF
C2129 a_11337_25071# nmat.col_n[1] 0.63fF
C2130 nmat.col[18] comp_latch 0.60fF
C2131 a_35230_63158# a_35230_62154# 1.00fF
C2132 a_30210_71190# m2_29980_72014# 1.00fF
C2133 VDD a_7578_48553# 0.50fF
C2134 _1183_.A2 a_32687_46607# 0.73fF
C2135 _1196_.B1 a_9411_2215# 2.52fF
C2136 VDD a_18546_23546# 32.78fF
C2137 a_25190_67174# ctopp 3.58fF
C2138 a_19166_63158# m2_17932_62978# 0.96fF
C2139 a_18546_70228# a_45178_70186# 0.35fF
C2140 VDD a_34226_67174# 0.52fF
C2141 a_14491_51969# a_14452_51843# 0.72fF
C2142 a_13432_62581# a_12003_52815# 0.36fF
C2143 VDD a_26515_38007# 0.59fF
C2144 a_41254_22544# a_41254_21540# 1.00fF
C2145 a_48282_66170# a_48282_65166# 1.00fF
C2146 VDD a_23182_14512# 0.52fF
C2147 a_40250_14512# a_41254_14512# 0.97fF
C2148 a_44266_62154# vcm 0.62fF
C2149 m2_51064_12234# vcm 0.51fF
C2150 VDD a_22178_64162# 0.52fF
C2151 pmat.sample a_21032_44007# 0.31fF
C2152 VDD a_4831_40303# 0.40fF
C2153 a_39246_64162# a_40250_64162# 0.97fF
C2154 a_18546_17522# a_40158_17930# 0.35fF
C2155 a_45270_68178# a_46274_68178# 0.97fF
C2156 a_18546_57176# a_36142_57134# 0.35fF
C2157 nmat.sw nmat.col_n[29] 0.51fF
C2158 a_34226_13508# a_34226_12504# 1.00fF
C2159 a_5687_71829# a_5081_53135# 2.65fF
C2160 a_6283_31591# nmat.col_n[12] 0.86fF
C2161 a_10949_43124# a_10781_42364# 1.48fF
C2162 pmat.col_n[6] pmat.col[7] 6.01fF
C2163 a_18546_15514# a_40158_15922# 0.35fF
C2164 a_9983_32385# a_9944_32259# 0.42fF
C2165 VDD a_34243_32143# 0.51fF
C2166 _1196_.B1 a_7939_31591# 0.32fF
C2167 VDD a_15144_36165# 1.08fF
C2168 a_43262_70186# vcm 0.62fF
C2169 a_30210_11500# vcm 0.65fF
C2170 a_12461_29673# a_8443_20719# 0.34fF
C2171 pmat.row_n[4] a_17397_48463# 0.33fF
C2172 nmat.sw a_11149_40188# 0.42fF
C2173 pmat.col_n[11] vcm 2.80fF
C2174 a_10873_39605# a_11681_35823# 0.81fF
C2175 a_6283_31591# a_35559_30209# 0.37fF
C2176 a_32218_19532# ctopn 3.58fF
C2177 VDD a_13719_43177# 0.57fF
C2178 VDD a_25190_65166# 0.52fF
C2179 a_10055_31591# a_2411_33749# 0.80fF
C2180 VDD a_4516_21531# 6.43fF
C2181 ANTENNA__1190__B1.DIODE a_28704_29568# 1.06fF
C2182 VDD a_32218_21540# 0.52fF
C2183 _1194_.A2 ANTENNA__1395__A2.DIODE 6.12fF
C2184 ANTENNA__1197__A.DIODE _1194_.B1 0.32fF
C2185 a_41254_65166# a_41254_64162# 1.00fF
C2186 a_31214_10496# ctopn 3.58fF
C2187 a_18546_68220# a_27106_68178# 0.35fF
C2188 VDD a_41227_29423# 1.87fF
C2189 a_2149_45717# a_4259_73807# 0.72fF
C2190 a_38242_58138# ctopp 3.58fF
C2191 a_34226_68178# vcm 0.62fF
C2192 VDD a_1643_69653# 0.37fF
C2193 VDD a_47278_58138# 0.52fF
C2194 cgen.dlycontrol3_in[0] a_11565_39061# 0.45fF
C2195 a_13655_26703# nmat.col_n[1] 0.66fF
C2196 VDD a_1757_27797# 0.62fF
C2197 nmat.rowon_n[14] ctopn 1.40fF
C2198 a_3746_58487# a_8907_48437# 0.31fF
C2199 a_30210_16520# a_30210_15516# 1.00fF
C2200 a_23182_62154# a_24186_62154# 0.97fF
C2201 a_49286_71190# m2_49056_72014# 1.00fF
C2202 VDD a_2935_38279# 3.43fF
C2203 a_21174_66170# a_22178_66170# 0.97fF
C2204 a_18546_60188# a_32126_60146# 0.35fF
C2205 pmat.rowon_n[7] pmat.row_n[7] 22.00fF
C2206 nmat.sw a_11921_41814# 0.37fF
C2207 VDD a_18546_66212# 32.63fF
C2208 a_17139_30503# a_45019_38645# 0.32fF
C2209 VDD a_35244_32411# 9.15fF
C2210 pmat.rowon_n[10] pmat.rowoff_n[10] 20.76fF
C2211 a_10873_38517# clk_ena 1.49fF
C2212 m2_47048_7214# m3_47180_7346# 2.79fF
C2213 VDD a_51202_64162# 0.30fF
C2214 VDD nmat.rowon_n[4] 4.01fF
C2215 a_10515_15055# pmat.rowoff_n[4] 2.32fF
C2216 nmat.col_n[24] m2_43032_24282# 0.37fF
C2217 m2_24960_54946# m3_25092_55078# 2.79fF
C2218 pmat.sample_n a_18823_50247# 0.68fF
C2219 a_39246_23548# vcm 0.65fF
C2220 a_9583_10121# a_12257_8527# 0.49fF
C2221 a_30210_69182# ctopp 3.58fF
C2222 a_41254_9492# vcm 0.65fF
C2223 VDD a_39246_69182# 0.52fF
C2224 ANTENNA__1187__B1.DIODE nmat.col_n[10] 0.34fF
C2225 m2_19940_72014# m2_20944_72014# 0.96fF
C2226 a_19233_41479# a_19689_41317# 0.32fF
C2227 a_2007_25597# a_29163_29423# 0.53fF
C2228 a_42258_65166# a_43262_65166# 0.97fF
C2229 a_39246_59142# ctopp 3.58fF
C2230 pmat.rowoff_n[4] a_14379_6567# 0.75fF
C2231 a_33222_11500# ctopn 3.58fF
C2232 a_10515_15055# nmat.col_n[3] 1.89fF
C2233 VDD a_48282_59142# 0.52fF
C2234 a_49286_21540# a_50290_21540# 0.97fF
C2235 _1184_.A2 a_2835_13077# 0.43fF
C2236 a_3866_57399# a_4265_71543# 0.90fF
C2237 a_22199_30287# nmat.col_n[29] 0.75fF
C2238 a_19166_16520# vcm 0.65fF
C2239 a_15667_27239# a_25879_31591# 1.05fF
C2240 a_18546_16518# a_44174_16926# 0.35fF
C2241 m2_37008_24282# vcm 0.42fF
C2242 a_6787_47607# a_10055_31591# 0.82fF
C2243 comp.adc_comp_circuit_0.adc_comp_buffer_1.in a_53622_39932# 0.44fF
C2244 a_22178_70186# a_23182_70186# 0.97fF
C2245 nmat.col[28] nmat.col[18] 3.57fF
C2246 a_50290_71190# a_50290_70186# 1.00fF
C2247 VDD a_13432_62581# 3.98fF
C2248 VDD a_25190_61150# 0.52fF
C2249 a_14773_38306# a_24015_36911# 0.38fF
C2250 a_3305_15823# a_3688_17179# 1.10fF
C2251 VDD a_28131_50069# 3.80fF
C2252 a_37238_13508# vcm 0.65fF
C2253 VDD a_27947_41245# 1.27fF
C2254 a_2007_25597# a_1586_18231# 0.85fF
C2255 a_13091_52047# a_13459_28111# 1.55fF
C2256 _1194_.A2 ANTENNA__1196__A2.DIODE 6.62fF
C2257 a_35230_18528# vcm 0.65fF
C2258 VDD a_18162_20536# 2.74fF
C2259 ANTENNA__1195__A1.DIODE nmat.col[29] 0.47fF
C2260 ANTENNA__1197__B.DIODE a_21371_50087# 0.83fF
C2261 a_9545_66567# a_10499_67503# 0.34fF
C2262 VDD a_35520_30083# 0.30fF
C2263 a_44382_40847# a_44444_32233# 0.53fF
C2264 VDD a_9827_53379# 0.63fF
C2265 a_48282_13508# a_49286_13508# 0.97fF
C2266 cgen.enable_dlycontrol_in a_11057_35836# 0.52fF
C2267 a_46274_15516# vcm 0.65fF
C2268 VDD a_31214_17524# 0.52fF
C2269 VDD vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 44.59fF
C2270 a_2215_47375# cgen.enable_dlycontrol_in 0.56fF
C2271 a_18546_8486# a_24094_8894# 0.35fF
C2272 a_18546_65208# a_21082_65166# 0.35fF
C2273 m2_39016_72014# m3_39148_72146# 2.79fF
C2274 a_46274_18528# a_47278_18528# 0.97fF
C2275 nmat.rowon_n[7] a_2389_45859# 1.04fF
C2276 VDD a_32218_8488# 0.55fF
C2277 a_13091_52047# a_12044_49641# 0.34fF
C2278 a_8443_20719# a_9741_28585# 0.38fF
C2279 a_18546_21538# a_35138_21946# 0.35fF
C2280 _1154_.X clk_comp 1.04fF
C2281 nmat.rowon_n[7] a_12447_16143# 1.07fF
C2282 a_33222_62154# a_33222_61150# 1.00fF
C2283 a_42258_23548# ctopn 3.40fF
C2284 VDD a_48282_19532# 0.52fF
C2285 a_44266_9492# ctopn 3.57fF
C2286 a_18546_67216# a_21082_67174# 0.35fF
C2287 a_7847_56085# a_8013_56085# 0.75fF
C2288 VDD a_3325_23439# 0.64fF
C2289 a_42258_60146# vcm 0.62fF
C2290 VDD a_47278_10496# 0.52fF
C2291 VDD a_11497_40719# 6.01fF
C2292 a_12116_40871# a_11921_41814# 0.97fF
C2293 a_11041_40948# a_14149_39747# 0.52fF
C2294 a_4383_7093# a_9583_10121# 0.41fF
C2295 a_33222_15516# a_33222_14512# 1.00fF
C2296 pmat.col_n[25] m2_44036_54946# 0.32fF
C2297 a_3615_71631# a_12263_50959# 0.32fF
C2298 VDD a_36453_29199# 1.14fF
C2299 a_36234_55126# ctopp 0.65fF
C2300 a_16800_47213# a_12263_50959# 0.68fF
C2301 a_46274_63158# pmat.col[27] 0.31fF
C2302 a_35230_69182# a_35230_68178# 1.00fF
C2303 VDD a_28803_31055# 0.76fF
C2304 a_34226_24552# m3_34128_24414# 2.08fF
C2305 a_19166_19532# m2_17932_19262# 0.96fF
C2306 a_43262_21540# a_43262_20536# 1.00fF
C2307 a_30111_47911# a_30999_48071# 0.66fF
C2308 VDD a_27198_12504# 0.52fF
C2309 VDD a_5521_72373# 0.73fF
C2310 a_48282_16520# vcm 0.65fF
C2311 VDD a_18546_58180# 32.63fF
C2312 a_40250_13508# ctopn 3.58fF
C2313 cgen.dlycontrol2_in[0] a_12237_36596# 0.75fF
C2314 a_35230_57134# vcm 0.62fF
C2315 a_27603_34191# cgen.dlycontrol1_in[3] 0.62fF
C2316 VDD a_6265_37039# 0.65fF
C2317 a_34226_71190# vcm 0.60fF
C2318 a_38242_18528# ctopn 3.58fF
C2319 a_18546_12502# vcm 0.40fF
C2320 VDD a_25393_41317# 1.19fF
C2321 a_21174_58138# vcm 0.62fF
C2322 ANTENNA__1190__A2.DIODE a_10593_15823# 0.62fF
C2323 VDD a_17959_41001# 0.60fF
C2324 a_2007_25597# a_3325_26159# 0.37fF
C2325 ANTENNA__1190__B1.DIODE ANTENNA__1190__A2.DIODE 0.77fF
C2326 a_49286_15516# ctopn 3.57fF
C2327 VDD a_49286_11500# 0.52fF
C2328 ANTENNA__1395__B1.DIODE a_38913_31055# 0.83fF
C2329 VDD a_1591_15829# 0.44fF
C2330 a_30543_40721# a_12116_40871# 0.36fF
C2331 VDD nmat.col_n[31] 13.20fF
C2332 ANTENNA__1184__B1.DIODE a_18563_27791# 3.95fF
C2333 a_18546_69224# a_49194_69182# 0.35fF
C2334 VDD a_2163_31741# 0.50fF
C2335 nmat.col[6] m2_24960_24282# 0.39fF
C2336 pmat.col_n[19] ctopp 2.02fF
C2337 a_37238_11500# a_37238_10496# 1.00fF
C2338 VDD a_44763_34293# 1.66fF
C2339 VDD a_45178_72194# 0.32fF
C2340 a_38793_49007# nmat.col[15] 0.39fF
C2341 nmat.en_bit_n[1] nmat.col[15] 0.40fF
C2342 pmat.row_n[12] a_12263_50959# 0.37fF
C2343 cgen.dlycontrol3_in[0] a_11113_39747# 6.20fF
C2344 a_13091_28327# a_22199_30287# 0.46fF
C2345 a_2007_25597# nmat.col_n[1] 0.67fF
C2346 a_18546_9490# a_23090_9898# 0.35fF
C2347 pmat.rowon_n[11] pmat.rowoff_n[11] 21.06fF
C2348 a_46274_22544# vcm 0.65fF
C2349 a_42258_61150# a_43262_61150# 0.97fF
C2350 a_44266_68178# ctopp 3.58fF
C2351 a_12067_67279# a_12152_66415# 1.67fF
C2352 a_12309_38659# a_36161_37462# 0.50fF
C2353 a_22178_59142# vcm 0.62fF
C2354 VDD nmat.col[4] 4.93fF
C2355 a_27198_12504# a_27198_11500# 1.00fF
C2356 a_4128_64391# a_9963_13967# 3.73fF
C2357 m2_17932_15246# vcm 0.44fF
C2358 cgen.dlycontrol3_in[4] cgen.dlycontrol4_in[2] 0.90fF
C2359 a_24374_29941# nmat.col[10] 0.60fF
C2360 a_10515_75895# a_11823_74895# 0.39fF
C2361 cgen.dlycontrol1_in[1] cgen.dlycontrol1_in[0] 1.28fF
C2362 VDD a_26194_56130# 0.55fF
C2363 a_36234_20536# a_37238_20536# 0.97fF
C2364 a_6283_31591# a_28621_47381# 0.60fF
C2365 VDD a_7276_11739# 0.81fF
C2366 a_24591_28327# a_29937_31055# 0.33fF
C2367 a_18546_72236# a_22086_72194# 0.35fF
C2368 a_19405_28853# nmat.col_n[1] 0.71fF
C2369 VDD m2_40020_7214# 1.04fF
C2370 pmat.col[17] ctopp 2.01fF
C2371 a_13275_48783# a_7717_14735# 0.33fF
C2372 cgen.enable_dlycontrol_in a_11113_36483# 4.48fF
C2373 VDD a_4048_74549# 0.65fF
C2374 a_18546_62196# a_40158_62154# 0.35fF
C2375 VDD a_42292_47893# 0.39fF
C2376 pmat.rowon_n[11] nmat.rowon_n[5] 0.80fF
C2377 a_49286_67174# a_49286_66170# 1.00fF
C2378 a_18546_66212# a_36142_66170# 0.35fF
C2379 a_35230_9492# a_35230_8488# 1.00fF
C2380 VDD a_13798_22351# 0.47fF
C2381 a_20170_66170# ctopp 3.57fF
C2382 a_50290_63158# m2_51064_62978# 0.96fF
C2383 a_11067_64015# a_14839_54599# 0.48fF
C2384 VDD a_2953_33237# 0.31fF
C2385 VDD a_29206_66170# 0.52fF
C2386 a_50290_56130# m2_50060_54946# 0.99fF
C2387 VDD a_22178_63158# 0.52fF
C2388 ANTENNA__1190__A1.DIODE a_20439_27247# 1.32fF
C2389 a_48282_17524# a_49286_17524# 0.97fF
C2390 a_46274_57134# a_47278_57134# 0.97fF
C2391 a_25575_31055# clk_ena 1.30fF
C2392 a_18546_61192# a_21082_61150# 0.35fF
C2393 a_13459_28111# a_24407_31375# 0.69fF
C2394 ANTENNA__1395__B1.DIODE a_21739_29415# 1.03fF
C2395 a_45270_71190# a_46274_71190# 0.97fF
C2396 a_1923_31743# a_1591_27797# 0.57fF
C2397 a_9963_28111# a_9075_28023# 0.76fF
C2398 a_14641_57711# a_10055_31591# 0.30fF
C2399 VDD a_28116_38567# 1.26fF
C2400 cgen.dlycontrol4_in[5] a_2046_30184# 0.89fF
C2401 a_32218_58138# a_33222_58138# 0.97fF
C2402 nmat.rowon_n[7] a_11435_58791# 1.24fF
C2403 a_10515_15055# a_11067_16359# 1.11fF
C2404 VDD a_30913_44219# 1.30fF
C2405 a_19166_69182# m2_17932_69002# 0.96fF
C2406 a_22178_19532# vcm 0.65fF
C2407 a_49286_8488# a_50290_8488# 0.97fF
C2408 a_9411_2215# a_8861_24527# 0.45fF
C2409 VDD a_7619_30485# 0.58fF
C2410 a_11435_58791# a_14653_53458# 0.32fF
C2411 VDD a_11711_58261# 0.45fF
C2412 m3_19068_23410# ctopn 0.46fF
C2413 a_6467_29415# a_19541_28879# 2.57fF
C2414 a_11067_30287# a_29076_48695# 0.58fF
C2415 a_24591_28327# a_15667_27239# 1.42fF
C2416 a_21174_10496# vcm 0.65fF
C2417 VDD a_12967_12863# 0.42fF
C2418 a_22357_39141# a_22085_38550# 0.31fF
C2419 _1192_.B1 a_31263_28309# 0.34fF
C2420 a_49286_22544# ctopn 3.56fF
C2421 ANTENNA__1183__B1.DIODE nmat.col[18] 11.65fF
C2422 a_17139_30503# a_22199_30287# 1.56fF
C2423 VDD a_20503_48981# 0.35fF
C2424 pmat.row_n[8] a_18162_16520# 25.57fF
C2425 a_10515_15055# nmat.rowoff_n[13] 0.75fF
C2426 a_9135_60967# a_9231_32117# 0.33fF
C2427 a_4259_73807# a_4266_63303# 0.37fF
C2428 a_32218_61150# a_32218_60146# 1.00fF
C2429 VDD a_13559_23439# 0.37fF
C2430 a_40250_19532# a_40250_18528# 1.00fF
C2431 pmat.row_n[4] cgen.dlycontrol1_in[4] 0.66fF
C2432 a_18546_70228# a_38150_70186# 0.35fF
C2433 VDD a_27198_67174# 0.52fF
C2434 pmat.row_n[15] pmat.row_n[4] 2.43fF
C2435 ANTENNA__1195__A1.DIODE pmat.col[1] 2.51fF
C2436 VDD a_4127_37013# 0.81fF
C2437 a_20170_18528# ctopn 3.57fF
C2438 pmat.rowoff_n[7] ctopp 0.60fF
C2439 VDD a_20251_42089# 0.59fF
C2440 a_37238_62154# vcm 0.62fF
C2441 a_13091_52047# a_19541_28879# 1.01fF
C2442 a_28704_29568# nmat.col_n[21] 0.58fF
C2443 a_18546_17522# a_33130_17930# 0.35fF
C2444 a_3923_68021# a_9643_66389# 0.46fF
C2445 _1179_.X a_29937_31055# 1.19fF
C2446 a_18546_57176# a_29114_57134# 0.35fF
C2447 VDD a_10815_55785# 0.52fF
C2448 a_33222_59142# a_33222_58138# 1.00fF
C2449 a_18162_67214# vcm 6.95fF
C2450 a_50290_8488# m2_51064_8218# 0.96fF
C2451 a_39246_8488# m2_39016_7214# 1.00fF
C2452 a_6283_31591# a_25681_46831# 0.31fF
C2453 a_33423_47695# a_29937_31055# 0.50fF
C2454 pmat.rowoff_n[15] pmat.rowon_n[15] 20.82fF
C2455 a_2879_57487# a_4991_69831# 1.23fF
C2456 a_18546_15514# a_33130_15922# 0.35fF
C2457 a_25190_15516# a_26194_15516# 0.97fF
C2458 a_24186_69182# a_25190_69182# 0.97fF
C2459 a_13158_71285# a_3615_71631# 0.60fF
C2460 a_36234_70186# vcm 0.62fF
C2461 VDD pmat.col_n[12] 5.48fF
C2462 a_23182_11500# vcm 0.65fF
C2463 VDD m2_51064_17254# 1.00fF
C2464 VDD a_1591_18005# 0.41fF
C2465 a_38242_17524# a_38242_16520# 1.00fF
C2466 a_2648_29397# a_2021_9563# 0.89fF
C2467 VDD a_20078_24958# 0.39fF
C2468 ANTENNA__1197__B.DIODE _1183_.A2 16.96fF
C2469 pmat.row_n[14] pmat.row_n[0] 1.18fF
C2470 VDD config_2_in[10] 1.21fF
C2471 a_44266_12504# a_45270_12504# 0.97fF
C2472 ANTENNA__1190__A1.DIODE a_27763_27221# 1.46fF
C2473 a_25190_19532# ctopn 3.58fF
C2474 a_21395_50857# a_10883_3303# 0.48fF
C2475 a_1591_27797# a_1757_27797# 0.60fF
C2476 VDD a_18546_15514# 32.63fF
C2477 nmat.rowon_n[9] a_18162_14512# 1.33fF
C2478 VDD a_25190_21540# 0.52fF
C2479 a_5363_33551# nmat.col_n[12] 1.13fF
C2480 a_18546_59184# a_49194_59142# 0.35fF
C2481 a_33222_59142# a_34226_59142# 0.97fF
C2482 a_24186_10496# ctopn 3.58fF
C2483 a_45270_57134# ctopp 3.57fF
C2484 pmat.row_n[12] pmat.rowon_n[11] 1.04fF
C2485 a_44266_71190# ctopp 3.40fF
C2486 VDD a_3225_55509# 0.63fF
C2487 a_31214_58138# ctopp 3.58fF
C2488 a_27198_68178# vcm 0.62fF
C2489 a_37820_30485# a_31675_47695# 0.32fF
C2490 VDD result_out[3] 0.73fF
C2491 pmat.rowoff_n[7] a_1586_50247# 0.40fF
C2492 nmat.rowon_n[5] a_18162_18528# 1.33fF
C2493 VDD a_40250_58138# 0.52fF
C2494 nmat.sw a_9411_2215# 0.60fF
C2495 a_22178_23548# a_22178_22544# 1.00fF
C2496 a_21174_60146# a_22178_60146# 0.97fF
C2497 a_18546_60188# a_25098_60146# 0.35fF
C2498 pmat.col_n[7] a_24867_53135# 0.34fF
C2499 a_11339_39319# a_11681_35823# 2.12fF
C2500 VDD a_1591_65327# 0.85fF
C2501 a_16311_28327# pmat.col[8] 0.39fF
C2502 a_26891_28327# a_22199_30287# 0.69fF
C2503 a_18563_27791# a_13641_23439# 0.61fF
C2504 VDD a_3045_19093# 0.35fF
C2505 nmat.col[29] nmat.col_n[28] 6.80fF
C2506 a_29206_68178# a_29206_67174# 1.00fF
C2507 a_32218_23548# vcm 0.65fF
C2508 a_23182_69182# ctopp 3.58fF
C2509 m2_51064_56954# m2_51064_55950# 0.99fF
C2510 a_4991_69831# a_7730_69109# 0.79fF
C2511 a_34226_9492# vcm 0.65fF
C2512 VDD a_32218_69182# 0.52fF
C2513 VDD a_21371_50087# 7.02fF
C2514 a_49286_23548# m2_49056_24282# 0.99fF
C2515 a_18546_22542# a_51202_22950# 0.35fF
C2516 a_11067_30287# a_13479_26935# 0.66fF
C2517 VDD a_31978_43439# 0.52fF
C2518 VDD a_26155_46831# 0.39fF
C2519 a_22365_32149# a_18241_31698# 0.58fF
C2520 pmat.rowon_n[0] a_2835_13077# 0.70fF
C2521 a_50290_20536# vcm 0.65fF
C2522 nmat.sw a_15049_36374# 1.30fF
C2523 a_32218_59142# ctopp 3.58fF
C2524 a_26194_11500# ctopn 3.58fF
C2525 VDD a_45589_31599# 0.34fF
C2526 a_10515_61839# nmat.rowoff_n[14] 0.71fF
C2527 VDD a_41254_59142# 0.52fF
C2528 VDD a_1591_56623# 1.16fF
C2529 VDD a_17959_35561# 0.60fF
C2530 pmat.rowon_n[6] ctopp 1.57fF
C2531 a_10441_21263# nmat.col[0] 0.34fF
C2532 a_1674_57711# pmat.rowoff_n[7] 0.31fF
C2533 pmat.sw a_2952_25045# 0.35fF
C2534 a_2263_43719# a_15899_47939# 0.42fF
C2535 a_19584_52423# a_11711_50959# 0.38fF
C2536 nmat.rowoff_n[6] a_12245_21807# 0.46fF
C2537 a_27198_16520# a_28202_16520# 0.97fF
C2538 a_18546_16518# a_37146_16926# 0.35fF
C2539 nmat.col[19] vcm 8.27fF
C2540 a_18546_70228# a_20078_70186# 0.35fF
C2541 a_7415_29397# a_9075_28023# 0.96fF
C2542 a_30210_13508# vcm 0.65fF
C2543 VDD a_14497_42658# 1.69fF
C2544 a_19166_62154# vcm 0.61fF
C2545 m2_46044_7214# m2_47048_7214# 0.96fF
C2546 cgen.dlycontrol3_in[4] a_12228_40693# 3.63fF
C2547 a_28202_18528# vcm 0.65fF
C2548 VDD a_18484_29967# 0.44fF
C2549 a_12815_74581# a_12981_74581# 0.75fF
C2550 a_30571_50959# nmat.col_n[21] 0.47fF
C2551 a_12235_39913# a_12228_39605# 0.41fF
C2552 a_6283_31591# a_29937_31055# 0.37fF
C2553 VDD a_1959_10615# 0.52fF
C2554 pmat.row_n[15] a_3305_27791# 1.15fF
C2555 VDD m3_35132_72146# 0.40fF
C2556 nmat.rowon_n[7] a_12044_49641# 0.31fF
C2557 a_10515_15055# a_11067_49871# 0.48fF
C2558 a_39246_15516# vcm 0.65fF
C2559 VDD a_24186_17524# 0.52fF
C2560 VDD a_4409_74183# 0.58fF
C2561 ANTENNA__1395__A1.DIODE ANTENNA__1197__B.DIODE 1.89fF
C2562 VDD a_18162_22544# 2.74fF
C2563 a_36234_70186# a_36234_69182# 1.00fF
C2564 VDD a_25190_8488# 0.55fF
C2565 a_18546_21538# a_28110_21946# 0.35fF
C2566 VDD a_46636_36469# 0.40fF
C2567 a_18546_70228# vcm 0.40fF
C2568 VDD a_9871_53903# 0.31fF
C2569 a_25190_14512# a_25190_13508# 1.00fF
C2570 VDD a_34705_51959# 1.32fF
C2571 a_25575_31055# a_27001_30511# 1.59fF
C2572 a_35230_23548# ctopn 3.51fF
C2573 VDD a_41254_19532# 0.52fF
C2574 a_37238_9492# ctopn 3.57fF
C2575 m2_20944_24282# m3_21076_24414# 2.79fF
C2576 _1194_.A2 ANTENNA__1190__B1.DIODE 6.63fF
C2577 ANTENNA__1197__A.DIODE ANTENNA__1190__A1.DIODE 0.86fF
C2578 a_29206_57134# a_29206_56130# 1.00fF
C2579 a_25695_28111# a_7717_14735# 1.13fF
C2580 pmat.col[0] a_15667_27239# 1.60fF
C2581 pmat.row_n[14] nmat.sample 0.34fF
C2582 a_33222_19532# a_34226_19532# 0.97fF
C2583 a_35230_60146# vcm 0.62fF
C2584 VDD a_40250_10496# 0.52fF
C2585 a_10873_38517# a_22537_36911# 0.95fF
C2586 a_10515_61839# a_11067_16359# 1.90fF
C2587 a_18243_28327# clk_ena 0.63fF
C2588 a_10515_13967# a_7644_16341# 0.37fF
C2589 pmat.col_n[21] m2_40020_54946# 0.37fF
C2590 VDD dummypin[7] 1.01fF
C2591 VDD a_1895_20346# 0.53fF
C2592 pmat.col[29] m2_48052_54946# 0.39fF
C2593 a_1923_31743# a_2787_33237# 0.35fF
C2594 a_18546_58180# a_47186_58138# 0.35fF
C2595 a_6795_76989# a_6975_76823# 2.53fF
C2596 VDD nmat.col[10] 8.99fF
C2597 VDD m2_17932_18258# 1.00fF
C2598 a_4259_31375# a_9307_31068# 0.31fF
C2599 a_32218_10496# a_33222_10496# 0.97fF
C2600 a_18546_10494# a_47186_10902# 0.35fF
C2601 a_21215_48071# a_15899_47939# 0.32fF
C2602 a_38391_48469# a_38557_48469# 0.42fF
C2603 a_47278_62154# ctopp 3.58fF
C2604 a_41254_16520# vcm 0.65fF
C2605 a_10883_3303# nmat.rowon_n[2] 0.43fF
C2606 a_10515_61839# nmat.rowoff_n[13] 0.72fF
C2607 a_43262_56130# a_44266_56130# 0.97fF
C2608 a_5731_58951# a_3746_58487# 0.54fF
C2609 pmat.row_n[4] pmat.rowon_n[3] 0.33fF
C2610 a_19166_18528# a_20170_18528# 0.97fF
C2611 a_33222_13508# ctopn 3.58fF
C2612 a_12263_50959# a_18547_51565# 1.03fF
C2613 a_28202_57134# vcm 0.62fF
C2614 VDD a_34887_38007# 0.63fF
C2615 a_27198_71190# vcm 0.60fF
C2616 a_31214_18528# ctopn 3.58fF
C2617 VDD a_1895_41018# 0.53fF
C2618 pmat.rowon_n[0] a_13091_7655# 0.34fF
C2619 inn_analog ANTENNA__1190__A2.DIODE 1.47fF
C2620 a_24861_29673# a_10147_29415# 1.27fF
C2621 VDD a_4533_38279# 1.17fF
C2622 a_28704_29568# clk_ena 0.86fF
C2623 a_46274_70186# ctopp 3.57fF
C2624 VDD a_14163_55295# 0.37fF
C2625 a_20170_63158# pmat.col[1] 0.31fF
C2626 a_42258_15516# ctopn 3.58fF
C2627 pmat.col_n[31] clk_ena 0.56fF
C2628 VDD a_42258_11500# 0.52fF
C2629 a_25190_22544# a_26194_22544# 0.97fF
C2630 a_32687_46607# a_2007_25597# 0.34fF
C2631 a_48282_62154# a_49286_62154# 0.97fF
C2632 m2_51064_12234# m2_51064_11230# 0.99fF
C2633 pmat.rowoff_n[7] cgen.start_conv_in 0.83fF
C2634 a_2021_26677# rst_n 0.41fF
C2635 VDD a_9213_53903# 1.18fF
C2636 nmat.col[10] nmat.rowoff_n[2] 4.53fF
C2637 a_46274_66170# a_47278_66170# 0.97fF
C2638 pmat.row_n[4] a_2648_29397# 3.05fF
C2639 pmat.rowon_n[7] pmat.rowoff_n[7] 20.57fF
C2640 a_5363_70543# a_9405_66627# 0.58fF
C2641 a_18546_69224# a_42166_69182# 0.35fF
C2642 VDD a_38727_32447# 0.32fF
C2643 VDD a_8105_7125# 0.67fF
C2644 VDD a_24937_36039# 1.22fF
C2645 a_25839_49783# a_13275_48783# 1.11fF
C2646 a_18162_17524# ctopn 1.49fF
C2647 _1154_.X nmat.col[19] 0.47fF
C2648 a_21739_29415# nmat.col[18] 1.02fF
C2649 VDD a_17007_50613# 0.30fF
C2650 a_4719_30287# a_4533_38279# 0.92fF
C2651 a_24591_28327# a_11067_27239# 0.46fF
C2652 ANTENNA__1184__B1.DIODE _1194_.B1 1.72fF
C2653 ANTENNA__1197__B.DIODE ANTENNA__1395__A2.DIODE 0.86fF
C2654 a_39246_63158# a_40250_63158# 0.97fF
C2655 m2_51064_55950# vcm 0.51fF
C2656 a_7026_24527# nmat.col_n[1] 0.52fF
C2657 a_39246_22544# vcm 0.65fF
C2658 a_37238_68178# ctopp 3.58fF
C2659 a_35230_55126# m3_35132_55078# 1.39fF
C2660 VDD a_46274_68178# 0.52fF
C2661 VDD a_12213_53359# 0.41fF
C2662 pmat.col_n[14] vcm 2.80fF
C2663 VDD a_25061_43132# 1.18fF
C2664 a_18546_14510# a_20078_14918# 0.35fF
C2665 a_50290_69182# m2_51064_69002# 0.96fF
C2666 a_18546_20534# a_48190_20942# 0.35fF
C2667 a_44266_16520# ctopn 3.58fF
C2668 a_14887_46377# a_32687_46607# 2.34fF
C2669 VDD a_2283_27221# 1.18fF
C2670 VDD m2_25964_7214# 0.93fF
C2671 VDD a_10515_75895# 2.44fF
C2672 a_18546_62196# a_33130_62154# 0.35fF
C2673 a_13091_28327# a_34942_51701# 0.32fF
C2674 VDD a_8079_46519# 0.66fF
C2675 a_18546_66212# a_29114_66170# 0.35fF
C2676 pmat.col_n[15] ANTENNA__1197__B.DIODE 0.35fF
C2677 a_47278_70186# a_48282_70186# 0.97fF
C2678 VDD a_22178_66170# 0.52fF
C2679 VDD a_1591_8213# 0.41fF
C2680 a_24867_53135# a_28915_50959# 1.60fF
C2681 a_18546_11498# a_51202_11906# 0.35fF
C2682 a_9675_10396# a_12705_10389# 0.59fF
C2683 a_34226_11500# a_35230_11500# 0.97fF
C2684 VDD a_1757_36501# 0.62fF
C2685 a_2315_44124# a_2659_35015# 0.51fF
C2686 ANTENNA_fanout52_A.DIODE vcm 0.75fF
C2687 a_7415_29397# a_33515_31055# 0.42fF
C2688 a_20170_17524# a_20170_16520# 1.00fF
C2689 a_36234_64162# a_36234_63158# 1.00fF
C2690 m2_29980_54946# m3_30112_55078# 2.79fF
C2691 a_6927_30503# a_6559_33767# 0.59fF
C2692 a_39246_10496# a_39246_9492# 1.00fF
C2693 a_6634_26133# a_5320_27023# 0.43fF
C2694 m2_17932_54946# m2_18936_54946# 0.96fF
C2695 a_36234_58138# a_36234_57134# 1.00fF
C2696 a_3339_59879# a_10239_77295# 0.34fF
C2697 a_1923_69823# a_7658_71543# 0.78fF
C2698 a_47278_14512# vcm 0.65fF
C2699 a_46274_64162# vcm 0.62fF
C2700 a_2007_25597# a_37471_32149# 0.57fF
C2701 a_40250_60146# a_40250_59142# 1.00fF
C2702 a_28202_18528# a_28202_17524# 1.00fF
C2703 a_19166_58138# vcm 0.61fF
C2704 VDD a_45396_31849# 0.39fF
C2705 a_12309_36483# a_11921_35286# 2.64fF
C2706 pmat.row_n[4] nmat.rowoff_n[5] 0.38fF
C2707 VDD pmat.rowon_n[1] 3.91fF
C2708 _1179_.X a_11067_27239# 0.60fF
C2709 ANTENNA_fanout52_A.DIODE _1194_.B1 3.57fF
C2710 ANTENNA__1197__B.DIODE ANTENNA__1196__A2.DIODE 0.79fF
C2711 a_24867_53135# ANTENNA__1395__B1.DIODE 1.14fF
C2712 _1192_.B1 a_21739_29415# 0.33fF
C2713 VDD a_49286_13508# 0.52fF
C2714 pmat.rowon_n[0] cgen.dlycontrol2_in[2] 0.38fF
C2715 a_42258_22544# ctopn 3.57fF
C2716 cgen.dlycontrol4_in[4] a_11497_40719# 0.45fF
C2717 VDD a_47278_18528# 0.52fF
C2718 a_28202_63158# a_28202_62154# 1.00fF
C2719 VDD a_37820_30485# 5.89fF
C2720 pmat.row_n[6] ANTENNA__1196__A2.DIODE 0.58fF
C2721 pmat.col[13] vcm 5.88fF
C2722 a_44266_67174# a_45270_67174# 0.97fF
C2723 a_18546_70228# a_31122_70186# 0.35fF
C2724 VDD a_20170_67174# 0.52fF
C2725 VDD a_5325_9269# 0.57fF
C2726 a_3615_71631# a_11435_58791# 1.58fF
C2727 a_33423_47695# a_35312_31599# 4.38fF
C2728 a_2411_43301# cgen.dlycontrol4_in[5] 0.71fF
C2729 a_34226_22544# a_34226_21540# 1.00fF
C2730 a_41254_66170# a_41254_65166# 1.00fF
C2731 _1154_.X ANTENNA__1184__B1.DIODE 1.15fF
C2732 VDD _1183_.A2 25.11fF
C2733 VDD a_38927_42359# 0.57fF
C2734 a_33222_14512# a_34226_14512# 0.97fF
C2735 a_18546_14510# a_49194_14918# 0.35fF
C2736 a_30210_62154# vcm 0.62fF
C2737 a_14653_53458# a_19541_28879# 0.51fF
C2738 a_18546_17522# a_26102_17930# 0.35fF
C2739 a_18546_64204# a_47186_64162# 0.35fF
C2740 a_32218_64162# a_33222_64162# 0.97fF
C2741 a_38242_68178# a_39246_68178# 0.97fF
C2742 a_2124_74299# a_2163_74173# 0.79fF
C2743 a_18546_57176# a_22086_57134# 0.35fF
C2744 a_4339_27804# clk_dig 1.54fF
C2745 a_14533_39631# a_19409_40719# 0.46fF
C2746 a_27198_13508# a_27198_12504# 1.00fF
C2747 a_11435_58791# a_2952_25045# 0.44fF
C2748 ANTENNA__1395__A2.DIODE a_14691_27399# 0.38fF
C2749 a_18546_15514# a_26102_15922# 0.35fF
C2750 a_49286_65166# vcm 0.62fF
C2751 a_45270_60146# ctopp 3.58fF
C2752 m2_44036_72014# m3_44168_72146# 2.79fF
C2753 VDD a_3956_59317# 0.39fF
C2754 a_6451_67655# a_5307_67655# 1.63fF
C2755 a_29206_70186# vcm 0.62fF
C2756 a_25839_49783# a_25850_48981# 0.90fF
C2757 pmat.en_bit_n[0] a_17702_29967# 0.52fF
C2758 a_20310_28029# a_10441_21263# 0.69fF
C2759 a_14943_26703# nmat.col[7] 0.37fF
C2760 nmat.col[30] nmat.col[21] 0.62fF
C2761 m2_17932_56954# vcm 0.44fF
C2762 VDD a_12463_22351# 1.12fF
C2763 a_19166_68178# ctopp 3.43fF
C2764 pmat.row_n[13] a_14641_57167# 0.63fF
C2765 a_50290_14512# ctopn 3.43fF
C2766 a_2199_13887# a_5654_9527# 0.30fF
C2767 a_8197_20871# a_8305_20871# 0.35fF
C2768 a_1781_9308# a_9963_28111# 0.71fF
C2769 VDD a_3229_14741# 0.66fF
C2770 a_4351_55527# a_6451_67655# 0.37fF
C2771 a_18546_59184# a_42166_59142# 0.35fF
C2772 a_34226_65166# a_34226_64162# 1.00fF
C2773 a_4075_31591# a_13091_7655# 0.35fF
C2774 a_1923_53055# a_2163_56765# 0.35fF
C2775 pmat.col[15] ctopp 1.99fF
C2776 pmat.rowoff_n[8] a_13091_52047# 0.56fF
C2777 a_38242_57134# ctopp 3.57fF
C2778 VDD a_34204_27765# 1.97fF
C2779 pmat.col_n[19] _1187_.A2 0.43fF
C2780 a_37238_71190# ctopp 3.40fF
C2781 VDD a_47278_57134# 0.52fF
C2782 a_24186_58138# ctopp 3.58fF
C2783 a_20170_68178# vcm 0.62fF
C2784 VDD a_46274_71190# 0.55fF
C2785 VDD a_33222_58138# 0.52fF
C2786 VDD a_14439_72703# 0.36fF
C2787 a_43262_23548# a_44266_23548# 0.97fF
C2788 a_23182_16520# a_23182_15516# 1.00fF
C2789 a_45270_9492# a_46274_9492# 0.97fF
C2790 pmat.row_n[4] a_5363_33551# 0.36fF
C2791 _1154_.X ANTENNA_fanout52_A.DIODE 2.09fF
C2792 pmat.row_n[11] a_5271_35407# 0.32fF
C2793 pmat.row_n[9] a_14825_50095# 0.59fF
C2794 VDD a_11007_58229# 1.37fF
C2795 cgen.dlycontrol2_in[0] a_14773_37218# 0.54fF
C2796 pmat.col[23] vcm 5.88fF
C2797 a_11067_64015# a_9983_32385# 0.63fF
C2798 a_11041_40948# a_11297_36091# 0.44fF
C2799 a_2263_43719# cgen.dlycontrol3_in[4] 1.41fF
C2800 a_33222_56130# m2_32992_54946# 0.99fF
C2801 ANTENNA__1395__B1.DIODE a_38851_28327# 1.54fF
C2802 a_18546_24550# a_47186_24958# 0.35fF
C2803 nmat.en_bit_n[0] a_22628_30485# 0.94fF
C2804 VDD a_30913_39867# 1.55fF
C2805 a_25190_23548# vcm 0.65fF
C2806 a_19166_65166# m2_17932_64986# 0.96fF
C2807 a_6200_70919# a_2407_49289# 0.83fF
C2808 a_27198_9492# vcm 0.65fF
C2809 VDD a_25190_69182# 0.52fF
C2810 a_49286_61150# vcm 0.62fF
C2811 _1224_.X clk_vcm 0.46fF
C2812 a_18546_22542# a_44174_22950# 0.35fF
C2813 VDD config_1_in[12] 1.41fF
C2814 a_1957_43567# a_1739_47893# 0.77fF
C2815 VDD m2_23956_24282# 0.62fF
C2816 VDD nmat.rowon_n[12] 19.54fF
C2817 a_43262_20536# vcm 0.65fF
C2818 pmat.rowon_n[7] a_11067_64015# 0.87fF
C2819 a_35230_65166# a_36234_65166# 0.97fF
C2820 a_25190_59142# ctopp 3.58fF
C2821 a_35244_32411# a_41949_30761# 1.11fF
C2822 a_18162_11500# ctopn 1.49fF
C2823 a_14287_70543# pmat.row_n[10] 1.08fF
C2824 VDD ANTENNA__1395__A1.DIODE 16.76fF
C2825 VDD a_34226_59142# 0.52fF
C2826 pmat.col_n[22] ctopp 2.02fF
C2827 a_21371_50087# a_22499_49783# 1.53fF
C2828 a_10883_3303# a_20475_49783# 0.50fF
C2829 a_42258_21540# a_43262_21540# 0.97fF
C2830 VDD a_5823_34863# 0.40fF
C2831 a_82863_64213# _1224_.X 0.48fF
C2832 VDD a_48190_72194# 0.32fF
C2833 a_10441_21263# a_9741_28585# 0.41fF
C2834 VDD config_2_in[4] 0.85fF
C2835 a_18546_16518# a_30118_16926# 0.35fF
C2836 a_5087_18543# a_5253_18543# 0.69fF
C2837 a_43262_71190# a_43262_70186# 1.00fF
C2838 VDD a_10499_67503# 0.34fF
C2839 pmat.col[0] m2_18936_54946# 0.39fF
C2840 a_23182_13508# vcm 0.65fF
C2841 pmat.rowon_n[11] a_18546_19530# 4.09fF
C2842 m2_39016_7214# m2_40020_7214# 0.96fF
C2843 a_10883_3303# a_25802_48169# 0.38fF
C2844 a_21174_18528# vcm 0.65fF
C2845 pmat.rowon_n[1] pmat.rowoff_n[1] 20.66fF
C2846 a_18823_50247# a_11711_50959# 0.55fF
C2847 a_4259_73807# a_4351_55527# 0.57fF
C2848 a_7658_71543# a_11232_73211# 0.60fF
C2849 a_4976_16091# a_7131_19407# 0.40fF
C2850 a_26891_28327# a_18563_27791# 0.65fF
C2851 m2_17932_58962# m2_17932_57958# 0.99fF
C2852 a_41254_13508# a_42258_13508# 0.97fF
C2853 _1154_.X a_25681_28879# 0.39fF
C2854 a_18546_72236# a_25098_72194# 0.35fF
C2855 a_32218_15516# vcm 0.65fF
C2856 VDD a_11881_16911# 0.49fF
C2857 _1179_.X _1196_.B1 6.89fF
C2858 VDD m2_51064_58962# 1.14fF
C2859 a_2787_33237# a_2953_33237# 0.72fF
C2860 a_10878_58487# pmat.rowon_n[3] 0.32fF
C2861 a_10239_14183# a_6467_29415# 0.86fF
C2862 a_39246_18528# a_40250_18528# 0.97fF
C2863 VDD a_3866_57399# 3.83fF
C2864 a_26194_62154# a_26194_61150# 1.00fF
C2865 nmat.col_n[29] vcm 4.09fF
C2866 a_28202_23548# ctopn 3.40fF
C2867 VDD a_34226_19532# 0.52fF
C2868 a_30210_9492# ctopn 3.57fF
C2869 VDD m2_43032_72014# 1.39fF
C2870 nmat.col[24] nmat.col_n[30] 8.32fF
C2871 a_40105_47375# a_43720_32143# 1.26fF
C2872 a_28202_60146# vcm 0.62fF
C2873 _1179_.X a_9785_28879# 0.39fF
C2874 VDD a_33222_10496# 0.52fF
C2875 ANTENNA__1184__B1.DIODE nmat.col_n[7] 1.15fF
C2876 m2_17932_72014# m2_17932_71010# 0.99fF
C2877 VDD a_36341_39141# 1.47fF
C2878 VDD result_out[14] 0.80fF
C2879 a_46274_20536# ctopn 3.58fF
C2880 a_26194_15516# a_26194_14512# 1.00fF
C2881 a_18546_58180# a_40158_58138# 0.35fF
C2882 a_49286_69182# a_50290_69182# 0.97fF
C2883 a_28202_69182# a_28202_68178# 1.00fF
C2884 a_3866_57399# a_4719_30287# 0.45fF
C2885 a_19166_71190# ctopp 3.24fF
C2886 a_4075_31591# nmat.sw 0.36fF
C2887 a_18546_10494# a_40158_10902# 0.35fF
C2888 a_36234_21540# a_36234_20536# 1.00fF
C2889 a_4075_50087# a_5682_56311# 0.54fF
C2890 a_40250_62154# ctopp 3.58fF
C2891 VDD a_49286_62154# 0.52fF
C2892 a_25681_28879# a_27995_30287# 0.75fF
C2893 a_34226_16520# vcm 0.65fF
C2894 a_11041_39860# cgen.dlycontrol4_in[1] 3.78fF
C2895 nmat.col[15] a_35244_32411# 0.35fF
C2896 VDD a_44774_48695# 0.76fF
C2897 a_4843_54826# a_1769_47919# 0.44fF
C2898 VDD ANTENNA__1395__A2.DIODE 16.64fF
C2899 a_26194_13508# ctopn 3.58fF
C2900 VDD a_34887_40183# 0.64fF
C2901 a_21174_57134# vcm 0.62fF
C2902 VDD a_20848_38341# 1.14fF
C2903 a_20170_71190# vcm 0.60fF
C2904 a_24186_18528# ctopn 3.58fF
C2905 VDD a_28999_42089# 0.63fF
C2906 pmat.row_n[2] a_16083_50069# 0.70fF
C2907 VDD a_18162_64202# 2.74fF
C2908 a_14917_23983# a_9785_28879# 1.83fF
C2909 VDD a_44382_40847# 1.09fF
C2910 a_39246_70186# ctopp 3.57fF
C2911 a_14839_20871# a_8861_24527# 0.40fF
C2912 VDD a_48282_70186# 0.52fF
C2913 a_35230_15516# ctopn 3.58fF
C2914 VDD a_35230_11500# 0.52fF
C2915 a_32218_23548# m2_31988_24282# 0.99fF
C2916 a_47278_23548# a_47278_22544# 1.00fF
C2917 VDD a_1849_45205# 0.64fF
C2918 a_46274_60146# a_47278_60146# 0.97fF
C2919 a_4075_68583# a_2315_44124# 0.37fF
C2920 a_18546_69224# a_35138_69182# 0.35fF
C2921 VDD a_3938_58229# 0.80fF
C2922 a_30210_11500# a_30210_10496# 1.00fF
C2923 a_50290_56130# vcm 0.62fF
C2924 VDD pmat.col_n[15] 4.97fF
C2925 VDD a_2499_13077# 0.44fF
C2926 VDD a_6175_60039# 2.74fF
C2927 a_2835_13077# a_2907_22522# 0.33fF
C2928 _1194_.A2 a_12263_50959# 0.48fF
C2929 a_4068_25615# a_3305_27791# 0.36fF
C2930 a_3325_36495# a_4127_37013# 0.63fF
C2931 a_32218_22544# vcm 0.65fF
C2932 a_35230_61150# a_36234_61150# 0.97fF
C2933 a_30210_68178# ctopp 3.58fF
C2934 VDD a_39246_68178# 0.52fF
C2935 pmat.rowon_n[3] cgen.dlycontrol4_in[1] 2.34fF
C2936 a_32687_46607# nmat.col_n[21] 0.43fF
C2937 VDD a_6173_42479# 0.57fF
C2938 a_46274_63158# vcm 0.62fF
C2939 ANTENNA__1190__A1.DIODE nmat.col[19] 0.42fF
C2940 a_16113_52271# pmat.rowoff_n[3] 0.34fF
C2941 a_3938_58229# a_4719_30287# 0.30fF
C2942 _1196_.B1 a_6830_22895# 0.34fF
C2943 _1196_.B1 pmat.col[0] 0.33fF
C2944 ANTENNA__1395__B1.DIODE pmat.col[28] 0.32fF
C2945 a_29206_20536# a_30210_20536# 0.97fF
C2946 a_18546_20534# a_41162_20942# 0.35fF
C2947 a_37238_16520# ctopn 3.58fF
C2948 a_6175_60039# a_4719_30287# 0.82fF
C2949 _1154_.A vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.30fF
C2950 a_6451_67655# a_3615_71631# 0.62fF
C2951 VDD ANTENNA__1196__A2.DIODE 26.95fF
C2952 a_10873_39605# cgen.dlycontrol2_in[4] 2.07fF
C2953 _1183_.A2 a_7840_27247# 0.88fF
C2954 a_18546_62196# a_26102_62154# 0.35fF
C2955 m2_51064_20266# vcm 0.51fF
C2956 a_42258_67174# a_42258_66170# 1.00fF
C2957 a_18546_66212# a_22086_66170# 0.35fF
C2958 a_9668_10651# comp_latch 0.39fF
C2959 _1154_.X nmat.col_n[29] 0.74fF
C2960 a_28202_9492# a_28202_8488# 1.00fF
C2961 pmat.rowon_n[3] nmat.rowoff_n[3] 0.34fF
C2962 a_10883_3303# ANTENNA__1183__B1.DIODE 0.43fF
C2963 a_4259_31375# a_11067_30287# 1.60fF
C2964 pmat.col_n[9] nmat.en_bit_n[1] 0.47fF
C2965 VDD a_44266_23548# 0.55fF
C2966 VDD a_46274_9492# 0.52fF
C2967 VDD a_18546_60188# 32.63fF
C2968 a_18546_11498# a_44174_11906# 0.35fF
C2969 VDD a_32947_37737# 0.60fF
C2970 a_13432_62581# a_12429_62607# 0.61fF
C2971 a_10515_61839# pmat.rowoff_n[5] 0.42fF
C2972 VDD a_82818_69135# 1.62fF
C2973 nmat.rowon_n[2] a_10839_11989# 0.49fF
C2974 a_41254_17524# a_42258_17524# 0.97fF
C2975 a_39246_57134# a_40250_57134# 0.97fF
C2976 nmat.col_n[26] nmat.col_n[24] 0.33fF
C2977 a_8385_51727# a_9463_50877# 0.39fF
C2978 a_44266_20536# a_44266_19532# 1.00fF
C2979 cgen.dlycontrol1_in[2] clk_ena 4.36fF
C2980 a_38242_71190# a_39246_71190# 0.97fF
C2981 ANTENNA__1197__B.DIODE a_19405_28853# 0.65fF
C2982 a_5547_77295# a_1923_69823# 0.60fF
C2983 a_25190_58138# a_26194_58138# 0.97fF
C2984 a_40250_14512# vcm 0.65fF
C2985 cgen.dlycontrol2_in[3] a_3983_41941# 0.58fF
C2986 a_39246_64162# vcm 0.62fF
C2987 VDD m2_47048_24282# 0.62fF
C2988 VDD a_41926_46983# 1.55fF
C2989 a_42258_8488# a_43262_8488# 0.97fF
C2990 a_36234_62154# pmat.col[17] 0.31fF
C2991 VDD a_11337_25071# 1.51fF
C2992 _1194_.B1 a_13091_28327# 2.04fF
C2993 a_4025_54965# pmat.rowon_n[3] 0.30fF
C2994 VDD a_42258_13508# 0.52fF
C2995 a_50290_14512# a_50290_13508# 1.00fF
C2996 a_1591_38677# a_1757_38677# 0.75fF
C2997 pmat.row_n[12] pmat.row_n[9] 1.95fF
C2998 a_35230_22544# ctopn 3.58fF
C2999 cgen.dlycontrol4_in[3] a_2021_26677# 2.68fF
C3000 VDD a_40250_18528# 0.52fF
C3001 a_37820_30485# a_43533_30761# 0.99fF
C3002 m2_28976_24282# vcm 0.42fF
C3003 a_25190_61150# a_25190_60146# 1.00fF
C3004 nmat.col[30] nmat.col_n[28] 5.08fF
C3005 a_33222_19532# a_33222_18528# 1.00fF
C3006 a_18546_70228# a_24094_70186# 0.35fF
C3007 _1187_.A2 _1192_.A2 2.14fF
C3008 a_24867_53135# _1192_.B1 0.33fF
C3009 a_18546_14510# a_42166_14918# 0.35fF
C3010 a_23182_62154# vcm 0.62fF
C3011 _1184_.A2 nmat.col[1] 0.31fF
C3012 a_18546_64204# a_40158_64162# 0.35fF
C3013 a_39246_62154# pmat.col[20] 0.31fF
C3014 a_11051_8903# a_11731_8751# 0.34fF
C3015 a_26194_59142# a_26194_58138# 1.00fF
C3016 a_2263_43719# a_13091_18535# 0.45fF
C3017 _1224_.X ANTENNA__1195__A1.DIODE 0.54fF
C3018 VDD a_7099_74313# 0.83fF
C3019 a_42258_65166# vcm 0.62fF
C3020 a_23395_53135# a_24867_53135# 0.77fF
C3021 ANTENNA__1190__A1.DIODE ANTENNA__1184__B1.DIODE 0.75fF
C3022 VDD a_8453_46287# 0.39fF
C3023 a_7415_29397# a_12987_26159# 0.42fF
C3024 cgen.dlycontrol3_in[1] a_3325_40847# 0.33fF
C3025 a_49286_21540# vcm 0.65fF
C3026 a_10515_13967# pmat.rowon_n[3] 0.77fF
C3027 cgen.dlycontrol4_in[3] a_2839_38101# 1.01fF
C3028 a_38242_60146# ctopp 3.58fF
C3029 VDD a_47278_60146# 0.52fF
C3030 VDD a_12069_36341# 3.20fF
C3031 a_22178_70186# vcm 0.62fF
C3032 a_9411_2215# a_41731_49525# 0.46fF
C3033 cgen.enable_dlycontrol_in config_2_in[15] 0.56fF
C3034 a_23021_29199# a_16478_29423# 1.41fF
C3035 nmat.rowon_n[6] vcm 0.53fF
C3036 a_31214_17524# a_31214_16520# 1.00fF
C3037 m2_25964_24282# m3_26096_24414# 2.79fF
C3038 cgen.dlycontrol3_in[1] cgen.dlycontrol3_in[0] 1.73fF
C3039 a_50290_65166# m2_51064_64986# 0.96fF
C3040 a_43262_14512# ctopn 3.58fF
C3041 a_37238_12504# a_38242_12504# 0.97fF
C3042 a_22199_30287# a_25879_31591# 2.00fF
C3043 VDD a_17996_41831# 1.29fF
C3044 nmat.sample_n a_9785_28879# 1.00fF
C3045 VDD a_13655_26703# 0.65fF
C3046 a_26194_59142# a_27198_59142# 0.97fF
C3047 a_18546_59184# a_35138_59142# 0.35fF
C3048 a_18243_28327# a_13459_28111# 0.89fF
C3049 a_1858_25615# a_14839_20871# 0.35fF
C3050 a_9411_2215# nmat.col[1] 0.39fF
C3051 a_31214_57134# ctopp 3.57fF
C3052 VDD a_29455_31293# 0.77fF
C3053 pmat.row_n[14] pmat.row_n[3] 10.48fF
C3054 a_30210_71190# ctopp 3.40fF
C3055 VDD a_40250_57134# 0.52fF
C3056 a_20170_20536# a_21174_20536# 0.97fF
C3057 VDD a_39246_71190# 0.55fF
C3058 VDD a_26194_58138# 0.52fF
C3059 a_10781_42869# a_24833_40719# 0.82fF
C3060 nmat.col_n[26] ctopn 2.03fF
C3061 a_19166_16520# a_19166_15516# 1.00fF
C3062 a_12447_16143# nmat.col_n[1] 0.36fF
C3063 m2_17932_15246# m2_17932_14242# 0.99fF
C3064 a_35230_71190# m2_35000_72014# 1.00fF
C3065 VDD m2_17932_61974# 1.00fF
C3066 _1154_.X a_13091_28327# 1.05fF
C3067 a_34226_55126# vcm 0.58fF
C3068 VDD a_10867_41271# 0.60fF
C3069 m2_18936_7214# m3_19068_7346# 2.79fF
C3070 a_18546_24550# a_40158_24958# 0.35fF
C3071 a_9441_20189# a_2835_13077# 0.85fF
C3072 pmat.col[31] vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.51fF
C3073 a_3247_6037# a_3413_6037# 0.58fF
C3074 VDD a_13259_41001# 0.57fF
C3075 a_22178_68178# a_22178_67174# 1.00fF
C3076 a_42258_61150# vcm 0.62fF
C3077 a_2389_45859# a_1769_14735# 0.31fF
C3078 ANTENNA_fanout52_A.DIODE ANTENNA__1190__A1.DIODE 1.27fF
C3079 pmat.rowon_n[9] pmat.rowoff_n[9] 20.80fF
C3080 a_18546_22542# a_37146_22950# 0.35fF
C3081 VDD a_44966_43255# 0.75fF
C3082 pmat.en_bit_n[2] a_11067_27239# 0.43fF
C3083 VDD a_12053_27497# 0.70fF
C3084 VDD m2_43032_54946# 0.62fF
C3085 _1192_.B1 a_38851_28327# 0.52fF
C3086 a_9135_60967# a_10147_29415# 0.33fF
C3087 a_36234_20536# vcm 0.65fF
C3088 pmat.row_n[1] a_18162_9492# 25.57fF
C3089 a_12345_39100# a_12513_39100# 0.64fF
C3090 a_5651_66975# a_6559_33767# 1.08fF
C3091 a_2727_58470# a_1586_63927# 1.56fF
C3092 a_10515_15055# a_8305_20871# 0.46fF
C3093 VDD a_27198_59142# 0.52fF
C3094 VDD a_36193_35805# 1.44fF
C3095 a_25681_28879# a_21365_27247# 0.53fF
C3096 VDD a_10190_60663# 1.38fF
C3097 a_48282_17524# vcm 0.65fF
C3098 a_18546_16518# a_23090_16926# 0.35fF
C3099 m2_24960_54946# vcm 0.42fF
C3100 a_18546_9490# a_18162_9492# 2.61fF
C3101 ANTENNA__1187__B1.DIODE a_32405_32463# 0.40fF
C3102 a_49286_8488# vcm 0.64fF
C3103 a_31675_47695# a_7109_29423# 0.48fF
C3104 a_18162_59182# vcm 6.95fF
C3105 a_6664_26159# nmat.col_n[13] 1.48fF
C3106 pmat.col_n[17] vcm 2.79fF
C3107 a_2007_25597# a_11603_28335# 0.47fF
C3108 VDD a_34553_42658# 1.07fF
C3109 a_1923_31743# a_4075_28335# 0.35fF
C3110 m2_31988_7214# m2_32992_7214# 0.96fF
C3111 pmat.rowon_n[8] comp_latch 0.46fF
C3112 a_12585_39355# ndecision_finish 0.97fF
C3113 a_1858_25615# a_14287_31599# 0.35fF
C3114 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[26] 0.94fF
C3115 m2_51064_69002# vcm 0.51fF
C3116 pmat.row_n[3] a_18546_11498# 0.35fF
C3117 a_18546_72236# a_19074_72194# 0.35fF
C3118 VDD nmat.col_n[17] 5.25fF
C3119 a_25190_15516# vcm 0.65fF
C3120 VDD a_2983_48071# 2.13fF
C3121 a_9583_10121# comp_latch 0.75fF
C3122 a_1586_50247# a_2163_55233# 0.40fF
C3123 a_22199_30287# nmat.col_n[9] 0.90fF
C3124 _1154_.X a_17139_30503# 0.44fF
C3125 a_29206_70186# a_29206_69182# 1.00fF
C3126 VDD a_9731_8439# 0.46fF
C3127 pmat.rowon_n[3] a_3659_39733# 0.37fF
C3128 VDD a_12237_36596# 1.99fF
C3129 a_44266_12504# vcm 0.65fF
C3130 a_49286_64162# ctopp 3.57fF
C3131 a_13641_23439# a_21365_27247# 1.03fF
C3132 a_5651_66975# a_8385_51727# 0.59fF
C3133 m2_51064_8218# vcm 0.50fF
C3134 VDD a_18162_63198# 2.73fF
C3135 a_21174_23548# ctopn 3.39fF
C3136 VDD a_27198_19532# 0.52fF
C3137 nmat.rowon_n[7] a_10239_14183# 1.24fF
C3138 a_23182_9492# ctopn 3.57fF
C3139 VDD m2_28976_72014# 0.98fF
C3140 a_22178_57134# a_22178_56130# 1.00fF
C3141 a_26194_19532# a_27198_19532# 0.97fF
C3142 a_21174_60146# vcm 0.62fF
C3143 VDD a_26194_10496# 0.52fF
C3144 VDD a_19689_39141# 1.20fF
C3145 a_39246_20536# ctopn 3.58fF
C3146 VDD a_21124_42919# 1.24fF
C3147 a_18162_19532# vcm 6.95fF
C3148 a_18546_58180# a_33130_58138# 0.35fF
C3149 a_25190_10496# a_26194_10496# 0.97fF
C3150 a_18546_10494# a_33130_10902# 0.35fF
C3151 _1194_.B1 _1184_.A2 3.75fF
C3152 a_2419_53351# a_4991_69831# 0.38fF
C3153 a_13275_48783# a_11067_30287# 1.30fF
C3154 VDD a_8175_12533# 0.43fF
C3155 a_33222_62154# ctopp 3.58fF
C3156 a_5173_9839# a_5579_12394# 0.93fF
C3157 VDD a_42258_62154# 0.52fF
C3158 a_27198_16520# vcm 0.65fF
C3159 a_11041_39860# a_10873_39605# 3.94fF
C3160 a_11317_40188# a_14773_43746# 3.13fF
C3161 pmat.col[22] vcm 5.88fF
C3162 a_36234_56130# a_37238_56130# 0.97fF
C3163 a_18162_13508# ctopn 1.49fF
C3164 nmat.col[18] nmat.col_n[19] 8.01fF
C3165 a_2149_45717# a_1586_50247# 0.74fF
C3166 VDD a_16837_42043# 1.07fF
C3167 VDD a_4379_13818# 0.88fF
C3168 VDD a_8175_63669# 0.45fF
C3169 a_7717_14735# ANTENNA__1183__B1.DIODE 0.32fF
C3170 a_6743_31061# a_6909_31061# 0.59fF
C3171 a_19166_15516# m2_17932_15246# 0.96fF
C3172 a_21371_50087# nmat.col[15] 1.86fF
C3173 _1154_.A a_21371_50087# 1.08fF
C3174 a_32218_70186# ctopp 3.57fF
C3175 VDD a_41254_70186# 0.52fF
C3176 a_28202_15516# ctopn 3.58fF
C3177 VDD a_28202_11500# 0.52fF
C3178 pmat.rowoff_n[4] pmat.rowon_n[0] 1.10fF
C3179 VDD a_31015_29111# 0.46fF
C3180 a_48282_16520# a_48282_15516# 1.00fF
C3181 a_41254_62154# a_42258_62154# 0.97fF
C3182 a_13459_28111# a_30571_50959# 0.94fF
C3183 a_39246_66170# a_40250_66170# 0.97fF
C3184 m2_49056_72014# m3_49188_72146# 2.79fF
C3185 a_47278_12504# ctopn 3.58fF
C3186 a_18546_69224# a_28110_69182# 0.35fF
C3187 VDD a_2007_25597# 13.49fF
C3188 a_11317_36924# a_11297_36091# 0.54fF
C3189 a_43262_56130# vcm 0.62fF
C3190 VDD a_33489_36603# 1.17fF
C3191 _1194_.B1 a_9411_2215# 0.35fF
C3192 a_7415_29397# comp_latch 3.49fF
C3193 a_32218_63158# a_33222_63158# 0.97fF
C3194 a_18546_63200# a_47186_63158# 0.35fF
C3195 a_12044_49641# a_11948_49783# 0.47fF
C3196 _1154_.X a_26891_28327# 1.26fF
C3197 a_25190_22544# vcm 0.65fF
C3198 a_23182_68178# ctopp 3.58fF
C3199 a_46274_66170# vcm 0.62fF
C3200 VDD a_32218_68178# 0.52fF
C3201 a_8443_20719# a_8197_20871# 0.66fF
C3202 nmat.col[6] ctopn 1.97fF
C3203 a_11711_50959# a_21371_50087# 1.07fF
C3204 nmat.col[21] nmat.col[28] 13.72fF
C3205 a_18546_20534# nmat.rowoff_n[3] 4.09fF
C3206 a_39246_63158# vcm 0.62fF
C3207 VDD a_13979_65087# 0.36fF
C3208 VDD a_19405_28853# 3.94fF
C3209 pmat.rowoff_n[12] a_9441_20189# 0.89fF
C3210 a_19584_52423# a_18823_50247# 0.40fF
C3211 pmat.col_n[22] _1187_.A2 0.31fF
C3212 pmat.en_bit_n[2] _1196_.B1 0.53fF
C3213 a_18546_20534# a_34134_20942# 0.35fF
C3214 a_30210_16520# ctopn 3.58fF
C3215 a_30111_47911# a_13643_29415# 0.96fF
C3216 ANTENNA__1395__B1.DIODE a_46229_37583# 0.59fF
C3217 a_20438_35431# a_10873_38517# 0.41fF
C3218 nmat.col[4] m2_22952_24282# 0.40fF
C3219 VDD pmat.col[25] 4.35fF
C3220 VDD a_4951_76983# 0.39fF
C3221 a_1899_35051# a_2411_33749# 1.17fF
C3222 pmat.row_n[7] cgen.dlycontrol4_in[2] 0.83fF
C3223 VDD a_14887_46377# 5.04fF
C3224 a_10515_13967# nmat.col[3] 0.41fF
C3225 pmat.row_n[15] a_18162_23548# 25.57fF
C3226 VDD a_37238_23548# 0.55fF
C3227 _1154_.A a_34705_51959# 0.34fF
C3228 _1154_.X _1184_.A2 2.60fF
C3229 m2_51064_22274# m2_51064_21270# 0.99fF
C3230 a_40250_70186# a_41254_70186# 0.97fF
C3231 VDD a_39246_9492# 0.52fF
C3232 VDD a_4043_59861# 0.43fF
C3233 a_27198_11500# a_28202_11500# 0.97fF
C3234 a_18546_11498# a_37146_11906# 0.35fF
C3235 a_2411_16101# a_5087_18543# 0.70fF
C3236 a_2411_43301# a_2389_45859# 0.93fF
C3237 VDD a_31469_40726# 1.51fF
C3238 a_29206_64162# a_29206_63158# 1.00fF
C3239 a_32218_10496# a_32218_9492# 1.00fF
C3240 a_10515_13967# a_19283_49783# 0.98fF
C3241 pmat.col[26] ctopp 1.97fF
C3242 a_44266_67174# vcm 0.62fF
C3243 a_29206_58138# a_29206_57134# 1.00fF
C3244 nmat.rowon_n[7] ctopn 1.40fF
C3245 a_33222_14512# vcm 0.65fF
C3246 VDD a_10593_15823# 0.80fF
C3247 a_10781_42364# a_10949_42364# 3.41fF
C3248 cgen.start_conv_in a_30523_41245# 0.55fF
C3249 a_32218_64162# vcm 0.62fF
C3250 a_11337_25071# a_4523_21276# 0.35fF
C3251 a_33222_60146# a_33222_59142# 1.00fF
C3252 pmat.row_n[15] nmat.sw 0.58fF
C3253 a_21174_18528# a_21174_17524# 1.00fF
C3254 VDD a_31339_31787# 3.01fF
C3255 VDD ANTENNA__1190__B1.DIODE 21.06fF
C3256 pmat.col_n[25] ctopp 2.02fF
C3257 VDD a_35230_13508# 0.52fF
C3258 a_28202_22544# ctopn 3.57fF
C3259 nmat.col[13] vcm 5.78fF
C3260 VDD a_33222_18528# 0.52fF
C3261 a_38242_63158# pmat.col[19] 0.31fF
C3262 a_21174_63158# a_21174_62154# 1.00fF
C3263 m2_48052_54946# vcm 0.42fF
C3264 a_37238_67174# a_38242_67174# 0.97fF
C3265 a_34226_66170# a_34226_65166# 1.00fF
C3266 a_27198_22544# a_27198_21540# 1.00fF
C3267 VDD a_44266_15516# 0.52fF
C3268 a_1586_50247# cgen.dlycontrol3_in[3] 0.55fF
C3269 a_26194_14512# a_27198_14512# 0.97fF
C3270 a_18546_14510# a_35138_14918# 0.35fF
C3271 a_4128_64391# a_6175_60039# 0.70fF
C3272 a_25190_64162# a_26194_64162# 0.97fF
C3273 a_18546_64204# a_33130_64162# 0.35fF
C3274 a_31214_68178# a_32218_68178# 0.97fF
C3275 VDD a_14365_22351# 3.22fF
C3276 pmat.rowon_n[15] a_18162_71230# 1.19fF
C3277 a_24591_28327# nmat.col_n[30] 0.65fF
C3278 nmat.rowoff_n[11] ctopn 0.60fF
C3279 a_25190_8488# m2_24960_7214# 1.00fF
C3280 a_18546_72236# a_28110_72194# 0.35fF
C3281 a_11067_30287# a_23933_32143# 0.33fF
C3282 a_3746_58487# cgen.dlycontrol3_in[3] 0.62fF
C3283 a_30819_40191# a_10781_42364# 0.61fF
C3284 a_17996_41831# a_12658_42895# 0.40fF
C3285 a_10781_42869# a_10873_40693# 1.07fF
C3286 a_35230_65166# vcm 0.62fF
C3287 a_42258_21540# vcm 0.65fF
C3288 a_1586_63927# a_3136_59459# 0.62fF
C3289 a_31214_60146# ctopp 3.58fF
C3290 pmat.rowoff_n[7] a_1781_9308# 2.33fF
C3291 ANTENNA__1190__A2.DIODE a_9528_20407# 0.45fF
C3292 VDD a_40250_60146# 0.52fF
C3293 a_12197_38306# a_11921_35286# 0.31fF
C3294 _1196_.B1 nmat.col[3] 7.28fF
C3295 a_2124_72123# a_2163_71997# 0.79fF
C3296 a_25839_49783# a_25802_48169# 1.13fF
C3297 VDD a_1591_52815# 0.79fF
C3298 nmat.col_n[27] vcm 2.80fF
C3299 ANTENNA__1395__A2.DIODE nmat.col_n[2] 0.31fF
C3300 m2_50060_54946# m3_50768_55078# 0.82fF
C3301 a_7840_27247# a_12053_27497# 0.56fF
C3302 pmat.row_n[11] a_18162_67214# 25.57fF
C3303 a_17139_30503# a_40837_46261# 0.51fF
C3304 a_18546_19530# a_46182_19938# 0.35fF
C3305 a_36234_14512# ctopn 3.58fF
C3306 a_18547_51565# a_19541_28879# 0.74fF
C3307 ANTENNA__1395__B1.DIODE a_6664_26159# 0.86fF
C3308 a_18546_12502# a_50198_12910# 0.35fF
C3309 a_12585_39355# cgen.dlycontrol1_in[4] 0.32fF
C3310 VDD a_3879_42997# 0.40fF
C3311 VDD a_46274_16520# 0.52fF
C3312 VDD a_7109_29423# 9.20fF
C3313 a_18546_59184# a_28110_59142# 0.35fF
C3314 a_27198_65166# a_27198_64162# 1.00fF
C3315 a_44774_40821# a_35312_31599# 0.58fF
C3316 VDD a_35230_55126# 0.58fF
C3317 a_24186_57134# ctopp 3.57fF
C3318 ANTENNA__1187__B1.DIODE nmat.col_n[24] 0.46fF
C3319 a_23182_71190# ctopp 3.40fF
C3320 VDD a_33222_57134# 0.52fF
C3321 a_49286_69182# vcm 0.62fF
C3322 VDD a_32218_71190# 0.55fF
C3323 VDD a_5363_12015# 0.58fF
C3324 a_36234_23548# a_37238_23548# 0.97fF
C3325 a_32865_30199# a_33011_29941# 0.31fF
C3326 pmat.rowoff_n[4] a_4075_31591# 2.31fF
C3327 a_38242_9492# a_39246_9492# 0.97fF
C3328 VDD a_23663_38825# 0.60fF
C3329 a_45270_12504# a_45270_11500# 1.00fF
C3330 VDD a_28116_37479# 1.42fF
C3331 a_2419_69455# a_2659_35015# 0.44fF
C3332 VDD a_39193_42043# 1.19fF
C3333 a_6664_26159# a_8568_26703# 0.63fF
C3334 m2_17932_11230# vcm 0.44fF
C3335 a_18546_55168# a_44174_55126# 0.35fF
C3336 a_18546_24550# a_33130_24958# 0.35fF
C3337 a_41949_30761# a_34204_27765# 0.44fF
C3338 a_44266_8488# m2_44036_7214# 1.00fF
C3339 a_11067_30287# a_1781_9308# 0.95fF
C3340 a_35230_61150# vcm 0.62fF
C3341 a_4075_50087# a_4991_69831# 0.54fF
C3342 a_18546_72236# a_51202_72194# 0.35fF
C3343 a_18546_22542# a_30118_22950# 0.35fF
C3344 a_45270_21540# ctopn 3.58fF
C3345 pmat.rowon_n[0] clk_dig 0.52fF
C3346 VDD cgen.dlycontrol4_in[5] 7.48fF
C3347 a_10949_43124# a_11021_42619# 1.06fF
C3348 a_29206_20536# vcm 0.65fF
C3349 a_28202_65166# a_29206_65166# 0.97fF
C3350 VDD a_44266_22544# 0.52fF
C3351 nmat.rowon_n[13] nmat.rowoff_n[13] 21.98fF
C3352 VDD a_51202_8894# 0.30fF
C3353 VDD a_20170_59142# 0.52fF
C3354 a_2199_13887# a_8399_6037# 0.60fF
C3355 a_35230_21540# a_36234_21540# 0.97fF
C3356 VDD pmat.col_n[18] 5.22fF
C3357 a_37820_30485# nmat.col[15] 1.70fF
C3358 a_49286_63158# ctopp 3.57fF
C3359 a_1586_50247# a_1987_45370# 0.69fF
C3360 a_41254_17524# vcm 0.65fF
C3361 nmat.col[24] vcm 7.99fF
C3362 _1183_.A2 nmat.col[15] 3.63fF
C3363 a_18546_56172# a_19074_56130# 0.35fF
C3364 _1154_.A _1183_.A2 0.99fF
C3365 ANTENNA__1183__B1.DIODE nmat.col[21] 5.09fF
C3366 m2_29980_24282# m2_30984_24282# 0.96fF
C3367 nmat.sw a_11041_39860# 1.53fF
C3368 a_36234_71190# a_36234_70186# 1.00fF
C3369 a_42258_8488# vcm 0.64fF
C3370 a_4719_30287# cgen.dlycontrol4_in[5] 0.31fF
C3371 m2_24960_7214# m2_25964_7214# 0.96fF
C3372 nmat.rowon_n[13] vcm 0.53fF
C3373 a_13641_23439# _0467_ 1.11fF
C3374 VDD a_46723_30485# 0.35fF
C3375 a_18162_24552# vcm 7.69fF
C3376 a_4399_51157# a_4128_46983# 0.50fF
C3377 VDD a_2124_69947# 0.65fF
C3378 a_18546_13506# a_51202_13914# 0.35fF
C3379 a_34226_13508# a_35230_13508# 0.97fF
C3380 VDD nmat.col_n[8] 5.16fF
C3381 a_3746_58487# a_6467_29415# 0.52fF
C3382 VDD a_10795_47893# 0.53fF
C3383 a_11041_38772# a_11681_35823# 0.48fF
C3384 a_50290_61150# a_50290_60146# 1.00fF
C3385 a_35244_32411# a_46130_34319# 0.55fF
C3386 a_18546_18526# a_47186_18934# 0.35fF
C3387 a_32218_18528# a_33222_18528# 0.97fF
C3388 VDD a_18162_66210# 2.73fF
C3389 cgen.dlycontrol2_in[0] a_12309_36483# 1.06fF
C3390 a_1591_36501# a_1757_36501# 0.53fF
C3391 pmat.rowon_n[0] vcm 0.90fF
C3392 a_37238_12504# vcm 0.65fF
C3393 a_42258_64162# ctopp 3.58fF
C3394 a_11711_50959# _1183_.A2 0.78fF
C3395 nmat.col[26] m2_45040_24282# 0.39fF
C3396 pmat.sample a_18823_50247# 0.66fF
C3397 nmat.rowoff_n[9] ctopn 0.60fF
C3398 a_9411_2215# nmat.col_n[7] 1.14fF
C3399 pmat.en_bit_n[0] a_18243_28327# 0.82fF
C3400 VDD a_18162_10496# 2.74fF
C3401 a_2007_25597# a_7840_27247# 0.35fF
C3402 ANTENNA__1184__B1.DIODE nmat.col[12] 0.88fF
C3403 ANTENNA__1197__A.DIODE a_28915_50959# 0.69fF
C3404 ANTENNA__1190__A1.DIODE a_17139_30503# 0.46fF
C3405 VDD a_12513_39100# 1.88fF
C3406 a_32218_20536# ctopn 3.58fF
C3407 a_10223_26703# _0467_ 0.45fF
C3408 a_43262_15516# a_44266_15516# 0.97fF
C3409 _1196_.B1 nmat.col_n[18] 1.17fF
C3410 cgen.start_conv_in a_18975_40871# 0.61fF
C3411 a_18546_58180# a_26102_58138# 0.35fF
C3412 a_42258_69182# a_43262_69182# 0.97fF
C3413 a_21174_69182# a_21174_68178# 1.00fF
C3414 nmat.col[1] a_20170_24552# 0.38fF
C3415 a_18546_10494# a_26102_10902# 0.35fF
C3416 VDD a_2163_56765# 0.49fF
C3417 a_29206_21540# a_29206_20536# 1.00fF
C3418 VDD a_2511_34319# 0.45fF
C3419 a_44266_17524# ctopn 3.58fF
C3420 VDD a_13884_71311# 0.44fF
C3421 a_26194_62154# ctopp 3.58fF
C3422 cgen.dlycontrol3_in[4] a_24833_34191# 0.36fF
C3423 VDD a_35230_62154# 0.52fF
C3424 VDD m2_51064_13238# 0.99fF
C3425 _1192_.A2 a_25695_28111# 0.64fF
C3426 m2_38012_24282# vcm 0.42fF
C3427 a_45270_8488# ctopn 3.40fF
C3428 VDD a_32411_49559# 0.32fF
C3429 a_18546_56172# a_48190_56130# 0.35fF
C3430 VDD a_47186_24958# 0.44fF
C3431 nmat.col_n[22] vcm 2.80fF
C3432 a_24407_31375# nmat.col[14] 0.56fF
C3433 a_45270_65166# ctopp 3.58fF
C3434 ANTENNA__1197__A.DIODE ANTENNA__1395__B1.DIODE 18.55fF
C3435 _1194_.A2 a_13459_28111# 0.97fF
C3436 a_9217_23983# a_8861_24527# 1.20fF
C3437 a_18546_55168# a_27106_55126# 0.35fF
C3438 nmat.col_n[28] nmat.col[28] 6.07fF
C3439 a_31675_47695# clk_ena 1.25fF
C3440 VDD a_19166_20536# 0.56fF
C3441 a_10239_14183# a_2952_25045# 2.04fF
C3442 a_25190_70186# ctopp 3.57fF
C3443 a_3339_59879# a_8031_76757# 0.96fF
C3444 a_21174_15516# ctopn 3.58fF
C3445 cgen.dlycontrol3_in[3] cgen.dlycontrol3_in[1] 1.01fF
C3446 VDD a_34226_70186# 0.52fF
C3447 VDD a_21174_11500# 0.52fF
C3448 a_40250_23548# a_40250_22544# 1.00fF
C3449 a_10949_43124# a_11021_43011# 0.35fF
C3450 cgen.dlycontrol4_in[3] a_2411_33749# 0.60fF
C3451 a_39246_60146# a_40250_60146# 0.97fF
C3452 a_19166_65166# a_20170_65166# 0.97fF
C3453 a_40250_12504# ctopn 3.58fF
C3454 _1154_.X nmat.col[24] 0.96fF
C3455 a_18546_69224# a_21082_69182# 0.35fF
C3456 a_2683_22089# a_4703_24527# 0.38fF
C3457 a_23182_11500# a_23182_10496# 1.00fF
C3458 a_36234_56130# vcm 0.62fF
C3459 VDD a_17996_36391# 0.94fF
C3460 VDD a_7026_24527# 2.79fF
C3461 a_7415_29397# nmat.col[0] 0.39fF
C3462 pmat.col[26] m2_45040_54946# 0.39fF
C3463 a_23821_35279# a_24937_36039# 0.45fF
C3464 a_18546_63200# a_40158_63158# 0.35fF
C3465 m2_30984_24282# m3_31116_24414# 2.79fF
C3466 a_47278_68178# a_47278_67174# 1.00fF
C3467 a_4351_55527# a_5462_62215# 1.51fF
C3468 a_28202_61150# a_29206_61150# 0.97fF
C3469 a_2835_13077# a_10791_14191# 0.70fF
C3470 a_39246_66170# vcm 0.62fF
C3471 a_2419_53351# a_4075_68583# 0.47fF
C3472 VDD a_25190_68178# 0.52fF
C3473 a_14195_7351# nmat.rowoff_n[1] 2.54fF
C3474 m2_49056_72014# m2_50060_72014# 0.96fF
C3475 a_11711_50959# a_11416_50363# 0.46fF
C3476 VDD a_23479_43447# 0.65fF
C3477 a_39321_42333# a_39079_40947# 0.39fF
C3478 a_32218_63158# vcm 0.62fF
C3479 VDD a_8197_64789# 0.66fF
C3480 VDD a_41237_28585# 0.71fF
C3481 VDD a_7533_19087# 0.47fF
C3482 ANTENNA_fanout52_A.DIODE cgen.enable_dlycontrol_in 0.37fF
C3483 VDD a_46182_55126# 0.42fF
C3484 a_8031_76757# a_6292_69831# 0.33fF
C3485 VDD nmat.col_n[21] 14.98fF
C3486 a_22178_20536# a_23182_20536# 0.97fF
C3487 a_18546_20534# a_27106_20942# 0.35fF
C3488 VDD a_37823_34191# 0.35fF
C3489 a_23182_16520# ctopn 3.58fF
C3490 ANTENNA__1190__A1.DIODE a_26891_28327# 1.60fF
C3491 a_12053_27497# nmat.col_n[2] 0.36fF
C3492 a_2263_43719# a_38391_47381# 0.64fF
C3493 a_45270_16520# a_46274_16520# 0.97fF
C3494 nmat.rowon_n[5] ctopn 1.40fF
C3495 a_35230_67174# a_35230_66170# 1.00fF
C3496 a_21174_9492# a_21174_8488# 1.00fF
C3497 a_4075_31591# clk_dig 1.32fF
C3498 a_9135_60967# a_3746_58487# 0.70fF
C3499 VDD a_30210_23548# 0.55fF
C3500 VDD a_18162_58178# 2.73fF
C3501 a_45270_61150# ctopp 3.58fF
C3502 VDD a_32218_9492# 0.52fF
C3503 a_18546_11498# a_30118_11906# 0.35fF
C3504 a_5403_67655# a_3923_68021# 0.55fF
C3505 VDD a_23939_41271# 0.63fF
C3506 a_8583_29199# a_19405_28853# 0.59fF
C3507 m2_23956_7214# m3_24088_7346# 2.79fF
C3508 a_45019_38645# a_43776_30287# 0.55fF
C3509 VDD a_48282_20536# 0.52fF
C3510 VDD a_19409_40719# 0.92fF
C3511 a_34226_17524# a_35230_17524# 0.97fF
C3512 a_32218_57134# a_33222_57134# 0.97fF
C3513 a_2791_57703# a_1586_50247# 0.50fF
C3514 pmat.rowon_n[7] a_6467_29415# 0.52fF
C3515 a_37238_20536# a_37238_19532# 1.00fF
C3516 a_37238_67174# vcm 0.62fF
C3517 a_31214_71190# a_32218_71190# 0.97fF
C3518 a_18546_71232# a_45178_71190# 0.35fF
C3519 pmat.row_n[7] a_2411_16101# 1.59fF
C3520 _1187_.A2 a_16311_28327# 0.36fF
C3521 ANTENNA__1190__A1.DIODE _1184_.A2 2.96fF
C3522 a_37820_30485# a_37291_29397# 0.32fF
C3523 a_26194_14512# vcm 0.65fF
C3524 a_10239_14183# a_2683_22089# 0.66fF
C3525 nmat.rowon_n[6] nmat.rowoff_n[8] 0.55fF
C3526 VDD inn_analog 7.72fF
C3527 a_25190_64162# vcm 0.62fF
C3528 VDD m2_51064_54946# 1.20fF
C3529 a_35230_8488# a_36234_8488# 0.97fF
C3530 a_18546_65208# a_50198_65166# 0.35fF
C3531 cgen.dlycontrol4_in[1] a_2283_39189# 0.40fF
C3532 a_2411_33749# a_1591_33775# 0.34fF
C3533 VDD a_28202_13508# 0.52fF
C3534 a_24747_29967# nmat.col[30] 1.65fF
C3535 a_43262_14512# a_43262_13508# 1.00fF
C3536 pmat.rowon_n[7] a_13091_52047# 0.82fF
C3537 a_21174_22544# ctopn 3.57fF
C3538 VDD a_26194_18528# 0.52fF
C3539 a_18546_67216# a_50198_67174# 0.35fF
C3540 a_47278_57134# a_47278_56130# 1.00fF
C3541 pmat.rowon_n[8] a_2263_43719# 1.69fF
C3542 pmat.rowoff_n[12] a_5363_33551# 0.91fF
C3543 a_26194_19532# a_26194_18528# 1.00fF
C3544 VDD a_2944_67752# 0.48fF
C3545 m2_51064_71010# m2_51064_70006# 0.99fF
C3546 pmat.col_n[20] vcm 2.80fF
C3547 nmat.col_n[12] m2_30984_24282# 0.37fF
C3548 VDD a_37238_15516# 0.52fF
C3549 pmat.row_n[0] a_13643_29415# 0.85fF
C3550 a_18546_14510# a_28110_14918# 0.35fF
C3551 pmat.sw ANTENNA__1197__B.DIODE 1.64fF
C3552 a_18546_7482# a_50198_7890# 0.35fF
C3553 a_18546_64204# a_26102_64162# 0.35fF
C3554 a_13459_28111# a_32687_46607# 1.43fF
C3555 a_20170_24552# vcm 0.62fF
C3556 a_11057_35836# cgen.dlycontrol1_in[3] 0.46fF
C3557 a_4705_39759# cgen.dlycontrol2_in[2] 0.49fF
C3558 a_3866_57399# a_5497_62839# 0.59fF
C3559 VDD nmat.col[26] 9.13fF
C3560 VDD m2_41024_7214# 0.91fF
C3561 ANTENNA__1190__A1.DIODE a_9411_2215# 1.46fF
C3562 cgen.dlycontrol3_in[0] a_10767_39087# 0.43fF
C3563 a_2648_29397# a_4337_22351# 0.83fF
C3564 a_28202_65166# vcm 0.62fF
C3565 pmat.row_n[10] nmat.rowon_n[5] 20.68fF
C3566 a_35230_21540# vcm 0.65fF
C3567 a_24186_60146# ctopp 3.58fF
C3568 VDD a_33222_60146# 0.52fF
C3569 a_27794_28879# a_21365_27247# 0.38fF
C3570 VDD a_14773_37218# 2.05fF
C3571 VDD pmat.col_n[0] 5.43fF
C3572 a_13641_23439# nmat.col[12] 1.62fF
C3573 a_50290_58138# vcm 0.62fF
C3574 pmat.col[24] vcm 5.88fF
C3575 a_24186_17524# a_24186_16520# 1.00fF
C3576 pmat.sw a_24374_29941# 0.55fF
C3577 m2_41024_54946# m3_41156_55078# 2.79fF
C3578 a_19166_61150# a_20170_61150# 0.97fF
C3579 ANTENNA__1195__A1.DIODE a_21739_29415# 5.12fF
C3580 a_18546_19530# a_39154_19938# 0.35fF
C3581 m2_25964_54946# m2_26968_54946# 0.96fF
C3582 a_29206_14512# ctopn 3.58fF
C3583 pmat.en_bit_n[2] pmat.col[12] 0.37fF
C3584 a_30210_12504# a_31214_12504# 0.97fF
C3585 a_18546_12502# a_43170_12910# 0.35fF
C3586 VDD a_29864_39429# 1.15fF
C3587 a_43262_22544# a_44266_22544# 0.97fF
C3588 VDD a_32035_44265# 0.67fF
C3589 VDD a_39246_16520# 0.52fF
C3590 pmat.col[6] m2_24960_54946# 0.40fF
C3591 pmat.row_n[11] a_6821_18543# 0.39fF
C3592 m2_51064_10226# m2_51064_9222# 0.99fF
C3593 VDD a_12263_50959# 8.78fF
C3594 a_18546_59184# a_21082_59142# 0.35fF
C3595 pmat.row_n[12] ctopn 1.65fF
C3596 VDD a_29114_55126# 0.42fF
C3597 VDD a_49194_7890# 0.33fF
C3598 ANTENNA__1196__A2.DIODE nmat.col[15] 0.69fF
C3599 a_20170_24552# m3_20072_24702# 2.44fF
C3600 VDD a_26194_57134# 0.52fF
C3601 VDD a_27687_34967# 0.69fF
C3602 a_42258_69182# vcm 0.62fF
C3603 nmat.col[15] a_44697_48783# 0.74fF
C3604 VDD a_25190_71190# 0.55fF
C3605 a_18546_23546# a_48190_23954# 0.35fF
C3606 VDD a_21923_47919# 0.40fF
C3607 VDD a_14335_23439# 0.60fF
C3608 a_18546_67216# ctopp 1.59fF
C3609 a_10814_29111# a_5351_19913# 0.61fF
C3610 VDD a_28613_40229# 1.41fF
C3611 pmat.col[16] ctopp 2.03fF
C3612 ANTENNA__1183__B1.DIODE nmat.col_n[28] 5.05fF
C3613 VDD a_6403_37252# 0.61fF
C3614 a_1586_33927# a_4792_34435# 0.60fF
C3615 a_18546_55168# a_37146_55126# 0.35fF
C3616 a_18546_24550# a_26102_24958# 0.35fF
C3617 a_13091_52047# a_24602_48169# 0.66fF
C3618 a_5363_70543# a_9213_53903# 0.90fF
C3619 a_20605_40719# a_14712_37429# 0.60fF
C3620 a_46274_56130# ctopp 3.40fF
C3621 VDD a_5955_55223# 0.35fF
C3622 a_19166_67174# vcm 0.61fF
C3623 a_28202_61150# vcm 0.62fF
C3624 pmat.rowon_n[7] a_9135_60967# 5.28fF
C3625 pmat.row_n[9] pmat.rowoff_n[9] 0.32fF
C3626 a_18546_22542# a_23090_22950# 0.35fF
C3627 a_38242_21540# ctopn 3.58fF
C3628 VDD a_44635_46025# 0.33fF
C3629 a_11041_39860# a_20572_40517# 0.68fF
C3630 a_2407_49289# a_5779_71285# 1.68fF
C3631 a_11067_16359# a_7644_16341# 1.03fF
C3632 pmat.rowon_n[2] pmat.rowoff_n[2] 20.63fF
C3633 a_4707_32156# a_5179_31591# 0.69fF
C3634 VDD a_29711_47679# 0.53fF
C3635 a_22178_20536# vcm 0.65fF
C3636 VDD a_37238_22544# 0.52fF
C3637 a_49286_66170# ctopp 3.57fF
C3638 a_4068_25615# a_6579_29199# 0.35fF
C3639 a_11317_36924# a_11681_35823# 0.32fF
C3640 a_10873_36341# a_11113_36483# 0.33fF
C3641 a_42258_63158# ctopp 3.58fF
C3642 VDD m2_17932_16250# 1.11fF
C3643 a_11113_38659# cgen.dlycontrol2_in[1] 0.98fF
C3644 a_22186_30485# a_23352_30761# 0.36fF
C3645 a_34226_17524# vcm 0.65fF
C3646 a_3351_27249# a_2564_21959# 0.38fF
C3647 a_11202_55687# a_13091_54447# 0.40fF
C3648 a_6956_8965# a_6872_8725# 0.61fF
C3649 a_18546_61192# a_50198_61150# 0.35fF
C3650 nmat.col[13] m2_31988_24282# 0.39fF
C3651 nmat.en_bit_n[1] _1183_.A2 4.14fF
C3652 VDD config_2_in[8] 0.78fF
C3653 m2_22952_24282# m2_23956_24282# 0.96fF
C3654 a_35230_8488# vcm 0.64fF
C3655 a_20170_55126# m2_20944_54946# 0.96fF
C3656 a_1781_9308# a_18597_31599# 2.96fF
C3657 a_4259_73807# a_1923_61759# 0.40fF
C3658 a_3615_71631# a_5462_62215# 0.48fF
C3659 m2_17932_7214# m2_18936_7214# 0.96fF
C3660 VDD pmat.rowon_n[9] 3.51fF
C3661 _1192_.B1 a_12061_26703# 3.18fF
C3662 _1224_.X _1192_.A2 1.12fF
C3663 a_18243_28327# nmat.col_n[24] 0.31fF
C3664 VDD nmat.col_n[10] 7.27fF
C3665 a_46274_18528# a_46274_17524# 1.00fF
C3666 pmat.rowon_n[13] pmat.rowoff_n[13] 20.94fF
C3667 a_25755_34343# a_20534_35431# 1.24fF
C3668 a_50290_10496# vcm 0.65fF
C3669 VDD clk_ena 25.77fF
C3670 a_18546_13506# a_44174_13914# 0.35fF
C3671 nmat.rowoff_n[6] a_5899_21807# 0.32fF
C3672 a_46274_63158# a_46274_62154# 1.00fF
C3673 VDD a_29300_48463# 0.39fF
C3674 a_47278_67174# ctopp 3.58fF
C3675 a_4128_64391# a_7109_29423# 0.43fF
C3676 a_18546_18526# a_40158_18934# 0.35fF
C3677 a_7521_47081# a_4259_31375# 0.86fF
C3678 a_22178_70186# a_22178_69182# 1.00fF
C3679 VDD a_3207_65845# 0.45fF
C3680 VDD a_24015_36911# 0.62fF
C3681 a_10055_31591# a_9963_28111# 0.35fF
C3682 nmat.rowon_n[7] a_3746_58487# 2.09fF
C3683 pmat.en_bit_n[0] a_15667_28111# 1.13fF
C3684 a_30210_12504# vcm 0.65fF
C3685 a_35230_64162# ctopp 3.58fF
C3686 VDD a_45270_14512# 0.52fF
C3687 a_11067_64015# _1224_.X 0.57fF
C3688 VDD a_44266_64162# 0.52fF
C3689 a_18546_19530# a_21082_19938# 0.35fF
C3690 a_41731_49525# a_43659_28853# 0.56fF
C3691 VDD a_32371_50247# 0.38fF
C3692 a_45270_13508# a_45270_12504# 1.00fF
C3693 a_25190_20536# ctopn 3.58fF
C3694 a_5687_71829# a_2879_57487# 0.34fF
C3695 pmat.row_n[12] pmat.rowon_n[12] 20.09fF
C3696 pmat.col_n[28] ctopp 2.02fF
C3697 VDD a_20534_35431# 1.18fF
C3698 a_37238_17524# ctopn 3.58fF
C3699 a_41731_49525# a_33423_47695# 0.40fF
C3700 a_1923_61759# a_8695_63937# 0.36fF
C3701 pmat.row_n[15] pmat.rowoff_n[4] 0.88fF
C3702 VDD a_28202_62154# 0.52fF
C3703 a_19166_58138# a_19166_57134# 1.00fF
C3704 a_38242_8488# ctopn 3.40fF
C3705 a_12693_38543# a_12513_36924# 0.51fF
C3706 a_29206_56130# a_30210_56130# 0.97fF
C3707 a_18546_56172# a_41162_56130# 0.35fF
C3708 VDD a_40158_24958# 0.44fF
C3709 nmat.col_n[9] vcm 2.80fF
C3710 VDD pmat.rowon_n[11] 20.62fF
C3711 VDD pmat.rowon_n[5] 3.82fF
C3712 a_2879_57487# a_4583_68021# 0.54fF
C3713 pmat.rowon_n[8] a_10055_31591# 0.54fF
C3714 a_38242_65166# ctopp 3.58fF
C3715 VDD a_18272_42693# 1.04fF
C3716 a_18777_51183# _1192_.A2 0.41fF
C3717 VDD a_47278_65166# 0.52fF
C3718 _1154_.X a_25879_31591# 0.82fF
C3719 a_12116_39783# a_13909_39605# 0.62fF
C3720 a_1858_25615# nmat.col_n[12] 1.70fF
C3721 a_1923_31743# a_2163_31741# 0.58fF
C3722 a_18546_68220# a_49194_68178# 0.35fF
C3723 VDD a_23043_28335# 0.89fF
C3724 VDD a_27198_70186# 0.52fF
C3725 a_18546_72236# a_31122_72194# 0.35fF
C3726 a_20170_21540# ctopn 3.57fF
C3727 VDD a_4697_74005# 0.70fF
C3728 a_41254_16520# a_41254_15516# 1.00fF
C3729 a_34226_62154# a_35230_62154# 0.97fF
C3730 ANTENNA__1197__A.DIODE _1192_.B1 3.26fF
C3731 ANTENNA__1395__A1.DIODE nmat.en_bit_n[1] 0.50fF
C3732 _1196_.B1 a_15667_27239# 0.48fF
C3733 a_32218_66170# a_33222_66170# 0.97fF
C3734 VDD a_19166_22544# 0.56fF
C3735 cgen.dlycontrol3_in[4] a_1739_47893# 0.89fF
C3736 a_33222_12504# ctopn 3.58fF
C3737 a_7026_24527# a_4523_21276# 0.58fF
C3738 a_19166_11500# a_19166_10496# 1.00fF
C3739 a_29206_56130# vcm 0.62fF
C3740 a_18162_70226# vcm 6.95fF
C3741 VDD a_13158_71285# 0.92fF
C3742 nmat.col[18] m2_37008_24282# 0.40fF
C3743 a_4351_55527# a_4985_51433# 1.47fF
C3744 cgen.dlycontrol4_in[5] cgen.dlycontrol4_in[4] 10.00fF
C3745 a_18546_63200# a_33130_63158# 0.35fF
C3746 a_25190_63158# a_26194_63158# 0.97fF
C3747 ANTENNA__1197__A.DIODE a_23395_53135# 1.80fF
C3748 _1184_.A2 a_8305_20871# 0.47fF
C3749 a_32218_66170# vcm 0.62fF
C3750 a_4979_38127# a_5221_45199# 0.91fF
C3751 nmat.col[29] nmat.col_n[26] 3.06fF
C3752 a_13327_70741# pmat.row_n[13] 0.34fF
C3753 m2_42028_72014# m2_43032_72014# 0.96fF
C3754 a_14641_57711# a_10515_61839# 0.31fF
C3755 pmat.row_n[6] a_11435_58791# 0.55fF
C3756 a_19166_57134# m2_17932_56954# 0.96fF
C3757 a_25190_63158# vcm 0.62fF
C3758 VDD a_5495_65479# 0.58fF
C3759 a_23933_32143# a_24861_29673# 1.19fF
C3760 pmat.col_n[1] a_20170_55126# 0.31fF
C3761 VDD a_39154_55126# 0.42fF
C3762 VDD a_24160_30199# 0.63fF
C3763 a_7779_22583# a_7693_22365# 0.66fF
C3764 a_18546_20534# a_19074_20942# 0.35fF
C3765 VDD a_11271_73085# 0.52fF
C3766 nmat.rowon_n[14] cgen.dlycontrol4_in[2] 1.31fF
C3767 VDD a_23182_23548# 0.55fF
C3768 VDD a_36561_38780# 1.25fF
C3769 a_38242_61150# ctopp 3.58fF
C3770 a_33222_70186# a_34226_70186# 0.97fF
C3771 VDD a_25190_9492# 0.52fF
C3772 VDD a_47278_61150# 0.52fF
C3773 a_18546_11498# a_23090_11906# 0.35fF
C3774 VDD a_37776_37479# 1.35fF
C3775 a_1586_50247# a_1769_13103# 0.49fF
C3776 a_5779_71285# a_6568_59887# 0.36fF
C3777 a_34226_24552# ctopn 1.01fF
C3778 VDD a_41254_20536# 0.52fF
C3779 a_22178_64162# a_22178_63158# 1.00fF
C3780 VDD a_1895_38842# 0.49fF
C3781 a_17139_30503# a_44628_45717# 0.34fF
C3782 a_1923_31743# a_7619_30485# 0.81fF
C3783 a_25190_10496# a_25190_9492# 1.00fF
C3784 VDD pmat.sw 18.11fF
C3785 m2_17932_56954# m2_17932_55950# 0.99fF
C3786 a_18546_71232# a_38150_71190# 0.35fF
C3787 a_30210_67174# vcm 0.62fF
C3788 nmat.sw a_5266_17143# 0.60fF
C3789 a_22178_58138# a_22178_57134# 1.00fF
C3790 nmat.rowon_n[14] a_18162_9492# 1.33fF
C3791 a_35244_32411# nmat.col_n[31] 0.35fF
C3792 a_18162_14512# vcm 6.95fF
C3793 VDD a_1895_15994# 0.51fF
C3794 a_10239_14183# ANTENNA__1190__A2.DIODE 0.49fF
C3795 VDD a_13139_54599# 0.43fF
C3796 a_18546_8486# a_46182_8894# 0.35fF
C3797 a_26194_60146# a_26194_59142# 1.00fF
C3798 a_18546_65208# a_43170_65166# 0.35fF
C3799 VDD a_40567_32403# 0.35fF
C3800 nmat.col[1] a_9441_20189# 0.45fF
C3801 VDD a_26552_36165# 1.08fF
C3802 VDD pmat.col_n[21] 5.20fF
C3803 a_19166_17524# ctopn 3.43fF
C3804 a_44266_62154# a_44266_61150# 1.00fF
C3805 VDD a_21174_13508# 0.52fF
C3806 pmat.rowon_n[7] a_14653_53458# 0.77fF
C3807 a_19166_61150# m2_17932_60970# 0.96fF
C3808 cgen.dlycontrol4_in[3] a_36854_44527# 0.49fF
C3809 a_27789_44743# a_28245_44581# 0.48fF
C3810 VDD a_18162_18528# 2.74fF
C3811 a_18546_16518# a_18162_16520# 2.61fF
C3812 m2_17932_54946# vcm 0.42fF
C3813 a_20170_8488# ctopn 3.39fF
C3814 pmat.en_bit_n[0] _1194_.A2 0.41fF
C3815 a_30210_67174# a_31214_67174# 0.97fF
C3816 a_18546_67216# a_43170_67174# 0.35fF
C3817 a_4339_27804# nmat.col_n[13] 0.46fF
C3818 pmat.rowoff_n[7] cgen.dlycontrol3_in[2] 0.63fF
C3819 m2_17932_24282# m2_17932_23278# 0.99fF
C3820 a_27198_66170# a_27198_65166# 1.00fF
C3821 VDD a_23663_43177# 0.60fF
C3822 VDD a_30210_15516# 0.52fF
C3823 a_44266_15516# a_44266_14512# 1.00fF
C3824 cgen.dlycontrol3_in[4] cgen.dlycontrol4_in[0] 0.83fF
C3825 a_39939_29967# a_38913_31055# 0.43fF
C3826 pmat.col_n[26] pmat.col[27] 5.87fF
C3827 a_18546_7482# a_43170_7890# 0.35fF
C3828 a_46274_69182# a_46274_68178# 1.00fF
C3829 a_24186_68178# a_25190_68178# 0.97fF
C3830 VDD a_27001_30511# 0.65fF
C3831 a_2046_30184# cgen.dlycontrol1_in[0] 0.66fF
C3832 a_33957_48437# a_35186_47375# 0.43fF
C3833 VDD a_49286_12504# 0.52fF
C3834 VDD m2_26968_7214# 1.27fF
C3835 a_2603_22357# a_2769_22357# 0.75fF
C3836 VDD a_4871_17429# 0.47fF
C3837 cgen.dlycontrol4_in[2] a_11021_43011# 2.13fF
C3838 a_10781_42869# a_10781_42364# 4.11fF
C3839 a_22199_30287# nmat.col_n[18] 0.54fF
C3840 VDD a_10697_75218# 2.85fF
C3841 a_21174_65166# vcm 0.62fF
C3842 a_28202_21540# vcm 0.65fF
C3843 pmat.col_n[16] a_24867_53135# 0.93fF
C3844 pmat.rowoff_n[11] ctopp 0.60fF
C3845 VDD a_26194_60146# 0.52fF
C3846 ANTENNA__1184__B1.DIODE a_28915_50959# 0.66fF
C3847 a_24591_28327# pmat.col[10] 0.65fF
C3848 a_43262_58138# vcm 0.62fF
C3849 _1179_.X vcm 0.82fF
C3850 a_18546_19530# a_32126_19938# 0.35fF
C3851 a_22178_14512# ctopn 3.58fF
C3852 a_18546_12502# a_36142_12910# 0.35fF
C3853 VDD a_19873_44219# 1.23fF
C3854 VDD a_32218_16520# 0.52fF
C3855 a_6451_67655# a_13183_72405# 0.50fF
C3856 a_36345_42567# a_36801_42405# 0.39fF
C3857 VDD a_2389_45859# 3.69fF
C3858 a_20170_65166# a_20170_64162# 1.00fF
C3859 VDD a_22086_55126# 0.42fF
C3860 VDD a_42166_7890# 0.33fF
C3861 VDD a_12447_16143# 11.64fF
C3862 a_48282_11500# a_48282_10496# 1.00fF
C3863 _1179_.X _1194_.B1 0.80fF
C3864 ANTENNA__1197__B.DIODE a_13459_28111# 0.32fF
C3865 nmat.en_bit_n[1] ANTENNA__1196__A2.DIODE 0.34fF
C3866 a_24867_53135# ANTENNA__1195__A1.DIODE 0.67fF
C3867 ANTENNA__1184__B1.DIODE ANTENNA__1395__B1.DIODE 0.82fF
C3868 ANTENNA__1395__A1.DIODE a_19584_52423# 0.51fF
C3869 a_35230_69182# vcm 0.62fF
C3870 a_44774_48695# a_43315_48437# 0.36fF
C3871 a_30571_50959# a_40951_31599# 0.76fF
C3872 _1194_.B1 a_33423_47695# 2.13fF
C3873 a_29206_23548# a_30210_23548# 0.97fF
C3874 a_18546_23546# a_41162_23954# 0.35fF
C3875 a_18823_50247# a_21371_50087# 0.50fF
C3876 a_16083_50069# a_10883_3303# 0.38fF
C3877 a_5357_62779# a_6175_60039# 0.45fF
C3878 a_21174_71190# m2_20944_72014# 1.00fF
C3879 a_31214_9492# a_32218_9492# 0.97fF
C3880 a_18546_9490# a_45178_9898# 0.35fF
C3881 VDD a_5558_9527# 1.40fF
C3882 a_44266_59142# vcm 0.62fF
C3883 VDD a_5687_38279# 0.94fF
C3884 a_38242_12504# a_38242_11500# 1.00fF
C3885 a_11207_11079# a_9675_10396# 0.33fF
C3886 _1154_.X a_24591_28327# 1.99fF
C3887 _1187_.A2 a_24407_31375# 0.31fF
C3888 a_39246_56130# ctopp 3.40fF
C3889 VDD a_39127_29423# 0.67fF
C3890 a_6292_65479# a_7099_74313# 1.24fF
C3891 pmat.col[3] ctopp 1.97fF
C3892 VDD a_48282_56130# 0.55fF
C3893 nmat.rowon_n[1] nmat.rowon_n[6] 0.53fF
C3894 a_47278_20536# a_48282_20536# 0.97fF
C3895 a_18546_71232# a_20078_71190# 0.35fF
C3896 a_33839_46805# a_35186_47375# 0.50fF
C3897 a_21174_61150# vcm 0.62fF
C3898 a_31214_21540# ctopn 3.58fF
C3899 ANTENNA__1190__B1.DIODE nmat.col[15] 4.43fF
C3900 VDD a_20267_47375# 0.58fF
C3901 a_25879_31591# a_40837_46261# 0.32fF
C3902 a_46274_9492# a_46274_8488# 1.00fF
C3903 a_21174_65166# a_22178_65166# 0.97fF
C3904 VDD a_30210_22544# 0.52fF
C3905 a_42258_66170# ctopp 3.58fF
C3906 a_4719_30287# a_5687_38279# 0.62fF
C3907 a_10515_15055# a_9463_50877# 0.34fF
C3908 VDD a_5341_59317# 0.33fF
C3909 a_16890_36911# a_15049_36374# 0.75fF
C3910 a_6283_31591# clk_dig 0.67fF
C3911 a_28202_21540# a_29206_21540# 0.97fF
C3912 a_35230_63158# ctopp 3.58fF
C3913 VDD a_44266_63158# 0.52fF
C3914 a_27198_17524# vcm 0.65fF
C3915 a_1586_8439# a_1757_15829# 0.38fF
C3916 m2_37008_24282# m3_37140_24414# 2.79fF
C3917 nmat.col[7] nmat.rowoff_n[14] 1.51fF
C3918 a_2952_25045# a_7779_22583# 0.32fF
C3919 nmat.col_n[18] nmat.col_n[30] 0.87fF
C3920 a_18546_61192# a_43170_61150# 0.35fF
C3921 a_10055_31591# a_8907_48437# 0.30fF
C3922 m2_49056_54946# m2_50060_54946# 0.93fF
C3923 a_29206_71190# a_29206_70186# 1.00fF
C3924 a_28202_8488# vcm 0.64fF
C3925 a_17139_30503# a_22628_30485# 0.40fF
C3926 pmat.row_n[15] vcm 1.14fF
C3927 a_43262_58138# a_44266_58138# 0.97fF
C3928 a_18546_19530# ctopn 1.59fF
C3929 VDD a_31095_42367# 0.60fF
C3930 m2_17932_14242# m3_18064_14374# 2.76fF
C3931 VDD a_17748_29673# 0.47fF
C3932 a_44266_19532# vcm 0.65fF
C3933 VDD a_18546_21538# 32.65fF
C3934 ANTENNA_fanout52_A.DIODE ANTENNA__1395__B1.DIODE 0.71fF
C3935 a_11067_30287# a_30999_48071# 0.38fF
C3936 a_43262_10496# vcm 0.65fF
C3937 a_27198_13508# a_28202_13508# 0.97fF
C3938 a_18546_13506# a_37146_13914# 0.35fF
C3939 a_10699_72943# a_9279_71829# 0.35fF
C3940 cgen.start_conv_in a_10873_38517# 2.07fF
C3941 a_11149_40188# a_24833_40719# 0.48fF
C3942 a_40250_71190# m2_40020_72014# 1.00fF
C3943 pmat.row_n[4] nmat.sw 1.37fF
C3944 VDD a_28629_48437# 0.30fF
C3945 pmat.col[0] vcm 5.85fF
C3946 a_43262_61150# a_43262_60146# 1.00fF
C3947 a_2124_65595# a_2163_65469# 0.58fF
C3948 a_40250_67174# ctopp 3.58fF
C3949 _1154_.X _1179_.X 4.00fF
C3950 a_25190_18528# a_26194_18528# 0.97fF
C3951 a_18546_18526# a_33130_18934# 0.35fF
C3952 _1196_.B1 a_11067_27239# 0.45fF
C3953 VDD a_49286_67174# 0.52fF
C3954 a_3571_13627# comp_latch 0.65fF
C3955 VDD a_12513_36924# 1.37fF
C3956 a_20438_35431# cgen.dlycontrol1_in[2] 1.66fF
C3957 a_23182_12504# vcm 0.65fF
C3958 a_28202_64162# ctopp 3.58fF
C3959 VDD a_39387_41271# 0.60fF
C3960 VDD a_38242_14512# 0.52fF
C3961 ANTENNA__1195__A1.DIODE a_38851_28327# 0.34fF
C3962 a_16311_28327# a_25695_28111# 0.50fF
C3963 m2_28976_7214# m3_29108_7346# 2.79fF
C3964 VDD a_37238_64162# 0.52fF
C3965 pmat.col[3] m2_21948_54946# 0.40fF
C3966 VDD a_32035_39913# 0.68fF
C3967 a_8583_29199# clk_ena 0.58fF
C3968 a_18546_57176# a_51202_57134# 0.35fF
C3969 a_16311_28327# a_1781_9308# 5.38fF
C3970 pmat.row_n[12] ctopp 1.65fF
C3971 a_1769_13103# cgen.dlycontrol3_in[1] 0.33fF
C3972 a_44266_59142# a_44266_58138# 1.00fF
C3973 a_4075_50087# a_7436_58487# 0.30fF
C3974 cgen.dlycontrol3_in[2] nmat.rowon_n[14] 1.90fF
C3975 a_9411_2215# nmat.col[12] 0.65fF
C3976 VDD a_8481_10396# 1.56fF
C3977 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top ANTENNA__1190__A2.DIODE 0.38fF
C3978 VDD config_1_in[10] 0.79fF
C3979 VDD a_16745_44581# 1.17fF
C3980 cgen.dlycontrol4_in[2] a_3325_40847# 1.15fF
C3981 a_18546_21538# nmat.rowoff_n[2] 4.09fF
C3982 a_18546_18526# nmat.rowoff_n[5] 4.09fF
C3983 a_36234_15516# a_37238_15516# 0.97fF
C3984 VDD m2_24960_24282# 0.62fF
C3985 a_19439_32149# a_19605_32149# 0.58fF
C3986 a_1899_35051# cgen.dlycontrol3_in[4] 0.95fF
C3987 pmat.row_n[9] pmat.row_n[6] 9.53fF
C3988 a_19166_18528# a_19166_17524# 1.00fF
C3989 VDD nmat.col_n[14] 5.23fF
C3990 a_19166_11500# ctopn 3.43fF
C3991 a_35230_69182# a_36234_69182# 0.97fF
C3992 a_22178_21540# a_22178_20536# 1.00fF
C3993 VDD a_5989_34863# 0.63fF
C3994 a_33467_46261# a_30111_47911# 1.59fF
C3995 a_30210_17524# ctopn 3.58fF
C3996 a_45270_11500# vcm 0.65fF
C3997 pmat.col[5] ctopp 1.97fF
C3998 VDD a_21174_62154# 0.52fF
C3999 a_20170_23548# a_21174_23548# 0.97fF
C4000 cgen.dlycontrol4_in[3] a_14773_43746# 4.45fF
C4001 a_49286_17524# a_49286_16520# 1.00fF
C4002 a_31214_8488# ctopn 3.40fF
C4003 cgen.dlycontrol3_in[3] a_10767_39087# 1.30fF
C4004 a_18546_56172# a_34134_56130# 0.35fF
C4005 VDD a_33130_24958# 0.44fF
C4006 a_24747_29967# nmat.col[28] 1.96fF
C4007 m2_46044_24282# m2_47048_24282# 0.96fF
C4008 VDD a_11142_64783# 0.44fF
C4009 VDD a_11435_58791# 13.53fF
C4010 pmat.col_n[23] vcm 2.80fF
C4011 a_12069_38517# a_11681_35823# 4.10fF
C4012 a_47278_19532# ctopn 3.58fF
C4013 a_31214_65166# ctopp 3.58fF
C4014 a_2683_22089# a_7779_22583# 0.83fF
C4015 pmat.row_n[11] a_18162_19532# 25.57fF
C4016 a_50290_57134# m2_51064_56954# 0.96fF
C4017 pmat.rowon_n[3] nmat.rowoff_n[14] 0.30fF
C4018 m2_17932_11230# m3_18064_11362# 2.76fF
C4019 VDD a_40250_65166# 0.52fF
C4020 a_13091_52047# a_13275_48783# 0.63fF
C4021 nmat.col_n[1] ctopn 2.01fF
C4022 VDD a_47278_21540# 0.52fF
C4023 pmat.row_n[2] pmat.rowoff_n[3] 1.84fF
C4024 a_44266_59142# a_45270_59142# 0.97fF
C4025 a_46274_10496# ctopn 3.58fF
C4026 pmat.col[0] pmat.col[10] 0.38fF
C4027 a_32218_62154# pmat.col[13] 0.31fF
C4028 a_18546_68220# a_42166_68178# 0.35fF
C4029 a_3615_71631# a_1674_57711# 0.34fF
C4030 a_49286_68178# vcm 0.62fF
C4031 VDD a_20170_70186# 0.52fF
C4032 a_33222_23548# a_33222_22544# 1.00fF
C4033 a_24833_40719# a_30543_40721# 0.36fF
C4034 a_6787_47607# a_11115_71285# 0.71fF
C4035 VDD a_14071_74879# 0.39fF
C4036 m2_17932_13238# m2_17932_12234# 0.99fF
C4037 VDD m2_17932_57958# 1.00fF
C4038 a_32218_60146# a_33222_60146# 0.97fF
C4039 a_18546_60188# a_47186_60146# 0.35fF
C4040 a_11435_58791# a_4719_30287# 0.41fF
C4041 m2_20944_72014# m3_21076_72146# 2.79fF
C4042 a_26194_12504# ctopn 3.58fF
C4043 ANTENNA__1190__A1.DIODE a_25879_31591# 3.27fF
C4044 a_22178_56130# vcm 0.62fF
C4045 a_10515_13967# _1196_.B1 0.37fF
C4046 VDD a_22537_36911# 3.65fF
C4047 nmat.col[7] vcm 5.76fF
C4048 nmat.col[17] vcm 5.76fF
C4049 a_18563_27791# a_28336_29967# 0.53fF
C4050 nmat.col[18] nmat.col[19] 3.29fF
C4051 a_18546_63200# a_26102_63158# 0.35fF
C4052 m2_46044_54946# m3_46176_55078# 2.79fF
C4053 VDD m2_44036_72014# 1.11fF
C4054 a_40250_68178# a_40250_67174# 1.00fF
C4055 pmat.col[31] ANTENNA__1190__B1.DIODE 0.80fF
C4056 a_21174_61150# a_22178_61150# 0.97fF
C4057 a_45270_69182# ctopp 3.58fF
C4058 nmat.sample_n vcm 1.22fF
C4059 a_25190_66170# vcm 0.62fF
C4060 VDD a_10991_68591# 0.64fF
C4061 a_19166_22544# m2_18936_23278# 0.99fF
C4062 m2_35000_72014# m2_36004_72014# 0.96fF
C4063 VDD a_34887_39095# 0.63fF
C4064 pmat.rowoff_n[7] a_2263_43719# 0.82fF
C4065 VDD a_44791_43541# 0.51fF
C4066 a_48282_11500# ctopn 3.58fF
C4067 ANTENNA_fanout52_A.DIODE a_30111_47911# 0.57fF
C4068 _1154_.X pmat.col[0] 1.03fF
C4069 pmat.rowoff_n[4] a_5363_33551# 1.72fF
C4070 pmat.rowon_n[3] clk_dig 1.25fF
C4071 a_50290_61150# m2_51064_60970# 0.96fF
C4072 a_14457_15823# nmat.rowoff_n[11] 0.94fF
C4073 a_38242_16520# a_39246_16520# 0.97fF
C4074 VDD a_45450_48695# 0.57fF
C4075 a_28202_67174# a_28202_66170# 1.00fF
C4076 VDD a_7048_23277# 0.96fF
C4077 VDD a_16377_38779# 1.13fF
C4078 a_31214_61150# ctopp 3.58fF
C4079 nmat.col[12] nmat.col[13] 6.53fF
C4080 a_10814_29111# a_9075_28023# 0.36fF
C4081 a_2411_43301# a_1591_50095# 0.33fF
C4082 VDD a_40250_61150# 0.52fF
C4083 VDD a_40628_39429# 1.76fF
C4084 VDD a_29217_41570# 1.46fF
C4085 VDD a_20170_14512# 0.52fF
C4086 a_13641_23439# a_8568_26703# 0.53fF
C4087 m2_17932_8218# m3_18064_8350# 2.76fF
C4088 VDD a_19166_64162# 0.58fF
C4089 a_5351_19913# a_2683_22089# 0.46fF
C4090 nmat.rowon_n[7] a_4259_31375# 0.58fF
C4091 a_50290_18528# vcm 0.65fF
C4092 VDD a_34226_20536# 0.52fF
C4093 a_27198_17524# a_28202_17524# 0.97fF
C4094 pmat.sw a_4523_21276# 0.37fF
C4095 m2_51064_64986# vcm 0.51fF
C4096 a_25190_57134# a_26194_57134# 0.97fF
C4097 cgen.dlycontrol1_in[2] cgen.dlycontrol1_in[0] 0.81fF
C4098 cgen.dlycontrol4_in[1] a_2835_13077# 0.38fF
C4099 a_30210_20536# a_30210_19532# 1.00fF
C4100 a_24186_71190# a_25190_71190# 0.97fF
C4101 a_18546_71232# a_31122_71190# 0.35fF
C4102 a_23182_67174# vcm 0.62fF
C4103 a_7658_71543# a_6787_47607# 0.83fF
C4104 nmat.rowoff_n[6] nmat.rowon_n[6] 20.79fF
C4105 m3_20072_55078# ctopp 0.35fF
C4106 a_2648_29397# clk_dig 1.03fF
C4107 a_5363_70543# a_10190_60663# 0.58fF
C4108 nmat.rowon_n[14] a_6872_8725# 0.58fF
C4109 VDD a_46274_17524# 0.52fF
C4110 VDD a_5331_28309# 0.41fF
C4111 VDD m2_20944_54946# 0.61fF
C4112 a_28202_8488# a_29206_8488# 0.97fF
C4113 a_18546_8486# a_39154_8894# 0.35fF
C4114 a_18546_65208# a_36142_65166# 0.35fF
C4115 a_47278_70186# a_47278_69182# 1.00fF
C4116 VDD a_47278_8488# 0.55fF
C4117 nmat.col_n[6] vcm 2.80fF
C4118 a_2199_13887# a_3247_6037# 0.68fF
C4119 a_18546_21538# a_50198_21946# 0.35fF
C4120 VDD a_5131_13255# 0.34fF
C4121 a_36234_14512# a_36234_13508# 1.00fF
C4122 VDD a_7212_62607# 0.36fF
C4123 a_29455_31293# a_30603_29575# 0.56fF
C4124 a_2263_43719# a_11067_30287# 1.08fF
C4125 a_18546_67216# a_36142_67174# 0.35fF
C4126 a_40250_57134# a_40250_56130# 1.00fF
C4127 _1194_.A2 cgen.dlycontrol1_in[0] 0.45fF
C4128 a_44266_19532# a_45270_19532# 0.97fF
C4129 pmat.rowon_n[3] vcm 0.85fF
C4130 a_20170_12504# a_20170_11500# 1.00fF
C4131 VDD a_23182_15516# 0.52fF
C4132 nmat.col_n[3] nmat.col[3] 0.78fF
C4133 nmat.col[21] nmat.col_n[19] 5.25fF
C4134 ANTENNA__1184__B1.DIODE nmat.col[18] 0.95fF
C4135 a_7717_14735# nmat.en_bit_n[0] 0.55fF
C4136 ANTENNA__1195__A1.DIODE nmat.col_n[19] 2.14fF
C4137 a_18546_7482# a_36142_7890# 0.35fF
C4138 VDD a_15753_28879# 1.36fF
C4139 a_43262_10496# a_44266_10496# 0.97fF
C4140 pmat.col_n[30] pmat.col_n[31] 1.19fF
C4141 ANTENNA__1187__B1.DIODE nmat.col[29] 1.37fF
C4142 VDD a_42258_12504# 0.52fF
C4143 a_8491_47911# pmat.row_n[15] 0.33fF
C4144 VDD a_13459_28111# 20.48fF
C4145 m2_17932_19262# vcm 0.44fF
C4146 a_21174_21540# vcm 0.65fF
C4147 VDD a_5267_65479# 0.37fF
C4148 a_50290_57134# vcm 0.62fF
C4149 VDD a_36617_37691# 1.37fF
C4150 a_49286_71190# vcm 0.60fF
C4151 a_36234_58138# vcm 0.62fF
C4152 a_41254_56130# m2_41024_54946# 0.99fF
C4153 a_3387_22869# a_2835_13077# 0.44fF
C4154 a_12228_39605# a_15049_36374# 0.91fF
C4155 a_6568_59887# a_4025_54965# 0.46fF
C4156 a_10245_51335# a_9427_50095# 0.59fF
C4157 a_18546_19530# a_25098_19938# 0.35fF
C4158 a_33423_47695# a_40837_46261# 1.41fF
C4159 a_24407_31375# a_13275_48783# 0.34fF
C4160 VDD a_12044_49641# 0.89fF
C4161 a_23182_12504# a_24186_12504# 0.97fF
C4162 a_18546_12502# a_29114_12910# 0.35fF
C4163 a_36234_22544# a_37238_22544# 0.97fF
C4164 VDD a_25190_16520# 0.52fF
C4165 a_3983_41941# a_4149_41941# 0.41fF
C4166 VDD m2_48052_24282# 0.62fF
C4167 VDD a_6829_26703# 2.63fF
C4168 VDD a_35138_7890# 0.34fF
C4169 pmat.col_n[31] ctopp 1.92fF
C4170 VDD a_12341_57141# 0.66fF
C4171 a_28202_69182# vcm 0.62fF
C4172 a_6787_47607# a_11797_60431# 0.85fF
C4173 a_18546_23546# a_34134_23954# 0.35fF
C4174 a_28336_29967# a_39496_30199# 0.36fF
C4175 nmat.rowon_n[7] a_2564_21959# 2.96fF
C4176 a_15667_27239# a_22199_30287# 0.88fF
C4177 a_41731_49525# a_43776_30287# 0.31fF
C4178 a_37820_30485# a_35244_32411# 0.97fF
C4179 m2_29980_24282# vcm 0.42fF
C4180 cgen.dlycontrol3_in[2] a_3325_40847# 0.35fF
C4181 a_18546_9490# a_38150_9898# 0.35fF
C4182 ANTENNA__1190__A2.DIODE a_82736_4943# 0.32fF
C4183 pmat.rowoff_n[2] vcm 0.33fF
C4184 a_37238_59142# vcm 0.62fF
C4185 a_18563_27791# nmat.col_n[18] 0.38fF
C4186 ANTENNA__1184__B1.DIODE _1192_.B1 0.35fF
C4187 pmat.row_n[0] a_14379_6567# 1.26fF
C4188 a_7717_14735# a_37612_30663# 0.30fF
C4189 a_18546_24550# ctopn 0.38fF
C4190 a_23821_35279# a_28116_37479# 0.31fF
C4191 a_18546_17522# a_18162_17524# 2.61fF
C4192 VDD a_14471_4943# 0.39fF
C4193 a_2407_49289# a_4399_51157# 0.91fF
C4194 a_32218_56130# ctopp 3.40fF
C4195 a_7435_68021# a_5307_67655# 0.30fF
C4196 VDD a_41254_56130# 0.55fF
C4197 a_3615_71631# a_12067_67279# 0.31fF
C4198 a_30210_8488# m2_29980_7214# 1.00fF
C4199 a_9963_13967# ANTENNA__1196__A2.DIODE 0.56fF
C4200 a_18546_72236# a_34134_72194# 0.35fF
C4201 VDD a_8013_25615# 1.27fF
C4202 a_24186_21540# ctopn 3.58fF
C4203 a_2263_43719# nmat.rowon_n[14] 0.47fF
C4204 _1224_.X a_16311_28327# 0.71fF
C4205 a_1586_33927# a_3983_41941# 0.73fF
C4206 ANTENNA__1190__A1.DIODE a_24591_28327# 1.88fF
C4207 _1187_.A2 ANTENNA__1187__B1.DIODE 11.90fF
C4208 a_13091_28327# a_28915_50959# 0.35fF
C4209 a_18546_66212# a_51202_66170# 0.35fF
C4210 a_18546_8486# a_21082_8894# 0.35fF
C4211 VDD a_23182_22544# 0.52fF
C4212 a_35230_66170# ctopp 3.58fF
C4213 VDD a_9231_32117# 0.39fF
C4214 VDD a_44266_66170# 0.52fF
C4215 a_45270_11500# a_46274_11500# 0.97fF
C4216 VDD a_12309_36483# 2.60fF
C4217 a_9183_72007# a_9279_71829# 0.37fF
C4218 VDD pmat.col_n[1] 7.26fF
C4219 a_28202_63158# ctopp 3.58fF
C4220 VDD a_37238_63158# 0.52fF
C4221 a_47278_64162# a_47278_63158# 1.00fF
C4222 a_50290_10496# a_50290_9492# 1.00fF
C4223 a_18546_61192# a_36142_61150# 0.35fF
C4224 VDD a_9528_20407# 4.02fF
C4225 nmat.col_n[12] nmat.col[1] 10.19fF
C4226 m2_42028_54946# m2_43032_54946# 0.96fF
C4227 a_21174_8488# vcm 0.64fF
C4228 _1194_.A2 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top 0.92fF
C4229 a_47278_58138# a_47278_57134# 1.00fF
C4230 VDD a_19233_41479# 1.50fF
C4231 pmat.row_n[1] a_13643_29415# 4.76fF
C4232 nmat.col[3] nmat.rowoff_n[14] 0.45fF
C4233 VDD pmat.row_n[9] 22.23fF
C4234 cgen.dlycontrol3_in[4] cgen.dlycontrol4_in[3] 0.33fF
C4235 VDD m2_51064_21270# 1.13fF
C4236 pmat.sample_n a_13459_28111# 2.89fF
C4237 a_37238_19532# vcm 0.65fF
C4238 a_13091_28327# ANTENNA__1395__B1.DIODE 0.64fF
C4239 a_39246_18528# a_39246_17524# 1.00fF
C4240 a_35244_32411# a_34204_27765# 0.39fF
C4241 a_1923_61759# a_3727_66113# 0.36fF
C4242 a_9411_2215# nmat.col_n[13] 1.80fF
C4243 VDD a_34002_34191# 0.47fF
C4244 a_36234_10496# vcm 0.65fF
C4245 a_18546_13506# a_30118_13914# 0.35fF
C4246 VDD a_6451_67655# 7.85fF
C4247 pmat.col_n[29] pmat.col[29] 1.14fF
C4248 a_5363_33551# clk_dig 1.53fF
C4249 nmat.col[23] ctopn 1.97fF
C4250 a_39246_63158# a_39246_62154# 1.00fF
C4251 a_33222_67174# ctopp 3.58fF
C4252 VDD vcm.sky130_fd_sc_hd__buf_4_2.A 0.41fF
C4253 a_18546_18526# a_26102_18934# 0.35fF
C4254 VDD a_42258_67174# 0.52fF
C4255 VDD a_11921_37462# 1.52fF
C4256 a_45270_22544# a_45270_21540# 1.00fF
C4257 a_21174_64162# ctopp 3.58fF
C4258 VDD a_13985_41317# 1.31fF
C4259 VDD a_31214_14512# 0.52fF
C4260 a_44266_14512# a_45270_14512# 0.97fF
C4261 VDD a_30210_64162# 0.52fF
C4262 a_13479_26935# a_12851_28853# 0.42fF
C4263 a_18546_17522# a_48190_17930# 0.35fF
C4264 a_43262_64162# a_44266_64162# 0.97fF
C4265 a_49286_68178# a_50290_68178# 0.97fF
C4266 pmat.rowoff_n[12] nmat.rowoff_n[3] 20.42fF
C4267 a_18546_57176# a_44174_57134# 0.35fF
C4268 VDD pmat.rowon_n[13] 3.80fF
C4269 a_49286_8488# m2_49056_7214# 1.00fF
C4270 _1179_.X ANTENNA__1190__A1.DIODE 0.40fF
C4271 a_40250_23548# m2_40020_24282# 0.99fF
C4272 a_38242_13508# a_38242_12504# 1.00fF
C4273 a_13275_48783# a_17842_27497# 0.33fF
C4274 pmat.en_bit_n[0] ANTENNA__1197__B.DIODE 3.25fF
C4275 a_18546_15514# a_48190_15922# 0.35fF
C4276 a_32687_46607# a_40951_31599# 1.77fF
C4277 VDD m2_44036_54946# 0.62fF
C4278 a_17139_30503# a_28915_50959# 0.68fF
C4279 a_18546_59184# ctopp 1.59fF
C4280 a_11435_58791# a_10595_53361# 0.37fF
C4281 VDD a_34887_35831# 0.63fF
C4282 a_23182_17524# ctopn 3.58fF
C4283 VDD pmat.col_n[24] 5.38fF
C4284 a_38242_11500# vcm 0.65fF
C4285 a_25190_63158# pmat.col[6] 0.31fF
C4286 VDD a_2944_61493# 0.66fF
C4287 a_11317_36924# ndecision_finish 0.53fF
C4288 nmat.col_n[7] nmat.col[7] 0.78fF
C4289 m2_25964_54946# vcm 0.42fF
C4290 a_24186_8488# ctopn 3.40fF
C4291 a_18546_56172# a_27106_56130# 0.35fF
C4292 a_22178_56130# a_23182_56130# 0.97fF
C4293 a_13432_62581# a_11007_58229# 0.78fF
C4294 VDD a_26102_24958# 0.44fF
C4295 m2_39016_24282# m2_40020_24282# 0.96fF
C4296 a_19166_59142# vcm 0.61fF
C4297 a_25575_31055# nmat.col[29] 0.49fF
C4298 nmat.col_n[22] m2_41024_24282# 0.37fF
C4299 a_4257_34319# cgen.dlycontrol1_in[2] 0.40fF
C4300 a_40250_19532# ctopn 3.58fF
C4301 a_24186_65166# ctopp 3.58fF
C4302 VDD a_34611_43177# 0.63fF
C4303 VDD a_33222_65166# 0.52fF
C4304 ANTENNA__1395__B1.DIODE a_13145_26935# 0.69fF
C4305 VDD a_40250_21540# 0.52fF
C4306 a_45270_65166# a_45270_64162# 1.00fF
C4307 m2_17932_67998# vcm 0.44fF
C4308 a_39246_10496# ctopn 3.58fF
C4309 a_18546_68220# a_35138_68178# 0.35fF
C4310 a_2411_16101# a_3571_13627# 0.64fF
C4311 a_46274_58138# ctopp 3.58fF
C4312 a_42258_68178# vcm 0.62fF
C4313 VDD a_11487_69653# 0.68fF
C4314 a_1957_43567# a_4075_31591# 0.77fF
C4315 VDD a_2129_10383# 0.52fF
C4316 VDD nmat.col[22] 4.36fF
C4317 VDD a_6883_51335# 0.40fF
C4318 VDD a_4259_73807# 5.89fF
C4319 a_27198_62154# a_28202_62154# 0.97fF
C4320 a_34226_16520# a_34226_15516# 1.00fF
C4321 a_6835_51183# pmat.rowon_n[3] 0.48fF
C4322 VDD a_19541_28879# 7.36fF
C4323 a_25190_66170# a_26194_66170# 0.97fF
C4324 a_18546_60188# a_40158_60146# 0.35fF
C4325 a_18162_12504# ctopn 1.49fF
C4326 VDD a_46912_34319# 0.44fF
C4327 a_8305_20871# a_7644_16341# 0.98fF
C4328 VDD a_13837_36893# 1.40fF
C4329 VDD a_19166_63158# 0.56fF
C4330 pmat.en_bit_n[2] a_22186_30485# 0.55fF
C4331 VDD m2_29980_72014# 1.00fF
C4332 nmat.col_n[13] nmat.col[13] 0.85fF
C4333 a_41731_49525# a_44774_40821# 0.42fF
C4334 a_47278_23548# vcm 0.65fF
C4335 a_38242_69182# ctopp 3.58fF
C4336 a_49286_9492# vcm 0.65fF
C4337 VDD a_47278_69182# 0.52fF
C4338 nmat.col[3] vcm 5.76fF
C4339 m2_27972_72014# m2_28976_72014# 0.96fF
C4340 a_11948_49783# a_35186_47375# 0.43fF
C4341 VDD a_18235_39095# 0.63fF
C4342 a_45270_63158# pmat.col[26] 0.31fF
C4343 VDD a_23571_44265# 0.64fF
C4344 VDD a_9335_51727# 0.77fF
C4345 a_19166_19532# vcm 0.65fF
C4346 _1196_.B1 a_13091_7655# 0.31fF
C4347 a_46274_65166# a_47278_65166# 0.97fF
C4348 a_47278_59142# ctopp 3.58fF
C4349 a_41254_11500# ctopn 3.58fF
C4350 VDD a_7999_31359# 0.47fF
C4351 a_33309_36039# a_33765_35877# 0.39fF
C4352 VDD a_8695_12801# 0.48fF
C4353 cgen.dlycontrol3_in[4] a_11297_36091# 0.80fF
C4354 a_28915_50959# a_26891_28327# 2.37fF
C4355 VDD a_11113_38659# 0.62fF
C4356 a_24186_61150# ctopp 3.58fF
C4357 a_19166_13508# ctopn 3.43fF
C4358 nmat.col_n[12] vcm 2.80fF
C4359 a_26194_70186# a_27198_70186# 0.97fF
C4360 VDD a_33222_61150# 0.52fF
C4361 a_24407_31375# a_1781_9308# 1.47fF
C4362 VDD a_16111_40183# 0.58fF
C4363 a_37291_29397# inn_analog 0.36fF
C4364 a_45270_13508# vcm 0.65fF
C4365 VDD a_8695_63937# 0.52fF
C4366 a_5351_19913# ANTENNA__1190__A2.DIODE 0.41fF
C4367 nmat.col_n[28] nmat.col_n[19] 11.18fF
C4368 a_43262_18528# vcm 0.65fF
C4369 VDD a_27198_20536# 0.52fF
C4370 pmat.col[11] vcm 5.88fF
C4371 VDD dummypin[15] 0.78fF
C4372 a_1586_18231# a_7809_17705# 0.34fF
C4373 a_18546_71232# a_24094_71190# 0.35fF
C4374 a_4128_64391# a_11435_58791# 1.05fF
C4375 a_18546_22542# a_19074_22950# 0.35fF
C4376 a_14149_39747# a_13503_39069# 0.38fF
C4377 VDD a_39246_17524# 0.52fF
C4378 pmat.col_n[14] pmat.col[14] 0.76fF
C4379 VDD a_33775_29111# 0.43fF
C4380 a_18546_20534# vcm 0.40fF
C4381 a_18546_8486# a_32126_8894# 0.35fF
C4382 a_18546_65208# a_29114_65166# 0.35fF
C4383 a_10515_15055# a_13091_18535# 0.33fF
C4384 VDD a_23455_32447# 0.34fF
C4385 VDD a_40250_8488# 0.55fF
C4386 a_18546_21538# a_43170_21946# 0.35fF
C4387 a_37238_62154# a_37238_61150# 1.00fF
C4388 a_20170_11500# vcm 0.65fF
C4389 a_14365_22351# a_14691_29575# 0.41fF
C4390 a_10441_21263# a_4339_27804# 0.71fF
C4391 a_13641_23439# a_10441_21263# 0.34fF
C4392 a_50290_23548# ctopn 3.37fF
C4393 m2_42028_24282# m3_42160_24414# 2.79fF
C4394 VDD m2_51064_70006# 1.00fF
C4395 a_18546_67216# a_29114_67174# 0.35fF
C4396 a_23182_67174# a_24186_67174# 0.97fF
C4397 a_11067_27239# a_22199_30287# 4.28fF
C4398 a_50290_60146# vcm 0.62fF
C4399 a_7840_27247# a_6829_26703# 0.52fF
C4400 a_2199_13887# a_6956_8965# 0.52fF
C4401 pmat.rowoff_n[8] pmat.row_n[6] 1.71fF
C4402 a_20170_66170# a_20170_65166# 1.00fF
C4403 a_37238_15516# a_37238_14512# 1.00fF
C4404 VDD a_11203_62037# 0.59fF
C4405 a_18546_7482# a_29114_7890# 0.35fF
C4406 a_10055_31591# a_11067_64015# 2.28fF
C4407 ANTENNA__1395__B1.DIODE _1184_.A2 3.75fF
C4408 a_39246_69182# a_39246_68178# 1.00fF
C4409 VDD a_9899_30724# 0.43fF
C4410 a_47278_21540# a_47278_20536# 1.00fF
C4411 VDD a_35230_12504# 0.52fF
C4412 pmat.row_n[2] nmat.rowon_n[13] 20.76fF
C4413 VDD m2_51064_9222# 0.99fF
C4414 a_13479_26935# nmat.col_n[1] 0.39fF
C4415 VDD a_4429_76751# 0.59fF
C4416 pmat.rowon_n[6] a_18162_62194# 1.19fF
C4417 a_18546_62196# a_19074_62154# 0.35fF
C4418 _1192_.B1 nmat.col_n[29] 0.87fF
C4419 a_28915_50959# a_9411_2215# 0.64fF
C4420 a_48282_13508# ctopn 3.58fF
C4421 VDD a_5939_60137# 0.51fF
C4422 a_43262_57134# vcm 0.62fF
C4423 pmat.row_n[11] a_4075_31591# 1.47fF
C4424 a_42258_71190# vcm 0.60fF
C4425 pmat.rowoff_n[4] pmat.row_n[4] 20.93fF
C4426 a_46274_18528# ctopn 3.58fF
C4427 a_29206_58138# vcm 0.62fF
C4428 a_13459_28111# a_22499_49783# 1.84fF
C4429 m2_33996_7214# m3_34128_7346# 2.79fF
C4430 pmat.sample a_21124_42919# 0.50fF
C4431 nmat.en_bit_n[0] a_7415_29397# 0.84fF
C4432 VDD a_33047_41001# 0.63fF
C4433 VDD a_54136_39932# 0.36fF
C4434 ANTENNA__1197__A.DIODE a_7717_14735# 0.40fF
C4435 cgen.dlycontrol3_in[3] cgen.dlycontrol4_in[2] 2.29fF
C4436 a_5731_58951# a_5535_57993# 0.65fF
C4437 VDD a_11987_10089# 0.86fF
C4438 a_18546_12502# a_22086_12910# 0.35fF
C4439 cgen.dlycontrol2_in[4] a_12585_40443# 1.19fF
C4440 VDD m3_39148_7346# 0.38fF
C4441 VDD a_24937_43655# 2.07fF
C4442 a_11021_42619# a_10949_42364# 2.04fF
C4443 pmat.row_n[4] nmat.col_n[3] 0.42fF
C4444 nmat.rowoff_n[10] nmat.rowon_n[10] 20.94fF
C4445 VDD a_12079_9615# 6.42fF
C4446 a_31214_62154# pmat.col[12] 0.31fF
C4447 VDD a_33869_31599# 0.38fF
C4448 _1196_.B1 nmat.sw 0.58fF
C4449 VDD a_28110_7890# 0.33fF
C4450 a_12069_36341# a_15144_36165# 0.50fF
C4451 a_41254_11500# a_41254_10496# 1.00fF
C4452 a_11067_49871# a_19283_49783# 0.38fF
C4453 VDD a_14589_35286# 1.07fF
C4454 a_21174_69182# vcm 0.62fF
C4455 a_2727_58470# a_4509_62037# 0.42fF
C4456 a_4259_73807# a_1823_60949# 0.36fF
C4457 a_22178_23548# a_23182_23548# 0.97fF
C4458 a_18546_23546# a_27106_23954# 0.35fF
C4459 ANTENNA_fanout52_A.DIODE a_30663_50087# 0.50fF
C4460 nmat.col_n[18] vcm 3.48fF
C4461 m2_49056_54946# vcm 0.41fF
C4462 a_24186_9492# a_25190_9492# 0.97fF
C4463 a_18546_9490# a_31122_9898# 0.35fF
C4464 a_46274_61150# a_47278_61150# 0.97fF
C4465 VDD a_36234_24552# 0.58fF
C4466 a_11067_64015# a_13688_47893# 0.48fF
C4467 m2_50060_24282# m2_51064_24282# 0.59fF
C4468 pmat.col[31] clk_ena 16.07fF
C4469 a_30210_59142# vcm 0.62fF
C4470 a_31214_12504# a_31214_11500# 1.00fF
C4471 pmat.col_n[26] vcm 2.80fF
C4472 a_1591_40853# a_1757_40853# 0.46fF
C4473 pmat.rowon_n[7] a_2046_30184# 0.42fF
C4474 pmat.sw nmat.col[15] 0.92fF
C4475 a_1586_50247# a_1769_14735# 0.41fF
C4476 _1154_.A pmat.sw 15.24fF
C4477 a_9963_28111# a_6664_26159# 0.37fF
C4478 a_12345_39100# a_12197_38306# 2.10fF
C4479 a_21371_50087# a_37820_30485# 0.45fF
C4480 VDD a_6487_5629# 0.51fF
C4481 a_25190_56130# ctopp 3.40fF
C4482 a_6051_74183# a_5931_74183# 0.59fF
C4483 VDD a_34226_56130# 0.54fF
C4484 a_40250_20536# a_41254_20536# 0.97fF
C4485 _1194_.B1 nmat.col_n[18] 1.42fF
C4486 VDD a_4989_11079# 0.68fF
C4487 a_20170_13508# a_20170_12504# 1.00fF
C4488 VDD m3_24088_72146# 0.33fF
C4489 a_13275_48783# a_26479_32117# 0.41fF
C4490 a_11067_30287# a_25688_32117# 0.36fF
C4491 a_10515_15055# a_10883_3303# 1.01fF
C4492 pmat.col_n[10] a_13091_28327# 0.40fF
C4493 VDD a_1643_74005# 0.40fF
C4494 a_18546_62196# a_48190_62154# 0.35fF
C4495 a_18546_66212# a_44174_66170# 0.35fF
C4496 a_39246_9492# a_39246_8488# 1.00fF
C4497 a_28202_66170# ctopp 3.58fF
C4498 m2_25964_72014# m3_26096_72146# 2.79fF
C4499 VDD a_37238_66170# 0.52fF
C4500 a_32405_32463# a_44571_32143# 0.35fF
C4501 a_11149_36924# a_11225_35836# 4.87fF
C4502 a_21174_21540# a_22178_21540# 0.97fF
C4503 VDD a_30095_36919# 0.59fF
C4504 a_21174_63158# ctopp 3.58fF
C4505 nmat.col[9] m2_27972_24282# 0.41fF
C4506 VDD a_30210_63158# 0.52fF
C4507 nmat.col[8] nmat.col_n[8] 0.72fF
C4508 a_4523_21276# a_9528_20407# 0.47fF
C4509 a_2952_25045# a_2564_21959# 0.39fF
C4510 m2_51064_54946# m3_51196_55078# 2.79fF
C4511 a_18546_61192# a_29114_61150# 0.35fF
C4512 pmat.col[1] pmat.col[5] 0.44fF
C4513 a_22178_71190# a_22178_70186# 1.00fF
C4514 a_49286_71190# a_50290_71190# 0.97fF
C4515 a_28704_29568# nmat.col[29] 0.48fF
C4516 a_36234_58138# a_37238_58138# 0.97fF
C4517 a_13643_29415# a_9307_31068# 0.38fF
C4518 cgen.dlycontrol2_in[3] a_14149_39747# 1.29fF
C4519 a_5363_33551# a_11823_46973# 0.32fF
C4520 VDD a_46582_46519# 0.93fF
C4521 a_30210_19532# vcm 0.65fF
C4522 VDD pmat.en_bit_n[0] 11.33fF
C4523 VDD a_6559_6031# 1.06fF
C4524 VDD a_16745_34427# 1.13fF
C4525 a_29206_10496# vcm 0.65fF
C4526 a_18546_13506# a_23090_13914# 0.35fF
C4527 a_33395_43455# a_30819_40191# 0.41fF
C4528 comp.adc_nor_latch_0.R comp.adc_nor_latch_0.NOR_1/A 0.35fF
C4529 a_3339_59879# a_5535_57993# 0.60fF
C4530 a_36234_61150# a_36234_60146# 1.00fF
C4531 a_26194_67174# ctopp 3.58fF
C4532 a_44266_19532# a_44266_18528# 1.00fF
C4533 a_18546_70228# a_46182_70186# 0.35fF
C4534 VDD a_35230_67174# 0.52fF
C4535 a_10651_37683# a_11317_36924# 0.30fF
C4536 a_18546_11498# a_18162_11500# 2.61fF
C4537 VDD a_30913_38053# 1.29fF
C4538 m2_51064_69002# m2_51064_67998# 0.99fF
C4539 a_10781_42364# a_11297_36091# 0.53fF
C4540 a_17139_30503# nmat.col[18] 2.20fF
C4541 VDD a_32405_32463# 6.82fF
C4542 VDD a_24186_14512# 0.52fF
C4543 a_24186_56130# m2_23956_54946# 0.99fF
C4544 a_45270_62154# vcm 0.62fF
C4545 VDD a_23182_64162# 0.52fF
C4546 a_27763_27221# nmat.col[21] 0.40fF
C4547 a_18546_17522# a_41162_17930# 0.35fF
C4548 ANTENNA__1395__B1.DIODE nmat.col[13] 0.87fF
C4549 a_18546_57176# a_37146_57134# 0.35fF
C4550 a_37238_59142# a_37238_58138# 1.00fF
C4551 VDD a_3069_69367# 0.42fF
C4552 a_29163_38545# a_27603_34191# 0.41fF
C4553 m3_35132_55078# ctopp 0.31fF
C4554 a_23395_53135# a_13091_28327# 0.46fF
C4555 _1187_.A2 a_18243_28327# 2.87fF
C4556 a_3339_70759# a_5081_53135# 0.73fF
C4557 VDD a_44573_45173# 0.43fF
C4558 a_14839_20871# nmat.rowon_n[1] 0.72fF
C4559 a_29206_15516# a_30210_15516# 0.97fF
C4560 a_18546_15514# a_41162_15922# 0.35fF
C4561 a_6787_47607# a_4075_31591# 0.49fF
C4562 _1154_.X nmat.col_n[18] 0.59fF
C4563 a_28202_69182# a_29206_69182# 0.97fF
C4564 VDD a_33684_32143# 0.43fF
C4565 a_8305_20871# a_4976_16091# 0.61fF
C4566 VDD a_17113_35877# 1.22fF
C4567 a_30571_50959# a_45908_33749# 0.36fF
C4568 pmat.col_n[1] pmat.col_n[3] 0.56fF
C4569 a_44266_70186# vcm 0.62fF
C4570 a_31214_11500# vcm 0.65fF
C4571 a_13459_28111# nmat.col_n[2] 0.35fF
C4572 a_36234_24552# a_36234_23548# 1.00fF
C4573 nmat.rowoff_n[13] nmat.rowoff_n[10] 0.55fF
C4574 a_42258_17524# a_42258_16520# 1.00fF
C4575 nmat.sw a_10873_39605# 0.51fF
C4576 a_48282_12504# a_49286_12504# 0.97fF
C4577 a_18563_27791# a_21341_28585# 0.35fF
C4578 a_33222_19532# ctopn 3.58fF
C4579 a_2564_21959# a_2683_22089# 0.53fF
C4580 VDD a_26194_65166# 0.52fF
C4581 VDD a_33222_21540# 0.52fF
C4582 a_37238_59142# a_38242_59142# 0.97fF
C4583 pmat.rowon_n[0] a_18546_8486# 4.09fF
C4584 a_1923_31743# a_2007_25597# 1.19fF
C4585 a_32218_10496# ctopn 3.58fF
C4586 a_18546_68220# a_28110_68178# 0.35fF
C4587 a_39246_58138# ctopp 3.58fF
C4588 a_35230_68178# vcm 0.62fF
C4589 VDD a_48282_58138# 0.52fF
C4590 VDD nmat.col[11] 4.38fF
C4591 a_26194_23548# a_26194_22544# 1.00fF
C4592 VDD a_11508_48187# 0.31fF
C4593 a_18546_60188# a_33130_60146# 0.35fF
C4594 a_25190_60146# a_26194_60146# 0.97fF
C4595 pmat.col_n[12] ANTENNA__1395__A2.DIODE 0.32fF
C4596 a_16800_47213# a_13275_48783# 1.18fF
C4597 a_4075_68583# pmat.rowon_n[0] 1.03fF
C4598 VDD a_19166_66170# 0.56fF
C4599 a_2021_26677# a_2648_29397# 0.44fF
C4600 _1192_.B1 a_17139_30503# 0.88fF
C4601 a_13357_37429# a_15049_36374# 1.77fF
C4602 a_21981_34191# a_11057_35836# 0.97fF
C4603 a_19166_62154# a_19166_61150# 1.00fF
C4604 pmat.en_bit_n[2] a_21365_27247# 0.85fF
C4605 a_7415_29397# a_6664_26159# 0.67fF
C4606 a_20170_56130# a_20170_55126# 1.00fF
C4607 a_33222_68178# a_33222_67174# 1.00fF
C4608 a_40250_23548# vcm 0.65fF
C4609 a_31214_69182# ctopp 3.58fF
C4610 a_42258_9492# vcm 0.65fF
C4611 a_18546_14510# ctopn 1.59fF
C4612 VDD a_40250_69182# 0.52fF
C4613 VDD a_19166_10496# 0.56fF
C4614 VDD pmat.col[8] 5.38fF
C4615 a_1591_31599# cgen.dlycontrol3_in[0] 1.08fF
C4616 pmat.row_n[6] ctopn 1.65fF
C4617 m2_20944_72014# m2_21948_72014# 0.96fF
C4618 a_19541_28879# a_8583_29199# 0.52fF
C4619 VDD a_10985_44220# 1.16fF
C4620 a_3175_72641# a_3136_72515# 0.57fF
C4621 a_40837_46261# a_43776_30287# 0.37fF
C4622 nmat.en_bit_n[1] clk_ena 0.46fF
C4623 a_40250_59142# ctopp 3.58fF
C4624 VDD a_18162_55166# 27.52fF
C4625 a_34226_11500# ctopn 3.58fF
C4626 VDD a_49286_59142# 0.52fF
C4627 a_15667_27239# a_41731_49525# 1.18fF
C4628 ANTENNA__1395__A1.DIODE a_34705_51959# 1.07fF
C4629 cgen.dlycontrol3_in[2] cgen.dlycontrol3_in[3] 1.33fF
C4630 VDD a_4421_70741# 0.31fF
C4631 pmat.row_n[15] pmat.row_n[5] 1.35fF
C4632 VDD m2_17932_12234# 1.01fF
C4633 a_31214_16520# a_32218_16520# 0.97fF
C4634 a_18546_16518# a_45178_16926# 0.35fF
C4635 m2_39016_24282# vcm 0.42fF
C4636 a_21174_67174# a_21174_66170# 1.00fF
C4637 a_2411_43301# a_1586_50247# 1.24fF
C4638 pmat.rowoff_n[13] ctopp 0.60fF
C4639 nmat.col_n[25] vcm 2.80fF
C4640 pmat.rowoff_n[9] ctopp 0.60fF
C4641 VDD pmat.rowoff_n[8] 4.71fF
C4642 VDD a_26194_61150# 0.52fF
C4643 VDD a_11565_39061# 1.25fF
C4644 a_38242_13508# vcm 0.65fF
C4645 VDD a_31923_42367# 0.79fF
C4646 ANTENNA__1197__A.DIODE ANTENNA__1195__A1.DIODE 0.94fF
C4647 a_36234_18528# vcm 0.65fF
C4648 ANTENNA__1184__B1.DIODE a_10883_3303# 0.67fF
C4649 a_18546_57176# a_18162_57174# 2.62fF
C4650 a_23182_20536# a_23182_19532# 1.00fF
C4651 a_3339_59879# a_8197_76757# 0.64fF
C4652 pmat.row_n[4] vcm 1.15fF
C4653 a_23182_23548# m2_22952_24282# 0.99fF
C4654 a_18546_72236# a_37146_72194# 0.35fF
C4655 nmat.col[15] nmat.col_n[14] 6.59fF
C4656 VDD m3_51196_64114# 0.35fF
C4657 a_47278_15516# vcm 0.65fF
C4658 VDD a_32218_17524# 0.52fF
C4659 a_20170_15516# a_21174_15516# 0.97fF
C4660 VDD a_13830_47607# 0.54fF
C4661 pmat.rowon_n[0] a_3325_20175# 0.63fF
C4662 a_18546_8486# a_25098_8894# 0.35fF
C4663 a_21174_8488# a_22178_8488# 0.97fF
C4664 a_18546_65208# a_22086_65166# 0.35fF
C4665 a_40250_70186# a_40250_69182# 1.00fF
C4666 a_19166_69182# a_20170_69182# 0.97fF
C4667 VDD a_33222_8488# 0.55fF
C4668 a_14943_26703# nmat.col_n[3] 0.78fF
C4669 a_12934_35823# a_15049_36374# 0.37fF
C4670 a_18546_21538# a_36142_21946# 0.35fF
C4671 VDD a_19965_36603# 1.25fF
C4672 VDD a_23090_72194# 0.33fF
C4673 a_29206_14512# a_29206_13508# 1.00fF
C4674 a_10147_29415# a_19605_30511# 0.58fF
C4675 a_43262_23548# ctopn 3.40fF
C4676 VDD a_49286_19532# 0.52fF
C4677 pmat.rowon_n[11] nmat.en_bit_n[1] 1.10fF
C4678 a_45270_9492# ctopn 3.57fF
C4679 a_18546_67216# a_22086_67174# 0.35fF
C4680 a_33222_57134# a_33222_56130# 1.00fF
C4681 a_18546_22542# vcm 0.40fF
C4682 VDD a_4703_24527# 2.73fF
C4683 a_37238_19532# a_38242_19532# 0.97fF
C4684 a_11115_71285# a_5651_66975# 1.17fF
C4685 a_1923_61759# a_1674_57711# 0.56fF
C4686 a_12228_39605# ndecision_finish 1.89fF
C4687 a_43262_60146# vcm 0.62fF
C4688 VDD a_48282_10496# 0.52fF
C4689 pmat.row_n[10] pmat.row_n[6] 5.34fF
C4690 a_1781_9308# a_26479_32117# 1.55fF
C4691 VDD a_20438_35431# 2.77fF
C4692 pmat.col_n[13] pmat.col[13] 0.75fF
C4693 VDD a_41703_29423# 0.31fF
C4694 a_18546_7482# a_22086_7890# 0.35fF
C4695 VDD a_7935_20719# 0.47fF
C4696 a_19584_52423# a_12263_50959# 0.42fF
C4697 a_5682_56311# a_11202_55687# 0.58fF
C4698 a_36234_10496# a_37238_10496# 0.97fF
C4699 VDD a_17867_34473# 0.62fF
C4700 a_23395_53135# a_26891_28327# 0.52fF
C4701 _1187_.A2 a_30571_50959# 0.30fF
C4702 VDD a_28202_12504# 0.52fF
C4703 a_49286_16520# vcm 0.65fF
C4704 cgen.dlycontrol4_in[1] a_12237_38772# 0.48fF
C4705 a_47278_56130# a_48282_56130# 0.97fF
C4706 a_41254_13508# ctopn 3.58fF
C4707 _1192_.B1 _1184_.A2 0.48fF
C4708 a_36234_57134# vcm 0.62fF
C4709 a_35230_71190# vcm 0.60fF
C4710 a_39246_18528# ctopn 3.58fF
C4711 VDD a_28281_41245# 1.27fF
C4712 a_22178_58138# vcm 0.62fF
C4713 VDD a_20221_40835# 3.45fF
C4714 VDD a_23663_39913# 0.61fF
C4715 VDD vcm.sky130_fd_sc_hd__buf_4_3.X 0.74fF
C4716 a_1923_69823# a_2407_49289# 0.40fF
C4717 a_50290_15516# ctopn 3.43fF
C4718 VDD a_50290_11500# 0.56fF
C4719 VDD a_1591_50095# 0.43fF
C4720 nmat.rowoff_n[8] nmat.rowoff_n[5] 0.77fF
C4721 VDD m3_51196_11362# 0.34fF
C4722 a_29206_22544# a_30210_22544# 0.97fF
C4723 VDD a_3325_43023# 0.66fF
C4724 VDD a_2847_16127# 0.70fF
C4725 VDD m2_17932_24282# 1.23fF
C4726 ANTENNA__1190__A1.DIODE a_43776_30287# 1.40fF
C4727 ANTENNA__1190__B1.DIODE a_35244_32411# 0.58fF
C4728 a_18546_69224# a_50198_69182# 0.35fF
C4729 VDD a_1823_77821# 0.56fF
C4730 a_11051_8903# a_9583_10121# 0.68fF
C4731 pmat.sample_n pmat.rowoff_n[8] 1.11fF
C4732 VDD pmat.col_n[27] 5.49fF
C4733 a_10814_29111# comp_latch 1.35fF
C4734 ANTENNA__1197__B.DIODE a_21279_48999# 1.11fF
C4735 a_2149_45717# a_2263_43719# 1.37fF
C4736 VDD a_10239_14183# 17.04fF
C4737 a_18546_23546# a_19074_23954# 0.35fF
C4738 a_43262_63158# a_44266_63158# 0.97fF
C4739 a_18546_9490# a_24094_9898# 0.35fF
C4740 a_47278_22544# vcm 0.65fF
C4741 pmat.row_n[4] a_18162_60186# 25.57fF
C4742 a_45270_68178# ctopp 3.58fF
C4743 _1187_.A2 a_46947_39215# 0.51fF
C4744 a_23182_59142# vcm 0.62fF
C4745 _1192_.B1 a_9411_2215# 2.74fF
C4746 a_10515_15055# pmat.row_n[3] 0.75fF
C4747 a_20170_13508# vcm 0.65fF
C4748 a_2407_49289# a_3967_56311# 0.50fF
C4749 VDD a_46233_43023# 0.42fF
C4750 a_23933_32143# a_25575_31055# 0.51fF
C4751 pmat.rowoff_n[0] ctopp 0.51fF
C4752 VDD a_27198_56130# 0.55fF
C4753 pmat.row_n[15] pmat.row_n[13] 0.33fF
C4754 a_30999_48071# a_31152_48071# 0.80fF
C4755 VDD a_2021_11043# 5.85fF
C4756 a_1899_35051# pmat.rowon_n[8] 1.78fF
C4757 VDD nmat.col_n[24] 10.45fF
C4758 VDD m2_42028_7214# 0.93fF
C4759 a_1823_76181# a_2791_57703# 0.36fF
C4760 VDD a_9457_51163# 0.47fF
C4761 a_18546_62196# a_41162_62154# 0.35fF
C4762 VDD a_47407_47919# 0.43fF
C4763 a_18546_66212# a_37146_66170# 0.35fF
C4764 a_21174_66170# ctopp 3.58fF
C4765 VDD a_30210_66170# 0.52fF
C4766 ANTENNA__1395__A1.DIODE _1183_.A2 1.10fF
C4767 a_38242_11500# a_39246_11500# 0.97fF
C4768 a_18162_56170# vcm 6.97fF
C4769 VDD a_18769_36965# 1.27fF
C4770 a_27763_27221# nmat.col[9] 0.32fF
C4771 VDD a_1643_71829# 0.36fF
C4772 a_2648_29397# a_8305_20871# 0.36fF
C4773 VDD a_23182_63158# 0.52fF
C4774 a_40250_64162# a_40250_63158# 1.00fF
C4775 a_24407_31375# nmat.col[28] 0.46fF
C4776 a_43262_10496# a_43262_9492# 1.00fF
C4777 a_18546_61192# a_22086_61150# 0.35fF
C4778 a_16311_28327# a_21739_29415# 1.40fF
C4779 nmat.rowon_n[15] vcm 0.54fF
C4780 a_40250_58138# a_40250_57134# 1.00fF
C4781 pmat.rowon_n[8] a_6554_43255# 0.50fF
C4782 VDD a_26239_39095# 0.63fF
C4783 a_1781_9308# a_5179_31591# 0.52fF
C4784 VDD a_11113_39747# 5.09fF
C4785 a_10949_42364# a_10651_42035# 0.92fF
C4786 a_23182_19532# vcm 0.65fF
C4787 a_47278_62154# pmat.col[28] 0.31fF
C4788 a_20170_55126# ctopp 0.57fF
C4789 a_44266_60146# a_44266_59142# 1.00fF
C4790 a_32218_18528# a_32218_17524# 1.00fF
C4791 nmat.sw a_8031_13353# 0.79fF
C4792 VDD a_12079_31061# 0.46fF
C4793 a_13459_28111# nmat.col[15] 2.32fF
C4794 VDD cgen.dlycontrol1_in[0] 7.80fF
C4795 a_6927_30503# a_4075_31591# 2.51fF
C4796 a_22178_10496# vcm 0.65fF
C4797 a_50290_22544# ctopn 3.42fF
C4798 a_12197_43746# cgen.dlycontrol4_in[0] 0.44fF
C4799 a_32218_63158# a_32218_62154# 1.00fF
C4800 a_26194_71190# m2_25964_72014# 1.00fF
C4801 a_48282_67174# a_49286_67174# 0.97fF
C4802 VDD a_4043_22869# 0.42fF
C4803 VDD a_6061_38377# 0.35fF
C4804 nmat.col[2] vcm 5.76fF
C4805 a_21365_27247# nmat.col_n[18] 0.31fF
C4806 a_18546_70228# a_39154_70186# 0.35fF
C4807 pmat.row_n[15] pmat.row_n[11] 0.35fF
C4808 VDD a_28202_67174# 0.52fF
C4809 a_18546_57176# vcm 0.40fF
C4810 VDD a_12197_38306# 2.51fF
C4811 a_45270_66170# a_45270_65166# 1.00fF
C4812 a_38242_22544# a_38242_21540# 1.00fF
C4813 VDD a_12116_39783# 3.37fF
C4814 a_37238_14512# a_38242_14512# 0.97fF
C4815 a_38242_62154# vcm 0.62fF
C4816 a_36234_64162# a_37238_64162# 0.97fF
C4817 a_18546_17522# a_34134_17930# 0.35fF
C4818 a_4719_30287# cgen.dlycontrol1_in[0] 0.93fF
C4819 a_42258_68178# a_43262_68178# 0.97fF
C4820 a_5651_66975# a_11797_60431# 0.76fF
C4821 a_18546_57176# a_30118_57134# 0.35fF
C4822 a_31214_13508# a_31214_12504# 1.00fF
C4823 a_10471_12791# a_10443_12879# 0.34fF
C4824 a_20170_22544# a_21174_22544# 0.97fF
C4825 a_12116_39783# a_14773_39394# 1.81fF
C4826 nmat.rowon_n[9] vcm 0.56fF
C4827 a_18546_15514# a_34134_15922# 0.35fF
C4828 nmat.rowon_n[7] cgen.dlycontrol4_in[2] 0.33fF
C4829 a_5784_52423# cgen.enable_dlycontrol_in 0.74fF
C4830 cgen.dlycontrol2_in[2] a_12585_39355# 4.14fF
C4831 nmat.rowon_n[14] a_2199_13887# 1.61fF
C4832 a_11041_36596# a_11113_36483# 0.73fF
C4833 VDD a_40951_31599# 1.13fF
C4834 a_37238_70186# vcm 0.62fF
C4835 a_37820_30485# a_44774_48695# 0.80fF
C4836 a_24186_11500# vcm 0.65fF
C4837 ANTENNA__1395__A2.DIODE a_37820_30485# 1.36fF
C4838 _1179_.X _1519_.A 3.31fF
C4839 a_10515_15055# a_10839_11989# 0.42fF
C4840 VDD a_2847_18303# 0.65fF
C4841 a_1586_18231# a_2564_21959# 1.36fF
C4842 m2_47048_24282# m3_47180_24414# 2.79fF
C4843 a_25695_28111# a_42791_32375# 0.67fF
C4844 VDD ctopn 93.62fF
C4845 a_35186_47375# a_36539_47113# 0.46fF
C4846 ANTENNA__1190__A1.DIODE nmat.col_n[18] 5.26fF
C4847 a_26194_19532# ctopn 3.58fF
C4848 pmat.col_n[19] pmat.col[20] 6.04fF
C4849 VDD a_26194_21540# 0.52fF
C4850 nmat.sw a_1858_25615# 1.76fF
C4851 pmat.rowon_n[3] a_1957_43567# 0.66fF
C4852 a_18546_59184# a_50198_59142# 0.35fF
C4853 a_38242_65166# a_38242_64162# 1.00fF
C4854 a_25190_10496# ctopn 3.58fF
C4855 a_46274_57134# ctopp 3.57fF
C4856 a_18546_68220# a_21082_68178# 0.35fF
C4857 VDD a_10147_29415# 8.73fF
C4858 a_45270_71190# ctopp 3.40fF
C4859 a_32218_58138# ctopp 3.58fF
C4860 a_28202_68178# vcm 0.62fF
C4861 VDD a_1644_70197# 0.32fF
C4862 a_11067_30287# a_13643_29415# 0.30fF
C4863 a_5784_52423# a_5211_57172# 0.64fF
C4864 VDD a_41254_58138# 0.52fF
C4865 a_47278_23548# a_48282_23548# 0.97fF
C4866 a_12069_38517# a_15921_38550# 0.42fF
C4867 a_20170_62154# a_21174_62154# 0.97fF
C4868 a_27198_16520# a_27198_15516# 1.00fF
C4869 a_45270_71190# m2_45040_72014# 1.00fF
C4870 VDD a_33905_48463# 0.38fF
C4871 a_18546_66212# a_18162_66210# 2.62fF
C4872 a_49286_9492# a_50290_9492# 0.97fF
C4873 _1224_.X ANTENNA__1187__B1.DIODE 2.86fF
C4874 a_18546_60188# a_26102_60146# 0.35fF
C4875 _1154_.X a_15667_27239# 1.37fF
C4876 VDD a_3727_66113# 0.47fF
C4877 VDD a_26957_37691# 1.31fF
C4878 nmat.col[24] nmat.col[18] 3.19fF
C4879 a_44444_32233# a_45908_33749# 0.37fF
C4880 m2_39016_7214# m3_39148_7346# 2.79fF
C4881 a_26891_28327# a_30663_50087# 0.67fF
C4882 a_28915_50959# a_25879_31591# 0.75fF
C4883 a_15101_29423# a_22459_28879# 0.75fF
C4884 a_23821_35279# a_22537_36911# 1.59fF
C4885 a_1781_9308# a_2683_22089# 0.40fF
C4886 nmat.rowoff_n[2] ctopn 0.60fF
C4887 a_33222_23548# vcm 0.65fF
C4888 nmat.col[23] nmat.col_n[23] 0.73fF
C4889 nmat.col_n[26] nmat.col[25] 0.30fF
C4890 a_24186_69182# ctopp 3.58fF
C4891 a_19166_19532# a_20170_19532# 0.97fF
C4892 m2_17932_55950# m2_17932_54946# 0.99fF
C4893 a_35230_9492# vcm 0.65fF
C4894 VDD a_33222_69182# 0.52fF
C4895 a_16083_50069# a_11067_30287# 1.07fF
C4896 a_11067_30287# nmat.en_bit_n[0] 0.98fF
C4897 pmat.row_n[15] a_2659_35015# 0.74fF
C4898 a_11389_40443# a_11041_40948# 4.69fF
C4899 VDD a_27411_46805# 0.60fF
C4900 a_39246_65166# a_40250_65166# 0.97fF
C4901 a_33222_59142# ctopp 3.58fF
C4902 a_27198_11500# ctopn 3.58fF
C4903 VDD a_42258_59142# 0.52fF
C4904 a_46274_21540# a_47278_21540# 0.97fF
C4905 VDD a_21621_35515# 1.42fF
C4906 VDD a_7663_71317# 0.49fF
C4907 VDD vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top 114.92fF
C4908 ANTENNA__1196__A2.DIODE _1183_.A2 0.48fF
C4909 a_18546_16518# a_38150_16926# 0.35fF
C4910 nmat.rowon_n[14] config_1_in[0] 0.33fF
C4911 a_6283_31591# a_2411_33749# 1.40fF
C4912 a_47278_71190# a_47278_70186# 1.00fF
C4913 a_12309_38659# a_14600_37607# 1.93fF
C4914 VDD pmat.row_n[10] 16.25fF
C4915 pmat.col_n[29] vcm 2.80fF
C4916 a_31214_13508# vcm 0.65fF
C4917 VDD a_19689_42405# 1.17fF
C4918 a_24407_31375# a_38905_28853# 0.45fF
C4919 m2_47048_7214# m2_48052_7214# 0.96fF
C4920 a_29206_18528# vcm 0.65fF
C4921 a_10767_39087# a_13909_39605# 1.28fF
C4922 a_11113_40835# a_20221_40835# 1.86fF
C4923 VDD a_1761_4399# 0.69fF
C4924 nmat.col[7] nmat.rowon_n[1] 0.46fF
C4925 a_3663_9269# a_5558_9527# 0.50fF
C4926 pmat.rowoff_n[8] a_22499_49783# 0.42fF
C4927 pmat.rowon_n[14] ctopp 1.57fF
C4928 a_26583_34343# cgen.dlycontrol1_in[3] 0.83fF
C4929 a_1674_68047# a_6795_76989# 0.49fF
C4930 VDD a_8111_11209# 0.53fF
C4931 a_45270_13508# a_46274_13508# 0.97fF
C4932 VDD m3_39148_72146# 0.41fF
C4933 a_40250_15516# vcm 0.65fF
C4934 VDD a_25190_17524# 0.52fF
C4935 a_24833_40719# cgen.dlycontrol2_in[4] 2.20fF
C4936 a_6787_47607# pmat.row_n[15] 0.42fF
C4937 ANTENNA__1395__A1.DIODE ANTENNA__1395__A2.DIODE 0.35fF
C4938 _1183_.A2 a_41926_46983# 1.10fF
C4939 a_49286_63158# pmat.col[30] 0.31fF
C4940 a_11041_38772# a_16381_35286# 0.82fF
C4941 m2_30984_72014# m3_31116_72146# 2.79fF
C4942 a_30571_50959# a_13275_48783# 0.88fF
C4943 a_43262_18528# a_44266_18528# 0.97fF
C4944 VDD a_4707_32156# 1.72fF
C4945 _0467_ nmat.col[3] 0.41fF
C4946 VDD a_26194_8488# 0.55fF
C4947 a_18546_21538# a_29114_21946# 0.35fF
C4948 a_19166_70186# vcm 0.61fF
C4949 a_30210_62154# a_30210_61150# 1.00fF
C4950 a_36234_23548# ctopn 3.44fF
C4951 a_2263_43719# a_6467_29415# 1.08fF
C4952 VDD a_42258_19532# 0.52fF
C4953 a_38242_9492# ctopn 3.57fF
C4954 _1194_.A2 _1187_.A2 3.97fF
C4955 a_11091_26311# nmat.col[1] 0.41fF
C4956 VDD pmat.rowon_n[12] 3.84fF
C4957 a_4979_38127# a_5935_46983# 0.40fF
C4958 inp_analog _1179_.X 0.66fF
C4959 a_36234_60146# vcm 0.62fF
C4960 VDD a_41254_10496# 0.52fF
C4961 VDD a_17154_43671# 1.29fF
C4962 VDD a_51202_16926# 0.31fF
C4963 a_7693_22365# comp_latch 1.28fF
C4964 ANTENNA__1187__B1.DIODE comp_latch 0.45fF
C4965 a_30210_15516# a_30210_14512# 1.00fF
C4966 m2_51064_16250# m3_51196_16382# 2.76fF
C4967 VDD a_5462_62215# 3.80fF
C4968 a_18546_7482# a_18162_7484# 2.62fF
C4969 VDD a_10498_19631# 0.74fF
C4970 a_41254_63158# pmat.col[22] 0.31fF
C4971 a_18546_58180# a_48190_58138# 0.35fF
C4972 a_32218_69182# a_32218_68178# 1.00fF
C4973 VDD a_15101_29423# 2.27fF
C4974 a_18546_10494# a_48190_10902# 0.35fF
C4975 a_40250_21540# a_40250_20536# 1.00fF
C4976 a_18546_20534# a_20078_20942# 0.35fF
C4977 pmat.rowon_n[6] pmat.rowoff_n[6] 20.90fF
C4978 VDD a_21174_12504# 0.52fF
C4979 a_48282_62154# ctopp 3.58fF
C4980 a_42258_16520# vcm 0.65fF
C4981 nmat.col[20] ctopn 1.97fF
C4982 VDD a_21279_48999# 7.70fF
C4983 a_34226_13508# ctopn 3.58fF
C4984 a_16981_37462# a_21219_36885# 0.49fF
C4985 a_29206_57134# vcm 0.62fF
C4986 a_41227_29423# inn_analog 0.99fF
C4987 VDD a_39981_37462# 1.25fF
C4988 a_28202_71190# vcm 0.60fF
C4989 pmat.row_n[0] nmat.col[13] 0.31fF
C4990 a_32218_18528# ctopn 3.58fF
C4991 pmat.row_n[6] ctopp 1.65fF
C4992 a_13091_28327# a_10883_3303# 0.82fF
C4993 a_18243_28327# a_25695_28111# 3.52fF
C4994 nmat.col[21] nmat.col[19] 12.15fF
C4995 a_47278_70186# ctopp 3.57fF
C4996 nmat.rowoff_n[3] vcm 0.30fF
C4997 a_43262_15516# ctopn 3.58fF
C4998 VDD a_43262_11500# 0.52fF
C4999 m3_50192_55078# ctopp 0.37fF
C5000 ANTENNA__1395__A1.DIODE ANTENNA__1196__A2.DIODE 0.58fF
C5001 a_14641_57167# pmat.rowon_n[6] 0.38fF
C5002 VDD a_4257_34319# 1.75fF
C5003 a_19166_14512# vcm 0.65fF
C5004 a_18546_64204# vcm 0.40fF
C5005 m2_17932_11230# m2_17932_10226# 0.99fF
C5006 pmat.rowon_n[3] nmat.rowon_n[1] 0.91fF
C5007 VDD a_14839_54599# 0.37fF
C5008 pmat.row_n[7] a_10515_15055# 0.90fF
C5009 a_18546_69224# a_43170_69182# 0.35fF
C5010 VDD a_41427_31599# 0.44fF
C5011 a_5363_70543# a_11435_58791# 0.90fF
C5012 a_34226_11500# a_34226_10496# 1.00fF
C5013 nmat.col_n[13] a_9441_20189# 0.56fF
C5014 a_3866_57399# a_6175_60039# 0.44fF
C5015 a_11067_27239# _1194_.B1 0.90fF
C5016 VDD a_19166_18528# 0.56fF
C5017 m2_18936_54946# vcm 0.41fF
C5018 a_6559_33767# a_6007_33767# 1.05fF
C5019 a_40250_22544# vcm 0.65fF
C5020 a_11067_16359# a_10515_13967# 9.51fF
C5021 a_39246_61150# a_40250_61150# 0.97fF
C5022 a_38242_68178# ctopp 3.58fF
C5023 pmat.rowoff_n[7] a_1739_47893# 0.56fF
C5024 a_29937_31055# a_40837_46261# 1.02fF
C5025 VDD a_47278_68178# 0.52fF
C5026 a_24186_12504# a_24186_11500# 1.00fF
C5027 a_20170_22544# a_20170_21540# 1.00fF
C5028 a_7717_14735# a_4339_27804# 0.92fF
C5029 nmat.rowoff_n[6] a_6830_22895# 1.47fF
C5030 VDD a_25997_42902# 1.03fF
C5031 m2_51064_13238# m3_51196_13370# 2.76fF
C5032 a_7717_14735# a_13641_23439# 1.15fF
C5033 a_38905_28853# a_17842_27497# 0.93fF
C5034 VDD a_15299_28879# 0.31fF
C5035 a_18546_64204# a_19074_64162# 0.35fF
C5036 a_1957_43567# a_5363_33551# 0.48fF
C5037 a_11057_35836# a_6007_33767# 2.30fF
C5038 VDD a_20170_56130# 0.54fF
C5039 a_33222_20536# a_34226_20536# 0.97fF
C5040 a_18546_20534# a_49194_20942# 0.35fF
C5041 a_45270_16520# ctopn 3.58fF
C5042 a_8443_20719# a_9441_20189# 1.81fF
C5043 VDD m2_27972_7214# 1.06fF
C5044 a_2263_43719# a_18869_46831# 0.35fF
C5045 VDD a_5715_16911# 0.35fF
C5046 ANTENNA__1184__B1.DIODE a_9963_28111# 0.32fF
C5047 VDD a_1591_74031# 0.92fF
C5048 a_3571_13627# a_2199_13887# 0.33fF
C5049 a_18546_62196# a_34134_62154# 0.35fF
C5050 a_18546_66212# a_30118_66170# 0.35fF
C5051 a_46274_67174# a_46274_66170# 1.00fF
C5052 a_32218_9492# a_32218_8488# 1.00fF
C5053 VDD a_23182_66170# 0.52fF
C5054 VDD a_2847_8511# 0.44fF
C5055 a_32405_32463# a_18241_31698# 0.32fF
C5056 a_24591_28327# a_28915_50959# 2.18fF
C5057 a_14600_37607# cgen.dlycontrol1_in[4] 2.67fF
C5058 a_46274_56130# m2_46044_54946# 0.99fF
C5059 a_45270_17524# a_46274_17524# 0.97fF
C5060 m2_51064_60970# vcm 0.51fF
C5061 a_20170_9492# ctopn 3.56fF
C5062 a_1957_43567# a_11202_55687# 0.34fF
C5063 a_43262_57134# a_44266_57134# 0.97fF
C5064 a_48282_20536# a_48282_19532# 1.00fF
C5065 a_42258_71190# a_43262_71190# 0.97fF
C5066 a_22178_62154# pmat.col[3] 0.31fF
C5067 a_29206_58138# a_30210_58138# 0.97fF
C5068 VDD a_20995_44265# 0.64fF
C5069 a_48282_14512# vcm 0.65fF
C5070 a_11435_58791# a_3688_17179# 0.95fF
C5071 a_47278_64162# vcm 0.62fF
C5072 pmat.col_n[11] m2_29980_54946# 0.37fF
C5073 a_26479_32117# a_31263_32117# 0.43fF
C5074 a_46274_8488# a_47278_8488# 0.97fF
C5075 VDD vcm.sky130_fd_sc_hd__buf_4_2.X 0.72fF
C5076 a_13459_28111# a_38793_49007# 0.40fF
C5077 VDD a_13985_34789# 1.35fF
C5078 ANTENNA__1395__A2.DIODE ANTENNA__1196__A2.DIODE 19.84fF
C5079 ANTENNA__1184__B1.DIODE ANTENNA__1195__A1.DIODE 1.57fF
C5080 a_24867_53135# a_16311_28327# 1.26fF
C5081 a_24591_28327# ANTENNA__1395__B1.DIODE 0.91fF
C5082 VDD a_18546_71232# 32.69fF
C5083 VDD a_50290_13508# 0.54fF
C5084 a_14641_57167# a_11067_64015# 0.64fF
C5085 a_18546_58180# a_18162_58178# 2.62fF
C5086 a_12461_29673# a_17702_29967# 0.83fF
C5087 a_43262_22544# ctopn 3.57fF
C5088 VDD a_48282_18528# 0.52fF
C5089 pmat.col[18] vcm 5.88fF
C5090 a_29206_61150# a_29206_60146# 1.00fF
C5091 a_37238_19532# a_37238_18528# 1.00fF
C5092 a_18546_70228# a_32126_70186# 0.35fF
C5093 VDD a_21174_67174# 0.52fF
C5094 nmat.col_n[21] nmat.col_n[31] 1.12fF
C5095 pmat.rowon_n[8] a_10515_61839# 1.35fF
C5096 a_15667_27239# nmat.col_n[0] 0.49fF
C5097 ANTENNA__1197__A.DIODE pmat.col[17] 0.68fF
C5098 a_18546_14510# a_50198_14918# 0.35fF
C5099 a_31214_62154# vcm 0.62fF
C5100 m2_51064_10226# m3_51196_10358# 2.76fF
C5101 a_18546_64204# a_48190_64162# 0.35fF
C5102 a_18546_17522# a_27106_17930# 0.35fF
C5103 nmat.rowon_n[1] nmat.rowoff_n[5] 0.72fF
C5104 VDD a_82736_4943# 0.64fF
C5105 a_18546_57176# a_23090_57134# 0.35fF
C5106 a_30210_59142# a_30210_58138# 1.00fF
C5107 VDD a_2124_52931# 0.64fF
C5108 a_35230_8488# m2_35000_7214# 1.00fF
C5109 a_18546_72236# a_40158_72194# 0.35fF
C5110 ANTENNA__1395__A2.DIODE a_11337_25071# 0.55fF
C5111 a_22178_15516# a_23182_15516# 0.97fF
C5112 a_18546_15514# a_27106_15922# 0.35fF
C5113 a_50290_65166# vcm 0.62fF
C5114 _1179_.X a_28915_50959# 1.69fF
C5115 VDD a_22567_47381# 0.51fF
C5116 a_2149_45717# a_2215_47375# 0.58fF
C5117 a_46274_60146# ctopp 3.58fF
C5118 a_21174_69182# a_22178_69182# 0.97fF
C5119 a_30210_70186# vcm 0.62fF
C5120 VDD a_26102_72194# 0.32fF
C5121 a_10883_3303# a_11927_27399# 1.35fF
C5122 a_4703_24527# a_3305_15823# 1.10fF
C5123 a_1591_23445# a_1757_23445# 0.57fF
C5124 a_13357_37429# ndecision_finish 0.82fF
C5125 VDD a_1895_18170# 0.51fF
C5126 a_35230_17524# a_35230_16520# 1.00fF
C5127 nmat.col[30] ANTENNA__1190__A2.DIODE 11.44fF
C5128 nmat.col_n[31] inn_analog 0.34fF
C5129 pmat.rowon_n[0] pmat.row_n[0] 20.83fF
C5130 VDD a_13683_24847# 0.34fF
C5131 a_10055_31591# a_6467_29415# 1.25fF
C5132 a_41254_12504# a_42258_12504# 0.97fF
C5133 a_11948_49783# a_1781_9308# 0.79fF
C5134 a_30571_50959# a_25695_28111# 0.97fF
C5135 a_14839_54599# pmat.rowoff_n[1] 0.40fF
C5136 _1196_.B1 vcm 0.44fF
C5137 a_1781_9308# a_2046_30184# 0.34fF
C5138 a_2124_31867# a_2422_29575# 0.47fF
C5139 _1179_.X ANTENNA__1395__B1.DIODE 3.37fF
C5140 a_30210_59142# a_31214_59142# 0.97fF
C5141 a_9963_13967# a_12447_16143# 2.54fF
C5142 pmat.rowon_n[3] pmat.row_n[2] 0.37fF
C5143 a_18546_59184# a_43170_59142# 0.35fF
C5144 pmat.rowoff_n[4] a_13091_7655# 2.09fF
C5145 a_39246_57134# ctopp 3.57fF
C5146 a_4991_69831# a_5363_33551# 0.76fF
C5147 a_38242_71190# ctopp 3.40fF
C5148 VDD a_48282_57134# 0.52fF
C5149 a_35244_32411# clk_ena 0.48fF
C5150 a_25190_58138# ctopp 3.58fF
C5151 a_21174_68178# vcm 0.62fF
C5152 VDD a_47278_71190# 0.55fF
C5153 VDD a_34226_58138# 0.52fF
C5154 m2_18936_23278# ctopn 0.36fF
C5155 a_10055_31591# a_13091_52047# 0.97fF
C5156 a_10781_42869# a_11021_43011# 1.54fF
C5157 VDD a_29076_48695# 1.96fF
C5158 _1196_.B1 _1194_.B1 0.55fF
C5159 VDD pmat.rowon_n[4] 3.65fF
C5160 a_21739_29415# a_24407_31375# 2.90fF
C5161 VDD a_14719_37737# 0.61fF
C5162 nmat.col_n[12] nmat.col[12] 0.74fF
C5163 a_1586_50247# a_6082_46831# 0.38fF
C5164 _1184_.A2 a_10883_3303# 2.04fF
C5165 a_16311_28327# a_38851_28327# 0.31fF
C5166 a_18546_24550# a_48190_24958# 0.35fF
C5167 a_8583_29199# a_10147_29415# 0.36fF
C5168 nmat.col_n[31] nmat.col[26] 2.04fF
C5169 VDD a_26773_40955# 1.36fF
C5170 VDD a_35108_39655# 1.32fF
C5171 a_26194_68178# a_26194_67174# 1.00fF
C5172 a_26194_23548# vcm 0.65fF
C5173 a_10515_13967# a_11067_49871# 0.47fF
C5174 ANTENNA__1395__A1.DIODE nmat.col_n[17] 0.31fF
C5175 a_28202_9492# vcm 0.65fF
C5176 VDD a_26194_69182# 0.52fF
C5177 a_50290_61150# vcm 0.62fF
C5178 VDD a_11803_49551# 0.40fF
C5179 ANTENNA__1395__B1.DIODE a_14917_23983# 0.72fF
C5180 a_45270_23548# m2_45040_24282# 0.99fF
C5181 ANTENNA__1190__A1.DIODE a_15667_27239# 0.47fF
C5182 a_23395_53135# pmat.col[24] 0.47fF
C5183 a_18546_22542# a_45178_22950# 0.35fF
C5184 VDD config_1_in[4] 0.83fF
C5185 VDD a_15107_44535# 0.60fF
C5186 a_6664_26159# a_9303_22351# 0.34fF
C5187 VDD m2_25964_24282# 0.62fF
C5188 a_44266_20536# vcm 0.65fF
C5189 a_26194_59142# ctopp 3.58fF
C5190 VDD nmat.col[14] 4.44fF
C5191 VDD a_18199_52789# 0.35fF
C5192 VDD a_35230_59142# 0.52fF
C5193 VDD pmat.col_n[30] 5.06fF
C5194 cgen.dlycontrol4_in[3] a_12197_43746# 0.67fF
C5195 a_24186_16520# a_25190_16520# 0.97fF
C5196 a_18546_16518# a_31122_16926# 0.35fF
C5197 a_14287_69455# pmat.row_n[1] 0.54fF
C5198 _1192_.A2 a_27763_27221# 0.34fF
C5199 a_4339_27804# a_9339_28335# 0.34fF
C5200 VDD a_3891_61519# 0.59fF
C5201 a_41731_49525# a_45019_38645# 0.37fF
C5202 a_5403_67655# a_4583_68021# 0.31fF
C5203 a_24186_13508# vcm 0.65fF
C5204 a_27198_62154# pmat.col[8] 0.31fF
C5205 pmat.rowon_n[11] nmat.rowon_n[4] 21.19fF
C5206 m2_40020_7214# m2_41024_7214# 0.96fF
C5207 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot clk_ena 0.32fF
C5208 a_7521_47081# a_6559_33767# 0.64fF
C5209 a_22178_18528# vcm 0.65fF
C5210 a_10883_3303# a_9411_2215# 0.56fF
C5211 _1192_.B1 a_25879_31591# 0.71fF
C5212 ANTENNA__1395__A2.DIODE a_12053_27497# 0.51fF
C5213 a_2407_49289# a_5595_65301# 0.31fF
C5214 VDD a_7779_22583# 3.67fF
C5215 a_33222_15516# vcm 0.65fF
C5216 a_17154_43671# a_12658_42895# 0.31fF
C5217 nmat.rowon_n[7] a_18162_16520# 1.33fF
C5218 a_33222_70186# a_33222_69182# 1.00fF
C5219 VDD a_18162_8488# 2.79fF
C5220 ANTENNA__1190__B1.DIODE _1183_.A2 2.83fF
C5221 VDD ctopp 93.81fF
C5222 a_18546_21538# a_22086_21946# 0.35fF
C5223 a_2835_13077# clk_dig 0.37fF
C5224 a_15753_28879# a_14691_29575# 0.61fF
C5225 a_22178_14512# a_22178_13508# 1.00fF
C5226 cgen.dlycontrol4_in[2] a_2683_22089# 1.32fF
C5227 pmat.en_bit_n[2] a_23021_29199# 0.52fF
C5228 a_29206_23548# ctopn 3.40fF
C5229 VDD a_35230_19532# 0.52fF
C5230 a_31214_9492# ctopn 3.57fF
C5231 _1154_.X _1196_.B1 0.93fF
C5232 VDD m2_45040_72014# 0.98fF
C5233 a_26194_57134# a_26194_56130# 1.00fF
C5234 a_30210_19532# a_31214_19532# 0.97fF
C5235 VDD a_4985_51433# 3.91fF
C5236 a_29206_60146# vcm 0.62fF
C5237 nmat.col_n[28] nmat.col[19] 1.14fF
C5238 VDD a_34226_10496# 0.52fF
C5239 a_1586_63927# a_8031_64789# 0.80fF
C5240 VDD a_39469_39141# 1.42fF
C5241 comp.adc_comp_circuit_0.adc_comp_buffer_0.in a_54136_39932# 0.53fF
C5242 a_47278_20536# ctopn 3.58fF
C5243 VDD a_11261_43421# 1.16fF
C5244 ANTENNA__1187__B1.DIODE ANTENNA__1183__B1.DIODE 2.40fF
C5245 a_18546_63200# vcm 0.40fF
C5246 a_18546_58180# a_41162_58138# 0.35fF
C5247 VDD a_13479_26935# 1.97fF
C5248 VDD a_1761_6031# 0.64fF
C5249 ANTENNA__1187__B1.DIODE nmat.col[25] 0.59fF
C5250 a_13459_28111# a_38695_48634# 0.38fF
C5251 a_18546_10494# a_41162_10902# 0.35fF
C5252 a_29206_10496# a_30210_10496# 0.97fF
C5253 a_7521_47081# a_8385_51727# 0.52fF
C5254 a_30111_47911# a_33423_47695# 1.50fF
C5255 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top 0.43fF
C5256 a_41254_62154# ctopp 3.58fF
C5257 a_18546_13506# a_18162_13508# 2.61fF
C5258 VDD a_50290_62154# 0.54fF
C5259 a_35230_16520# vcm 0.65fF
C5260 VDD a_47591_49007# 0.45fF
C5261 nmat.rowon_n[14] cgen.dlycontrol4_in[0] 0.53fF
C5262 a_40250_56130# a_41254_56130# 0.97fF
C5263 a_4985_51433# a_4719_30287# 0.66fF
C5264 a_11435_58791# a_9963_13967# 0.98fF
C5265 a_27198_13508# ctopn 3.58fF
C5266 pmat.row_n[14] pmat.row_n[12] 14.77fF
C5267 VDD vcm.sky130_fd_sc_hd__buf_4_1.X 1.01fF
C5268 a_22178_57134# vcm 0.62fF
C5269 VDD a_23329_37462# 1.15fF
C5270 a_21174_71190# vcm 0.60fF
C5271 a_25190_18528# ctopn 3.58fF
C5272 VDD a_32035_42089# 0.65fF
C5273 nmat.col_n[31] clk_ena 0.43fF
C5274 a_2419_53351# pmat.rowoff_n[7] 0.81fF
C5275 m2_17932_63982# vcm 0.44fF
C5276 nmat.col_n[2] ctopn 2.02fF
C5277 a_40250_70186# ctopp 3.57fF
C5278 VDD a_1586_50247# 12.07fF
C5279 VDD a_49286_70186# 0.52fF
C5280 a_36234_15516# ctopn 3.58fF
C5281 a_37820_30485# a_7109_29423# 0.48fF
C5282 a_30111_47911# a_36324_46983# 0.30fF
C5283 a_8583_47381# a_8749_47381# 0.46fF
C5284 pmat.col_n[2] pmat.col[3] 6.03fF
C5285 VDD a_36234_11500# 0.52fF
C5286 a_7067_53511# a_7163_53333# 0.37fF
C5287 a_11067_27239# a_40837_46261# 0.62fF
C5288 a_6787_47607# a_5363_33551# 0.63fF
C5289 a_22178_22544# a_23182_22544# 0.97fF
C5290 a_19166_12504# m2_17932_12234# 0.96fF
C5291 a_12237_38772# a_12116_40871# 0.44fF
C5292 VDD a_5351_19913# 9.90fF
C5293 a_45270_62154# a_46274_62154# 0.97fF
C5294 VDD m2_21948_54946# 0.62fF
C5295 VDD a_35186_47375# 3.90fF
C5296 a_43262_66170# a_44266_66170# 0.97fF
C5297 VDD a_10239_77295# 0.88fF
C5298 a_18546_69224# a_36142_69182# 0.35fF
C5299 VDD a_3746_58487# 9.16fF
C5300 a_10873_36341# a_15049_36374# 0.77fF
C5301 a_40837_46261# a_35312_31599# 0.72fF
C5302 VDD a_4307_35639# 0.59fF
C5303 a_10883_3303# nmat.col[13] 0.45fF
C5304 a_20170_55126# pmat.col[1] 0.41fF
C5305 a_11113_38659# a_10927_37981# 1.06fF
C5306 ANTENNA__1197__A.DIODE _1192_.A2 1.53fF
C5307 VDD a_7809_17705# 0.52fF
C5308 a_36234_63158# a_37238_63158# 0.97fF
C5309 m2_17932_23278# m3_18064_23410# 2.76fF
C5310 nmat.rowon_n[12] a_10593_15823# 0.59fF
C5311 a_33222_22544# vcm 0.65fF
C5312 a_31214_68178# ctopp 3.58fF
C5313 VDD a_40250_68178# 0.52fF
C5314 pmat.col[20] m2_39016_54946# 0.39fF
C5315 a_18243_28327# comp_latch 0.41fF
C5316 pmat.en_bit_n[2] nmat.col_n[13] 0.37fF
C5317 a_4128_64391# a_4707_32156# 0.75fF
C5318 a_47278_63158# vcm 0.62fF
C5319 a_24591_28327# nmat.col[18] 0.30fF
C5320 a_24861_29673# a_20616_27791# 0.89fF
C5321 VDD a_2743_28853# 0.48fF
C5322 ANTENNA__1395__A1.DIODE ANTENNA__1190__B1.DIODE 3.12fF
C5323 a_3746_58487# a_4719_30287# 0.89fF
C5324 nmat.col[10] a_7026_24527# 1.22fF
C5325 a_13091_7655# clk_dig 0.67fF
C5326 a_18546_20534# a_42166_20942# 0.35fF
C5327 ANTENNA__1184__B1.DIODE nmat.col_n[28] 5.69fF
C5328 a_38242_16520# ctopn 3.58fF
C5329 VDD a_1674_57711# 10.46fF
C5330 a_13275_48783# a_32687_46607# 0.70fF
C5331 pmat.rowoff_n[15] pmat.row_n[15] 20.67fF
C5332 nmat.col_n[15] a_34226_24552# 0.31fF
C5333 ANTENNA__1395__A2.DIODE a_2007_25597# 1.16fF
C5334 a_18546_62196# a_27106_62154# 0.35fF
C5335 a_18546_66212# a_23090_66170# 0.35fF
C5336 VDD a_45270_23548# 0.55fF
C5337 a_5462_62215# a_4128_64391# 1.17fF
C5338 a_44266_70186# a_45270_70186# 0.97fF
C5339 VDD a_47278_9492# 0.52fF
C5340 a_13357_37429# cgen.dlycontrol1_in[4] 0.49fF
C5341 a_18546_11498# a_45178_11906# 0.35fF
C5342 a_31214_11500# a_32218_11500# 0.97fF
C5343 VDD a_39045_37692# 1.44fF
C5344 pmat.row_n[5] pmat.row_n[4] 0.37fF
C5345 a_7415_29397# a_4339_27804# 0.87fF
C5346 m2_44036_7214# m3_44168_7346# 2.79fF
C5347 a_13641_23439# a_7415_29397# 1.04fF
C5348 a_9307_31068# a_19439_30511# 0.44fF
C5349 nmat.rowon_n[5] ANTENNA__1183__B1.DIODE 0.43fF
C5350 VDD a_14011_19087# 0.43fF
C5351 a_2879_57487# a_3751_64757# 0.39fF
C5352 a_33222_64162# a_33222_63158# 1.00fF
C5353 nmat.col[25] m2_44036_24282# 0.39fF
C5354 m2_21948_54946# m3_22080_55078# 2.79fF
C5355 a_36234_10496# a_36234_9492# 1.00fF
C5356 a_31675_47695# nmat.col[29] 0.54fF
C5357 a_33222_58138# a_33222_57134# 1.00fF
C5358 ANTENNA__1395__A2.DIODE a_19405_28853# 0.85fF
C5359 VDD a_37731_44527# 0.39fF
C5360 a_41254_14512# vcm 0.65fF
C5361 a_40250_64162# vcm 0.62fF
C5362 pmat.col_n[7] m2_25964_54946# 0.38fF
C5363 VDD m2_49056_24282# 0.64fF
C5364 a_37238_60146# a_37238_59142# 1.00fF
C5365 pmat.rowoff_n[1] ctopp 0.60fF
C5366 a_25190_18528# a_25190_17524# 1.00fF
C5367 VDD a_18546_55168# 36.81fF
C5368 a_20170_10496# a_21174_10496# 0.97fF
C5369 a_26891_28327# a_7717_14735# 0.51fF
C5370 a_6283_31591# a_30111_47911# 0.42fF
C5371 VDD a_43262_13508# 0.52fF
C5372 cgen.dlycontrol3_in[4] a_22085_36374# 0.35fF
C5373 pmat.sw a_36453_29199# 0.74fF
C5374 a_36234_22544# ctopn 3.58fF
C5375 VDD a_41254_18528# 0.52fF
C5376 a_3571_13627# a_9319_15279# 0.42fF
C5377 a_25190_63158# a_25190_62154# 1.00fF
C5378 m2_30984_24282# vcm 0.42fF
C5379 VDD m2_51064_65990# 1.00fF
C5380 VDD a_25743_49783# 0.39fF
C5381 a_41254_67174# a_42258_67174# 0.97fF
C5382 a_2419_53351# a_4421_67477# 0.37fF
C5383 a_18546_70228# a_25098_70186# 0.35fF
C5384 a_7415_29397# a_10223_26703# 0.35fF
C5385 a_38242_66170# a_38242_65166# 1.00fF
C5386 a_31214_22544# a_31214_21540# 1.00fF
C5387 a_2411_33749# a_6099_37039# 0.31fF
C5388 _1194_.B1 a_45019_38645# 0.33fF
C5389 a_24591_28327# _1192_.B1 0.70fF
C5390 ANTENNA__1395__A1.DIODE a_7109_29423# 0.41fF
C5391 a_30210_14512# a_31214_14512# 0.97fF
C5392 a_18546_14510# a_43170_14918# 0.35fF
C5393 a_24186_62154# vcm 0.62fF
C5394 a_29206_64162# a_30210_64162# 0.97fF
C5395 a_18546_64204# a_41162_64162# 0.35fF
C5396 a_35230_68178# a_36234_68178# 0.97fF
C5397 a_1739_47893# cgen.dlycontrol3_in[0] 0.96fF
C5398 pmat.rowoff_n[12] a_11067_16359# 1.16fF
C5399 a_1586_18231# a_5253_18543# 0.49fF
C5400 ANTENNA__1196__A2.DIODE a_2007_25597# 0.71fF
C5401 a_24186_13508# a_24186_12504# 1.00fF
C5402 _1224_.X ANTENNA__1190__A2.DIODE 0.95fF
C5403 a_10873_39605# a_11041_40948# 0.40fF
C5404 a_3339_59879# a_10921_64786# 0.47fF
C5405 a_2648_29397# a_3325_20175# 0.40fF
C5406 a_18546_15514# a_19074_15922# 0.35fF
C5407 a_43262_65166# vcm 0.62fF
C5408 ANTENNA__1190__B1.DIODE ANTENNA__1395__A2.DIODE 20.12fF
C5409 _1187_.A2 ANTENNA__1197__B.DIODE 0.86fF
C5410 ANTENNA__1190__A1.DIODE a_11067_27239# 2.42fF
C5411 VDD a_9839_47679# 0.36fF
C5412 a_50290_21540# vcm 0.65fF
C5413 a_19166_8488# a_20170_8488# 0.97fF
C5414 pmat.row_n[3] a_18162_59182# 25.57fF
C5415 a_39246_60146# ctopp 3.58fF
C5416 m2_36004_72014# m3_36136_72146# 2.79fF
C5417 VDD a_48282_60146# 0.52fF
C5418 pmat.rowon_n[2] pmat.rowoff_n[4] 0.60fF
C5419 a_12237_36596# a_12069_36341# 1.44fF
C5420 a_9279_71829# a_9375_72007# 0.83fF
C5421 a_23182_70186# vcm 0.62fF
C5422 pmat.sw nmat.col_n[31] 1.28fF
C5423 a_22199_30287# a_41731_49525# 0.47fF
C5424 a_44266_14512# ctopn 3.58fF
C5425 a_30663_50087# a_25879_31591# 0.60fF
C5426 VDD cgen.start_conv_in 9.13fF
C5427 VDD pmat.rowon_n[7] 12.80fF
C5428 VDD m2_17932_20266# 1.01fF
C5429 VDD a_17306_28879# 0.80fF
C5430 _1196_.B1 a_40837_46261# 0.69fF
C5431 a_18546_59184# a_36142_59142# 0.35fF
C5432 a_10055_31591# nmat.rowon_n[7] 2.45fF
C5433 a_31214_65166# a_31214_64162# 1.00fF
C5434 a_32218_57134# ctopp 3.57fF
C5435 a_31214_71190# ctopp 3.40fF
C5436 VDD a_41254_57134# 0.52fF
C5437 pmat.rowoff_n[12] vcm 0.84fF
C5438 VDD a_40250_71190# 0.55fF
C5439 a_20170_16520# ctopn 3.57fF
C5440 nmat.sw clk_dig 0.84fF
C5441 VDD a_27198_58138# 0.52fF
C5442 VDD a_2655_72373# 0.41fF
C5443 a_10055_31591# a_14653_53458# 0.40fF
C5444 a_40250_23548# a_41254_23548# 0.97fF
C5445 cgen.dlycontrol4_in[1] a_2021_26677# 2.03fF
C5446 a_11041_38772# a_11225_35836# 3.80fF
C5447 a_42258_9492# a_43262_9492# 0.97fF
C5448 a_49286_12504# a_49286_11500# 1.00fF
C5449 _1192_.B1 a_33423_47695# 1.18fF
C5450 cgen.dlycontrol2_in[3] a_11681_35823# 0.44fF
C5451 a_4351_55527# a_4587_53505# 0.35fF
C5452 VDD a_17113_41317# 1.15fF
C5453 a_29206_56130# m2_28976_54946# 0.99fF
C5454 a_18546_24550# a_41162_24958# 0.35fF
C5455 a_19283_49783# a_28901_48437# 0.55fF
C5456 VDD a_16671_39913# 0.61fF
C5457 a_18162_23548# vcm 6.97fF
C5458 a_21174_9492# vcm 0.65fF
C5459 a_43262_61150# vcm 0.62fF
C5460 a_10515_15055# a_8831_24501# 0.88fF
C5461 ANTENNA__1395__A2.DIODE a_7109_29423# 1.18fF
C5462 ANTENNA__1190__B1.DIODE ANTENNA__1196__A2.DIODE 2.65fF
C5463 a_24867_53135# a_24407_31375# 0.91fF
C5464 ANTENNA__1187__B1.DIODE a_21739_29415# 0.64fF
C5465 a_18546_22542# a_38150_22950# 0.35fF
C5466 a_37820_30485# nmat.col_n[21] 1.01fF
C5467 VDD m2_45040_54946# 0.62fF
C5468 VDD cgen.dlycontrol3_in[1] 7.96fF
C5469 VDD dummypin[5] 0.91fF
C5470 a_37238_20536# vcm 0.65fF
C5471 a_32218_65166# a_33222_65166# 0.97fF
C5472 a_1923_61759# a_1823_66941# 0.56fF
C5473 _1183_.A2 nmat.col_n[21] 8.85fF
C5474 VDD nmat.rowoff_n[1] 3.27fF
C5475 VDD a_28202_59142# 0.52fF
C5476 a_39246_21540# a_40250_21540# 0.97fF
C5477 a_49286_17524# vcm 0.65fF
C5478 cgen.dlycontrol3_in[0] cgen.dlycontrol4_in[0] 0.47fF
C5479 a_18546_16518# a_24094_16926# 0.35fF
C5480 a_9963_13967# a_9528_20407# 0.62fF
C5481 m2_26968_54946# vcm 0.42fF
C5482 a_38851_28327# nmat.col_n[26] 0.41fF
C5483 a_7026_24527# a_12463_22351# 0.31fF
C5484 a_25695_28111# a_42307_31756# 0.33fF
C5485 ANTENNA__1190__A2.DIODE comp_latch 0.32fF
C5486 a_40250_71190# a_40250_70186# 1.00fF
C5487 a_50290_8488# vcm 0.64fF
C5488 ANTENNA__1196__A2.DIODE a_14365_22351# 1.42fF
C5489 a_1586_33927# a_5271_35407# 0.38fF
C5490 VDD a_36345_42567# 1.29fF
C5491 ANTENNA__1197__B.DIODE pmat.col[1] 0.57fF
C5492 pmat.col[29] vcm 5.88fF
C5493 m2_32992_7214# m2_33996_7214# 0.96fF
C5494 a_17139_30503# nmat.col[21] 1.52fF
C5495 ANTENNA__1195__A1.DIODE a_17139_30503# 0.36fF
C5496 a_4075_31591# a_13091_18535# 0.99fF
C5497 a_2659_35015# a_2563_34837# 1.03fF
C5498 a_4075_31591# a_5535_29980# 1.17fF
C5499 VDD a_12067_67279# 0.91fF
C5500 a_11067_30287# a_14379_6567# 2.72fF
C5501 pmat.rowon_n[8] nmat.rowon_n[6] 0.85fF
C5502 a_38242_13508# a_39246_13508# 0.97fF
C5503 a_18546_72236# a_20078_72194# 0.35fF
C5504 VDD nmat.col_n[23] 5.14fF
C5505 a_26194_15516# vcm 0.65fF
C5506 VDD a_11421_17455# 0.37fF
C5507 VDD a_24602_48169# 0.98fF
C5508 a_2163_55233# a_2124_55107# 0.67fF
C5509 cgen.dlycontrol4_in[2] a_1586_18231# 1.09fF
C5510 VDD a_6817_21807# 0.79fF
C5511 a_36234_18528# a_37238_18528# 0.97fF
C5512 a_19166_12504# ctopn 3.43fF
C5513 VDD a_45908_33749# 0.65fF
C5514 VDD a_12257_8527# 0.49fF
C5515 m2_51064_66994# m2_51064_65990# 0.99fF
C5516 a_23182_62154# a_23182_61150# 1.00fF
C5517 cgen.dlycontrol3_in[4] a_12309_38659# 0.44fF
C5518 a_45270_12504# vcm 0.65fF
C5519 a_50290_64162# ctopp 3.43fF
C5520 nmat.col[10] nmat.col_n[10] 0.72fF
C5521 nmat.rowoff_n[13] a_18546_10494# 4.09fF
C5522 nmat.col[15] ctopn 1.99fF
C5523 a_22178_23548# ctopn 3.40fF
C5524 a_25695_28111# a_32687_46607# 0.59fF
C5525 pmat.col[12] vcm 5.88fF
C5526 pmat.sample pmat.row_n[9] 0.44fF
C5527 VDD a_28202_19532# 0.52fF
C5528 a_18546_63200# a_19074_63158# 0.35fF
C5529 a_24186_9492# ctopn 3.57fF
C5530 VDD m2_30984_72014# 1.35fF
C5531 a_12155_27791# a_12175_27221# 0.31fF
C5532 a_5351_19913# a_7840_27247# 1.23fF
C5533 nmat.col[10] clk_ena 0.50fF
C5534 pmat.rowon_n[0] cgen.dlycontrol1_in[3] 1.39fF
C5535 a_13459_28111# a_18823_50247# 0.83fF
C5536 pmat.rowon_n[10] vcm 0.61fF
C5537 a_32687_46607# a_1781_9308# 0.65fF
C5538 a_22178_60146# vcm 0.62fF
C5539 pmat.en_bit_n[2] ANTENNA__1395__B1.DIODE 1.27fF
C5540 VDD a_27198_10496# 0.52fF
C5541 a_13091_28327# a_7415_29397# 0.50fF
C5542 VDD a_22357_39141# 1.26fF
C5543 a_40250_20536# ctopn 3.58fF
C5544 a_23182_15516# a_23182_14512# 1.00fF
C5545 a_47278_15516# a_48282_15516# 0.97fF
C5546 VDD a_9427_50095# 1.14fF
C5547 a_6927_30503# a_5363_33551# 0.34fF
C5548 a_18546_58180# a_34134_58138# 0.35fF
C5549 a_25190_69182# a_25190_68178# 1.00fF
C5550 a_46274_69182# a_47278_69182# 0.97fF
C5551 a_6559_33767# a_7163_53333# 0.40fF
C5552 a_18546_10494# a_34134_10902# 0.35fF
C5553 _1196_.B1 ANTENNA__1190__A1.DIODE 1.69fF
C5554 a_33222_21540# a_33222_20536# 1.00fF
C5555 VDD a_20811_34743# 0.59fF
C5556 a_24591_28327# pmat.col[14] 0.79fF
C5557 a_18546_10494# vcm 0.40fF
C5558 a_34226_62154# ctopp 3.58fF
C5559 _1183_.A2 nmat.col[26] 3.65fF
C5560 VDD a_43262_62154# 0.52fF
C5561 a_28202_16520# vcm 0.65fF
C5562 a_11149_40188# a_12197_43746# 0.45fF
C5563 VDD a_8267_49159# 0.54fF
C5564 pmat.col[27] vcm 5.88fF
C5565 a_8569_60405# a_8841_60405# 0.41fF
C5566 VDD a_19413_40229# 1.23fF
C5567 VDD a_45325_38127# 0.71fF
C5568 a_4337_22351# clk_dig 0.34fF
C5569 a_6787_47607# a_10497_54697# 0.40fF
C5570 VDD a_5331_13951# 0.34fF
C5571 VDD config_2_in[2] 0.57fF
C5572 a_6927_30503# a_11202_55687# 0.82fF
C5573 a_33222_70186# ctopp 3.57fF
C5574 VDD a_1591_54991# 1.62fF
C5575 a_10239_77295# a_11023_76359# 0.30fF
C5576 VDD a_42258_70186# 0.52fF
C5577 a_29206_15516# ctopn 3.58fF
C5578 VDD a_29206_11500# 0.52fF
C5579 a_28202_23548# m2_27972_24282# 0.99fF
C5580 a_5351_19913# a_4523_21276# 2.59fF
C5581 a_18546_72236# a_43170_72194# 0.35fF
C5582 a_44266_23548# a_44266_22544# 1.00fF
C5583 VDD a_4313_44111# 0.62fF
C5584 VDD nmat.col[29] 12.07fF
C5585 ANTENNA__1195__A1.DIODE a_26891_28327# 2.96fF
C5586 a_19166_60146# a_19166_59142# 1.00fF
C5587 a_43262_60146# a_44266_60146# 0.97fF
C5588 a_48282_12504# ctopn 3.58fF
C5589 a_18546_69224# a_29114_69182# 0.35fF
C5590 pmat.col_n[3] ctopp 2.02fF
C5591 a_27198_11500# a_27198_10496# 1.00fF
C5592 a_44266_56130# vcm 0.62fF
C5593 VDD a_36617_36603# 1.36fF
C5594 VDD a_29114_72194# 0.32fF
C5595 VDD a_4383_7093# 15.42fF
C5596 a_18546_63200# a_48190_63158# 0.35fF
C5597 VDD m2_17932_69002# 1.12fF
C5598 a_20475_49783# a_11948_49783# 0.45fF
C5599 a_26194_22544# vcm 0.65fF
C5600 a_32218_61150# a_33222_61150# 0.97fF
C5601 a_24186_68178# ctopp 3.58fF
C5602 a_47278_66170# vcm 0.62fF
C5603 VDD a_33222_68178# 0.52fF
C5604 nmat.en_bit_n[2] nmat.col_n[16] 0.30fF
C5605 ANTENNA__1395__A1.DIODE inn_analog 15.94fF
C5606 nmat.col[28] ANTENNA__1190__A2.DIODE 13.09fF
C5607 VDD a_40591_43447# 0.70fF
C5608 a_4075_13653# a_4241_13653# 0.72fF
C5609 a_40250_63158# vcm 0.62fF
C5610 a_5363_70543# a_11508_48187# 0.59fF
C5611 a_38905_28853# a_28704_29568# 0.33fF
C5612 pmat.col_n[1] a_18823_50247# 0.31fF
C5613 VDD a_33101_29673# 0.64fF
C5614 a_6927_30503# nmat.col_n[12] 0.69fF
C5615 a_1923_53055# a_1823_58237# 0.48fF
C5616 a_10515_15055# a_11067_64015# 1.15fF
C5617 ANTENNA__1195__A1.DIODE _1184_.A2 9.07fF
C5618 pmat.sample a_19541_28879# 0.43fF
C5619 a_2149_45717# a_5497_73719# 0.59fF
C5620 a_18546_20534# a_35138_20942# 0.35fF
C5621 a_26194_20536# a_27198_20536# 0.97fF
C5622 a_31214_16520# ctopn 3.58fF
C5623 VDD result_out[12] 0.54fF
C5624 a_8491_47911# a_13605_71017# 0.45fF
C5625 VDD m2_17932_8218# 1.03fF
C5626 a_13459_28111# a_35244_32411# 0.52fF
C5627 VDD a_6795_76989# 1.97fF
C5628 a_49286_16520# a_50290_16520# 0.97fF
C5629 VDD a_38391_48469# 0.38fF
C5630 a_39246_67174# a_39246_66170# 1.00fF
C5631 a_25190_9492# a_25190_8488# 1.00fF
C5632 _1192_.B1 nmat.col[7] 0.79fF
C5633 VDD a_38242_23548# 0.55fF
C5634 m2_17932_21270# m2_17932_20266# 0.99fF
C5635 VDD a_12993_66415# 0.45fF
C5636 VDD a_40250_9492# 0.52fF
C5637 a_18546_11498# a_38150_11906# 0.35fF
C5638 VDD a_19423_37737# 0.57fF
C5639 a_28704_29568# ANTENNA__1183__B1.DIODE 0.87fF
C5640 a_38242_17524# a_39246_17524# 0.97fF
C5641 a_36234_57134# a_37238_57134# 0.97fF
C5642 pmat.rowon_n[2] vcm 0.60fF
C5643 a_1899_35051# a_5221_45199# 0.59fF
C5644 a_41254_20536# a_41254_19532# 1.00fF
C5645 _1224_.X _1194_.A2 0.88fF
C5646 a_35230_71190# a_36234_71190# 0.97fF
C5647 a_45270_67174# vcm 0.62fF
C5648 VDD a_14249_49525# 0.63fF
C5649 a_22178_58138# a_23182_58138# 0.97fF
C5650 a_34226_14512# vcm 0.65fF
C5651 VDD a_14457_15823# 0.91fF
C5652 a_33222_64162# vcm 0.62fF
C5653 pmat.col_n[3] m2_21948_54946# 0.38fF
C5654 a_7939_31591# a_9963_28111# 6.82fF
C5655 a_39246_8488# a_40250_8488# 0.97fF
C5656 VDD a_37143_31573# 0.64fF
C5657 pmat.rowoff_n[15] nmat.rowoff_n[0] 20.39fF
C5658 VDD _1187_.A2 20.19fF
C5659 a_14600_37607# a_26767_34967# 0.44fF
C5660 VDD a_16837_35515# 1.24fF
C5661 VDD a_36234_13508# 0.52fF
C5662 cgen.dlycontrol3_in[4] cgen.dlycontrol1_in[4] 0.55fF
C5663 a_47278_14512# a_47278_13508# 1.00fF
C5664 a_4351_55527# a_5535_57993# 1.03fF
C5665 a_29206_22544# ctopn 3.57fF
C5666 nmat.col_n[30] vcm 6.70fF
C5667 VDD a_34226_18528# 0.52fF
C5668 pmat.sw nmat.col[10] 0.79fF
C5669 nmat.rowon_n[14] cgen.dlycontrol4_in[3] 0.50fF
C5670 a_22178_61150# a_22178_60146# 1.00fF
C5671 a_30210_19532# a_30210_18528# 1.00fF
C5672 a_11116_18695# a_4383_7093# 0.31fF
C5673 a_16311_28327# a_20439_27247# 3.62fF
C5674 a_7415_29397# a_11927_27399# 0.36fF
C5675 VDD a_45270_15516# 0.52fF
C5676 a_1591_40853# a_2411_33749# 0.34fF
C5677 a_18546_14510# a_36142_14918# 0.35fF
C5678 m2_51064_15246# vcm 0.55fF
C5679 _1154_.X a_22199_30287# 2.45fF
C5680 a_18546_64204# a_34134_64162# 0.35fF
C5681 a_2835_13077# a_12539_10389# 0.34fF
C5682 a_13432_62581# a_12044_49641# 0.45fF
C5683 a_23182_59142# a_23182_58138# 1.00fF
C5684 pmat.rowoff_n[15] a_5363_33551# 1.34fF
C5685 a_25879_31591# a_10883_3303# 0.51fF
C5686 VDD a_5070_26703# 0.47fF
C5687 a_1781_9308# a_1979_9334# 0.30fF
C5688 VDD a_2124_74299# 0.70fF
C5689 a_36234_65166# vcm 0.62fF
C5690 cgen.dlycontrol3_in[1] a_11113_40835# 1.99fF
C5691 a_43262_21540# vcm 0.65fF
C5692 a_5535_57993# a_10090_58093# 0.34fF
C5693 a_32218_60146# ctopp 3.58fF
C5694 a_11711_50959# a_21279_48999# 0.39fF
C5695 VDD a_41254_60146# 0.52fF
C5696 a_10239_14183# a_3305_17999# 0.59fF
C5697 VDD a_33765_36965# 1.14fF
C5698 a_11497_38543# ndecision_finish 1.40fF
C5699 VDD a_4259_31375# 4.71fF
C5700 a_19166_14512# m2_17932_14242# 0.96fF
C5701 pmat.row_n[6] a_18546_62196# 0.35fF
C5702 a_28202_17524# a_28202_16520# 1.00fF
C5703 a_24407_31375# nmat.col_n[19] 0.74fF
C5704 a_18546_19530# a_47186_19938# 0.35fF
C5705 a_37238_14512# ctopn 3.58fF
C5706 VDD a_7435_68021# 0.62fF
C5707 a_8491_47911# a_13091_54447# 0.46fF
C5708 a_18546_12502# a_51202_12910# 0.35fF
C5709 a_34226_12504# a_35230_12504# 0.97fF
C5710 a_47278_22544# a_48282_22544# 0.97fF
C5711 VDD a_47278_16520# 0.52fF
C5712 a_11041_40948# a_12116_40871# 2.52fF
C5713 a_6292_69831# a_4075_50087# 0.32fF
C5714 a_23182_59142# a_24186_59142# 0.97fF
C5715 a_18546_59184# a_29114_59142# 0.35fF
C5716 a_25190_57134# ctopp 3.57fF
C5717 VDD a_20591_31029# 0.44fF
C5718 VDD a_8703_6202# 1.13fF
C5719 a_24186_71190# ctopp 3.40fF
C5720 a_2149_45717# a_1739_47893# 0.38fF
C5721 VDD a_34226_57134# 0.52fF
C5722 a_4719_30287# a_4259_31375# 0.42fF
C5723 a_50290_69182# vcm 0.62fF
C5724 VDD a_33222_71190# 0.55fF
C5725 VDD a_20170_58138# 0.52fF
C5726 a_31214_71190# m2_30984_72014# 1.00fF
C5727 VDD a_20170_23548# 0.54fF
C5728 a_10055_31591# a_5179_31591# 0.41fF
C5729 cgen.dlycontrol4_in[2] cgen.dlycontrol1_in[2] 0.48fF
C5730 a_11021_42619# a_11297_36091# 0.57fF
C5731 VDD a_46753_41935# 1.26fF
C5732 a_18546_55168# a_45178_55126# 0.35fF
C5733 a_18546_24550# a_34134_24958# 0.39fF
C5734 a_13091_52047# a_13643_29415# 0.59fF
C5735 VDD a_5233_40553# 0.42fF
C5736 a_16311_28327# a_27763_27221# 1.43fF
C5737 VDD pmat.col[1] 5.55fF
C5738 VDD a_4243_54991# 0.40fF
C5739 a_30571_50959# ANTENNA__1183__B1.DIODE 0.33fF
C5740 a_36234_61150# vcm 0.62fF
C5741 a_30819_40191# a_29163_38545# 0.39fF
C5742 a_18546_22542# a_31122_22950# 0.35fF
C5743 a_46274_21540# ctopn 3.58fF
C5744 VDD a_9075_28023# 2.19fF
C5745 a_30210_20536# vcm 0.65fF
C5746 VDD a_45270_22544# 0.52fF
C5747 m2_17932_70006# m3_18064_70138# 2.76fF
C5748 _1154_.X nmat.col_n[30] 1.09fF
C5749 a_4991_69831# a_10878_58487# 1.65fF
C5750 VDD a_21174_59142# 0.52fF
C5751 a_50290_63158# ctopp 3.43fF
C5752 VDD a_4927_50613# 0.38fF
C5753 ANTENNA__1190__A1.DIODE a_45019_38645# 0.62fF
C5754 a_42258_17524# vcm 0.65fF
C5755 pmat.en_bit_n[2] nmat.col[18] 1.04fF
C5756 pmat.row_n[7] a_2191_25045# 0.43fF
C5757 pmat.rowoff_n[12] pmat.rowoff_n[5] 0.64fF
C5758 m2_30984_24282# m2_31988_24282# 0.96fF
C5759 a_43262_8488# vcm 0.64fF
C5760 pmat.row_n[0] nmat.col[7] 0.81fF
C5761 a_12197_38306# a_19233_38215# 0.34fF
C5762 VDD pmat.col[4] 4.45fF
C5763 VDD a_16689_43132# 1.12fF
C5764 m2_25964_7214# m2_26968_7214# 0.96fF
C5765 a_5687_38279# a_4533_38279# 0.52fF
C5766 ANTENNA__1195__A1.DIODE nmat.col_n[27] 0.76fF
C5767 pmat.col_n[8] a_24407_31375# 0.36fF
C5768 VDD a_9323_28879# 0.37fF
C5769 a_50290_18528# a_50290_17524# 1.00fF
C5770 a_10515_75895# a_10697_75218# 1.20fF
C5771 pmat.row_n[15] nmat.sample 0.33fF
C5772 VDD a_2944_69928# 0.48fF
C5773 VDD a_2564_21959# 5.41fF
C5774 a_2407_49289# a_5053_59575# 0.41fF
C5775 pmat.row_n[12] a_10055_31591# 1.01fF
C5776 VDD nmat.col_n[11] 5.28fF
C5777 a_18162_15516# vcm 6.95fF
C5778 a_12228_40693# a_22361_41479# 0.61fF
C5779 a_50290_63158# a_50290_62154# 1.00fF
C5780 a_18546_65208# vcm 0.40fF
C5781 a_50290_71190# m2_50060_72014# 1.00fF
C5782 a_10515_15055# a_3571_13627# 0.50fF
C5783 pmat.col_n[13] a_24591_28327# 0.35fF
C5784 pmat.rowon_n[7] a_4128_64391# 0.84fF
C5785 a_18546_18526# a_48190_18934# 0.35fF
C5786 a_26194_70186# a_26194_69182# 1.00fF
C5787 a_2021_11043# a_3663_9269# 0.31fF
C5788 a_2411_43301# cgen.dlycontrol4_in[2] 0.43fF
C5789 a_38242_12504# vcm 0.65fF
C5790 a_43262_64162# ctopp 3.58fF
C5791 a_6664_26159# a_25315_28335# 0.41fF
C5792 m2_49056_7214# m3_49188_7346# 2.79fF
C5793 a_35230_24552# a_36234_24552# 0.97fF
C5794 VDD a_21174_19532# 0.52fF
C5795 m2_26968_54946# m3_27100_55078# 2.79fF
C5796 a_3923_68021# a_12217_66389# 0.55fF
C5797 ANTENNA_fanout52_A.DIODE _1192_.A2 0.83fF
C5798 a_18243_28327# a_21739_29415# 0.43fF
C5799 a_23182_19532# a_24186_19532# 0.97fF
C5800 a_17842_27497# nmat.col_n[19] 2.93fF
C5801 a_18243_28327# a_20310_28029# 0.52fF
C5802 a_49286_13508# a_49286_12504# 1.00fF
C5803 a_1586_18231# a_2411_16101# 0.93fF
C5804 a_11067_27239# nmat.col[12] 1.13fF
C5805 a_10772_77563# a_10811_77437# 0.79fF
C5806 VDD a_1591_38677# 0.43fF
C5807 a_33222_20536# ctopn 3.58fF
C5808 VDD a_10927_43421# 1.19fF
C5809 a_19166_15516# a_19166_14512# 1.00fF
C5810 a_4707_32156# a_14453_31599# 0.77fF
C5811 a_23933_32143# a_24374_29941# 0.39fF
C5812 m2_17932_66994# m3_18064_67126# 2.76fF
C5813 a_18546_58180# a_27106_58138# 0.35fF
C5814 a_22178_10496# a_23182_10496# 0.97fF
C5815 a_18546_10494# a_27106_10902# 0.35fF
C5816 VDD a_4792_34435# 0.65fF
C5817 a_45270_17524# ctopn 3.58fF
C5818 VDD a_5081_53135# 6.40fF
C5819 pmat.rowon_n[3] cgen.dlycontrol3_in[4] 1.07fF
C5820 a_27198_62154# ctopp 3.58fF
C5821 pmat.col_n[5] pmat.col[5] 0.98fF
C5822 VDD a_36234_62154# 0.52fF
C5823 a_21174_16520# vcm 0.65fF
C5824 a_19166_71190# m2_18936_72014# 1.00fF
C5825 m2_40020_24282# vcm 0.42fF
C5826 a_46274_8488# ctopn 3.40fF
C5827 a_11041_38772# a_11149_36924# 0.68fF
C5828 a_18546_56172# a_49194_56130# 0.35fF
C5829 a_33222_56130# a_34226_56130# 0.97fF
C5830 VDD a_48190_24958# 0.44fF
C5831 a_46274_65166# ctopp 3.58fF
C5832 VDD a_33617_42333# 1.12fF
C5833 ANTENNA__1190__B1.DIODE a_7109_29423# 0.36fF
C5834 ANTENNA__1197__A.DIODE a_16311_28327# 0.66fF
C5835 a_18546_55168# a_28110_55126# 0.35fF
C5836 nmat.col[24] nmat.col[21] 1.39fF
C5837 pmat.en_bit_n[2] a_23395_53135# 1.21fF
C5838 ANTENNA__1197__B.DIODE a_25695_28111# 1.12fF
C5839 VDD a_24131_29967# 0.31fF
C5840 a_26194_70186# ctopp 3.57fF
C5841 pmat.rowon_n[0] a_5173_9839# 0.35fF
C5842 VDD a_35230_70186# 0.52fF
C5843 a_22178_15516# ctopn 3.58fF
C5844 a_18546_61192# vcm 0.40fF
C5845 VDD a_22178_11500# 0.52fF
C5846 pmat.col[7] ctopp 1.97fF
C5847 ANTENNA__1183__B1.DIODE nmat.col_n[1] 0.48fF
C5848 a_38242_62154# a_39246_62154# 0.97fF
C5849 a_45270_16520# a_45270_15516# 1.00fF
C5850 a_36234_66170# a_37238_66170# 0.97fF
C5851 m2_41024_72014# m3_41156_72146# 2.79fF
C5852 a_41254_12504# ctopn 3.58fF
C5853 a_18546_69224# a_22086_69182# 0.35fF
C5854 a_37238_56130# vcm 0.62fF
C5855 a_12851_28853# a_12461_29673# 1.08fF
C5856 a_25695_28111# a_31675_47695# 0.70fF
C5857 a_29206_63158# a_30210_63158# 0.97fF
C5858 a_18546_63200# a_41162_63158# 0.35fF
C5859 pmat.row_n[11] nmat.rowoff_n[3] 0.80fF
C5860 cgen.dlycontrol3_in[1] cgen.dlycontrol4_in[4] 1.22fF
C5861 VDD a_6173_22895# 1.19fF
C5862 a_40250_66170# vcm 0.62fF
C5863 VDD a_26194_68178# 0.52fF
C5864 m2_50060_72014# m2_51064_72014# 0.96fF
C5865 VDD a_28981_43493# 1.36fF
C5866 ANTENNA__1184__B1.DIODE a_24747_29967# 0.51fF
C5867 a_33222_63158# vcm 0.62fF
C5868 ANTENNA__1190__A1.DIODE nmat.sw 0.35fF
C5869 VDD a_47212_29673# 0.64fF
C5870 nmat.sample nmat.sample_n 11.16fF
C5871 m2_17932_63982# m3_18064_64114# 2.76fF
C5872 VDD a_47186_55126# 0.42fF
C5873 VDD a_33515_31055# 1.10fF
C5874 pmat.row_n[13] a_10515_13967# 0.48fF
C5875 VDD m2_51064_18258# 1.01fF
C5876 a_18546_20534# a_28110_20942# 0.35fF
C5877 a_24186_16520# ctopn 3.58fF
C5878 a_13091_18535# a_9441_20189# 0.89fF
C5879 a_10515_13967# cgen.enable_dlycontrol_in 3.80fF
C5880 nmat.rowon_n[1] nmat.rowoff_n[3] 2.52fF
C5881 a_2263_43719# a_11948_49783# 0.38fF
C5882 pmat.col_n[10] pmat.col[11] 6.00fF
C5883 VDD a_13275_48783# 14.21fF
C5884 VDD a_31214_23548# 0.55fF
C5885 a_46274_61150# ctopp 3.58fF
C5886 a_37238_70186# a_38242_70186# 0.97fF
C5887 VDD a_33222_9492# 0.52fF
C5888 a_24186_11500# a_25190_11500# 0.97fF
C5889 a_18546_11498# a_31122_11906# 0.35fF
C5890 a_2263_43719# a_30571_50959# 0.63fF
C5891 pmat.rowoff_n[4] a_11067_16359# 0.43fF
C5892 a_20170_12504# vcm 0.65fF
C5893 VDD a_26515_41271# 0.60fF
C5894 a_13459_28111# a_21371_50087# 1.65fF
C5895 VDD a_49286_20536# 0.52fF
C5896 a_26194_64162# a_26194_63158# 1.00fF
C5897 pmat.row_n[4] a_3325_20175# 0.65fF
C5898 a_29206_10496# a_29206_9492# 1.00fF
C5899 a_18546_71232# a_46182_71190# 0.35fF
C5900 a_38242_67174# vcm 0.62fF
C5901 a_26194_58138# a_26194_57134# 1.00fF
C5902 VDD a_1757_50095# 0.62fF
C5903 a_27198_14512# vcm 0.65fF
C5904 cgen.dlycontrol4_in[1] a_2411_33749# 0.76fF
C5905 pmat.col_n[28] pmat.col[28] 0.97fF
C5906 a_10441_21263# a_10513_24135# 1.01fF
C5907 a_26194_64162# vcm 0.62fF
C5908 VDD m2_18936_24282# 0.65fF
C5909 a_22199_30287# a_21365_27247# 0.39fF
C5910 a_30210_60146# a_30210_59142# 1.00fF
C5911 a_18546_65208# a_51202_65166# 0.35fF
C5912 VDD a_10985_35516# 1.27fF
C5913 a_48282_62154# a_48282_61150# 1.00fF
C5914 VDD a_29206_13508# 0.52fF
C5915 a_28812_29575# nmat.col[30] 0.60fF
C5916 VDD a_18546_62196# 32.63fF
C5917 a_18546_23546# a_20078_23954# 0.35fF
C5918 a_19166_66170# m2_17932_65990# 0.96fF
C5919 a_22178_22544# ctopn 3.57fF
C5920 VDD a_27198_18528# 0.52fF
C5921 a_24186_63158# pmat.col[5] 0.31fF
C5922 a_12309_38659# a_22153_37179# 0.30fF
C5923 a_18546_67216# a_51202_67174# 0.35fF
C5924 a_34226_67174# a_35230_67174# 0.97fF
C5925 m2_17932_70006# m2_17932_69002# 0.99fF
C5926 a_31214_66170# a_31214_65166# 1.00fF
C5927 a_24186_22544# a_24186_21540# 1.00fF
C5928 VDD a_38242_15516# 0.52fF
C5929 a_7717_14735# a_7644_16341# 0.97fF
C5930 a_48282_15516# a_48282_14512# 1.00fF
C5931 a_23182_14512# a_24186_14512# 0.97fF
C5932 a_18546_14510# a_29114_14918# 0.35fF
C5933 pmat.rowoff_n[4] vcm 0.81fF
C5934 pmat.sw ANTENNA__1395__A2.DIODE 0.35fF
C5935 a_18546_18526# vcm 0.40fF
C5936 a_18546_7482# a_51202_7890# 0.35fF
C5937 a_18546_64204# a_27106_64162# 0.35fF
C5938 a_22178_64162# a_23182_64162# 0.97fF
C5939 m2_17932_60970# m3_18064_61102# 2.76fF
C5940 pmat.col_n[17] a_36234_55126# 0.31fF
C5941 a_32319_50345# a_28915_50959# 0.35fF
C5942 a_28202_68178# a_29206_68178# 0.97fF
C5943 a_18546_56172# ctopp 1.36fF
C5944 a_50290_69182# a_50290_68178# 1.00fF
C5945 a_1674_68047# a_3175_72641# 0.57fF
C5946 a_1923_69823# a_8491_47911# 0.45fF
C5947 a_2149_45717# a_1899_35051# 2.55fF
C5948 pmat.col_n[14] pmat.col[15] 6.66fF
C5949 a_12069_36341# clk_ena 3.10fF
C5950 a_21174_8488# m2_20944_7214# 1.00fF
C5951 nmat.col[8] ctopn 1.97fF
C5952 VDD a_8479_11484# 0.54fF
C5953 a_14287_69455# a_11067_64015# 2.38fF
C5954 VDD m2_43032_7214# 1.32fF
C5955 a_6817_21807# a_3305_15823# 0.39fF
C5956 a_10071_17999# a_8197_20871# 0.32fF
C5957 pmat.col_n[5] a_18243_28327# 0.31fF
C5958 a_10781_42869# a_13227_42333# 0.30fF
C5959 a_3339_70759# a_2215_47375# 1.48fF
C5960 a_2149_45717# a_2419_53351# 0.64fF
C5961 a_29206_65166# vcm 0.62fF
C5962 nmat.col_n[3] vcm 2.80fF
C5963 a_36234_21540# vcm 0.65fF
C5964 a_25190_60146# ctopp 3.58fF
C5965 a_5497_62839# a_4985_51433# 2.86fF
C5966 VDD a_34226_60146# 0.52fF
C5967 a_32405_32463# a_34243_32143# 0.37fF
C5968 ANTENNA__1190__A1.DIODE a_22199_30287# 2.45fF
C5969 a_12237_36596# a_14773_37218# 0.98fF
C5970 nmat.col_n[18] nmat.col[18] 0.78fF
C5971 VDD a_2124_72123# 0.66fF
C5972 _1192_.A2 nmat.col_n[29] 4.32fF
C5973 a_18546_19530# a_40158_19938# 0.35fF
C5974 m2_26968_54946# m2_27972_54946# 0.96fF
C5975 pmat.col_n[30] pmat.col[31] 6.17fF
C5976 a_30210_14512# ctopn 3.58fF
C5977 a_7717_14735# a_8767_16055# 0.42fF
C5978 a_18546_12502# a_44174_12910# 0.35fF
C5979 a_1591_71855# a_1674_57711# 0.99fF
C5980 _1194_.B1 nmat.col_n[3] 1.13fF
C5981 VDD a_27603_34191# 2.52fF
C5982 VDD a_34611_44265# 0.64fF
C5983 VDD a_40250_16520# 0.52fF
C5984 m2_17932_9222# m2_17932_8218# 0.99fF
C5985 a_18546_59184# a_22086_59142# 0.35fF
C5986 a_24186_65166# a_24186_64162# 1.00fF
C5987 pmat.sample_n a_13275_48783# 0.77fF
C5988 a_30571_50959# a_40105_47375# 0.64fF
C5989 VDD a_30118_55126# 0.42fF
C5990 VDD a_12245_31061# 0.63fF
C5991 VDD a_50198_7890# 0.33fF
C5992 VDD a_12792_58633# 0.32fF
C5993 VDD a_27198_57134# 0.52fF
C5994 VDD a_46522_34293# 0.60fF
C5995 a_43262_69182# vcm 0.62fF
C5996 VDD a_26194_71190# 0.55fF
C5997 a_10239_14183# a_9963_13967# 2.02fF
C5998 a_33222_23548# a_34226_23548# 0.97fF
C5999 a_18546_23546# a_49194_23954# 0.35fF
C6000 VDD a_25850_48981# 1.13fF
C6001 _1194_.A2 ANTENNA__1183__B1.DIODE 1.25fF
C6002 a_35230_9492# a_36234_9492# 0.97fF
C6003 a_42258_12504# a_42258_11500# 1.00fF
C6004 a_18162_57174# vcm 6.95fF
C6005 VDD a_13837_37981# 1.27fF
C6006 a_32405_32463# a_35244_32411# 0.32fF
C6007 VDD a_10767_39087# 1.89fF
C6008 a_4351_55527# a_2315_44124# 1.07fF
C6009 a_18546_55168# a_38150_55126# 0.35fF
C6010 a_18546_24550# a_27106_24958# 0.35fF
C6011 m2_17932_57958# m3_18064_58090# 2.76fF
C6012 a_47278_56130# ctopp 3.40fF
C6013 pmat.col[31] ctopp 3.45fF
C6014 a_1674_68047# a_1823_74557# 0.30fF
C6015 a_40250_8488# m2_40020_7214# 1.00fF
C6016 a_29206_61150# vcm 0.62fF
C6017 a_20170_23548# m2_18936_23278# 0.96fF
C6018 a_18546_72236# a_46182_72194# 0.35fF
C6019 a_18546_22542# a_24094_22950# 0.35fF
C6020 a_39246_21540# ctopn 3.58fF
C6021 nmat.rowon_n[10] vcm 0.53fF
C6022 pmat.col_n[17] pmat.col[17] 0.64fF
C6023 a_23182_20536# vcm 0.65fF
C6024 a_50290_9492# a_50290_8488# 1.00fF
C6025 nmat.sw a_11317_36924# 0.33fF
C6026 VDD a_38242_22544# 0.52fF
C6027 a_25190_65166# a_26194_65166# 0.97fF
C6028 a_50290_66170# ctopp 3.43fF
C6029 VDD a_23933_32143# 1.50fF
C6030 pmat.col_n[6] ctopp 2.02fF
C6031 a_10873_36341# cgen.dlycontrol1_in[4] 3.16fF
C6032 a_32218_21540# a_33222_21540# 0.97fF
C6033 pmat.rowon_n[8] a_4075_31591# 0.38fF
C6034 a_3305_15823# a_4383_7093# 0.35fF
C6035 pmat.rowoff_n[15] pmat.row_n[4] 3.42fF
C6036 VDD a_32126_72194# 0.32fF
C6037 a_41731_49525# a_45370_48169# 0.36fF
C6038 a_43262_63158# ctopp 3.58fF
C6039 a_17702_29967# a_16478_29423# 0.62fF
C6040 _1194_.B1 a_41731_49525# 0.69fF
C6041 nmat.col[1] vcm 5.76fF
C6042 VDD a_1644_62581# 0.30fF
C6043 a_35230_17524# vcm 0.65fF
C6044 a_14712_37429# ndecision_finish 0.72fF
C6045 m2_51064_56954# vcm 0.52fF
C6046 a_18546_61192# a_51202_61150# 0.35fF
C6047 VDD a_8291_23983# 0.66fF
C6048 m2_23956_24282# m2_24960_24282# 0.96fF
C6049 a_33222_71190# a_33222_70186# 1.00fF
C6050 a_36234_8488# vcm 0.64fF
C6051 pmat.col[18] m2_37008_54946# 0.41fF
C6052 a_27763_27221# nmat.col_n[26] 0.43fF
C6053 nmat.col_n[12] a_5991_23983# 1.81fF
C6054 m2_17932_17254# a_19166_17524# 0.96fF
C6055 a_50290_62154# pmat.col[31] 0.31fF
C6056 a_47278_58138# a_48282_58138# 0.97fF
C6057 VDD a_10949_43124# 2.07fF
C6058 pmat.rowon_n[3] a_13091_18535# 0.86fF
C6059 VDD a_20170_15516# 0.52fF
C6060 a_1823_74557# a_1923_61759# 0.39fF
C6061 m2_18936_7214# m2_19940_7214# 0.96fF
C6062 VDD nmat.col[30] 11.34fF
C6063 ANTENNA__1395__B1.DIODE a_15667_27239# 0.86fF
C6064 a_19166_68178# a_20170_68178# 0.97fF
C6065 a_6292_69831# a_7092_74005# 0.62fF
C6066 a_5823_34863# a_5989_34863# 0.66fF
C6067 cgen.dlycontrol1_in[4] cgen.dlycontrol1_in[3] 1.34fF
C6068 a_1899_35051# cgen.dlycontrol3_in[3] 0.73fF
C6069 VDD a_8013_56085# 0.57fF
C6070 a_2564_21959# a_4523_21276# 0.46fF
C6071 VDD a_2387_70483# 0.52fF
C6072 a_31214_13508# a_32218_13508# 0.97fF
C6073 a_18546_13506# a_45178_13914# 0.35fF
C6074 pmat.rowoff_n[12] a_8305_20871# 0.62fF
C6075 a_20310_28029# nmat.col_n[1] 0.34fF
C6076 VDD a_8031_76757# 0.50fF
C6077 a_14691_27399# a_12987_26159# 0.89fF
C6078 a_22153_37179# cgen.dlycontrol1_in[4] 2.55fF
C6079 _1224_.X ANTENNA__1197__B.DIODE 4.01fF
C6080 a_47278_61150# a_47278_60146# 1.00fF
C6081 a_48282_67174# ctopp 3.58fF
C6082 a_18546_18526# a_41162_18934# 0.35fF
C6083 a_29206_18528# a_30210_18528# 0.97fF
C6084 a_11149_36924# a_11317_36924# 1.81fF
C6085 a_24407_31375# a_16478_29423# 0.38fF
C6086 a_10055_31591# a_11948_49783# 1.10fF
C6087 a_31214_12504# vcm 0.65fF
C6088 a_36234_64162# ctopp 3.58fF
C6089 a_15101_29423# a_14691_29575# 0.30fF
C6090 a_14917_23983# a_10589_22351# 0.31fF
C6091 VDD a_46274_14512# 0.52fF
C6092 a_10055_31591# a_2046_30184# 1.47fF
C6093 VDD a_45270_64162# 0.52fF
C6094 a_47147_44655# a_47290_45717# 0.49fF
C6095 cgen.enable_dlycontrol_in a_10873_39605# 0.32fF
C6096 nmat.col_n[28] nmat.col[24] 7.25fF
C6097 nmat.col_n[26] nmat.col[27] 6.51fF
C6098 a_48282_59142# a_48282_58138# 1.00fF
C6099 a_11067_30287# a_40741_46565# 0.30fF
C6100 VDD a_25695_28111# 12.74fF
C6101 a_50290_23548# m2_50060_24282# 0.99fF
C6102 a_12447_16143# ANTENNA__1196__A2.DIODE 0.72fF
C6103 a_26194_20536# ctopn 3.58fF
C6104 VDD a_34002_44527# 0.36fF
C6105 a_11389_40443# a_10873_40693# 4.47fF
C6106 inp_analog a_11067_27239# 0.39fF
C6107 a_40250_15516# a_41254_15516# 0.97fF
C6108 a_14839_20871# a_9963_28111# 0.56fF
C6109 VDD a_1781_9308# 25.73fF
C6110 pmat.sample_n a_25850_48981# 0.63fF
C6111 a_39246_69182# a_40250_69182# 0.97fF
C6112 pmat.col_n[0] ANTENNA__1190__B1.DIODE 1.18fF
C6113 a_18546_10494# a_19074_10902# 0.35fF
C6114 a_26194_21540# a_26194_20536# 1.00fF
C6115 a_24867_53135# a_18243_28327# 1.20fF
C6116 a_38242_17524# ctopn 3.58fF
C6117 a_20170_62154# ctopp 3.57fF
C6118 a_14641_57167# nmat.rowon_n[7] 1.30fF
C6119 a_1923_61759# a_7797_63151# 0.45fF
C6120 VDD a_29206_62154# 0.52fF
C6121 a_39246_8488# ctopn 3.40fF
C6122 a_18546_56172# a_42166_56130# 0.35fF
C6123 VDD a_41162_24958# 0.44fF
C6124 a_12309_38659# a_14712_37429# 1.00fF
C6125 VDD a_1823_66941# 3.66fF
C6126 m2_17932_18258# m3_18064_18390# 2.76fF
C6127 pmat.col_n[3] pmat.col[4] 6.54fF
C6128 a_39246_65166# ctopp 3.58fF
C6129 VDD a_48282_65166# 0.52fF
C6130 a_18546_55168# a_21082_55126# 0.35fF
C6131 a_48282_59142# a_49286_59142# 0.97fF
C6132 a_5462_62215# a_7457_62037# 0.59fF
C6133 VDD a_2219_4943# 0.45fF
C6134 a_18546_68220# a_50198_68178# 0.35fF
C6135 a_5363_33551# nmat.sample 0.34fF
C6136 a_2007_25597# clk_ena 0.80fF
C6137 pmat.col_n[22] pmat.col[23] 6.06fF
C6138 a_29076_48695# a_31105_46805# 0.30fF
C6139 VDD a_28202_70186# 0.52fF
C6140 a_10589_22351# a_9441_20189# 0.68fF
C6141 VDD a_1895_26372# 0.53fF
C6142 a_37238_23548# a_37238_22544# 1.00fF
C6143 a_33423_47695# a_7717_14735# 0.42fF
C6144 a_2879_57487# a_4520_60975# 0.38fF
C6145 VDD a_9831_74183# 0.69fF
C6146 VDD a_3793_47479# 0.47fF
C6147 a_36234_60146# a_37238_60146# 0.97fF
C6148 VDD a_20170_22544# 0.52fF
C6149 a_34226_12504# ctopn 3.58fF
C6150 a_30210_56130# vcm 0.62fF
C6151 a_18546_63200# a_34134_63158# 0.35fF
C6152 a_11619_16367# a_11785_16367# 0.62fF
C6153 ANTENNA__1197__A.DIODE nmat.col_n[26] 1.09fF
C6154 _1192_.A2 a_13145_26935# 0.37fF
C6155 m2_22952_24282# m3_23084_24414# 2.79fF
C6156 a_44266_68178# a_44266_67174# 1.00fF
C6157 a_25190_61150# a_26194_61150# 0.97fF
C6158 a_33222_66170# vcm 0.62fF
C6159 pmat.col_n[20] pmat.col[21] 6.10fF
C6160 m2_43032_72014# m2_44036_72014# 0.96fF
C6161 a_4351_55527# a_5320_57863# 0.30fF
C6162 a_26194_63158# vcm 0.62fF
C6163 nmat.rowoff_n[6] a_11091_26311# 0.52fF
C6164 a_14887_46377# clk_ena 2.88fF
C6165 VDD a_12155_20719# 0.34fF
C6166 VDD a_40158_55126# 0.42fF
C6167 pmat.row_n[15] a_18162_71230# 25.57fF
C6168 VDD a_10699_72943# 1.09fF
C6169 a_50290_66170# m2_51064_65990# 0.96fF
C6170 a_10873_39605# a_12069_38517# 0.54fF
C6171 a_42258_16520# a_43262_16520# 0.97fF
C6172 a_32218_67174# a_32218_66170# 1.00fF
C6173 a_11067_64015# a_17139_30503# 0.38fF
C6174 a_18546_61192# pmat.rowoff_n[5] 4.09fF
C6175 VDD a_24186_23548# 0.55fF
C6176 VDD a_39505_38780# 1.27fF
C6177 a_39246_61150# ctopp 3.58fF
C6178 a_20170_18528# a_21174_18528# 0.97fF
C6179 nmat.col[12] m2_30984_24282# 0.39fF
C6180 VDD a_26194_9492# 0.52fF
C6181 VDD a_48282_61150# 0.52fF
C6182 a_18546_11498# a_24094_11906# 0.35fF
C6183 ANTENNA__1190__B1.DIODE nmat.col_n[10] 6.31fF
C6184 a_35230_24552# ctopn 1.70fF
C6185 VDD a_42258_20536# 0.52fF
C6186 a_31214_17524# a_32218_17524# 0.97fF
C6187 a_4399_51157# a_2659_35015# 0.80fF
C6188 a_29206_57134# a_30210_57134# 0.97fF
C6189 ANTENNA__1190__B1.DIODE clk_ena 0.45fF
C6190 cgen.dlycontrol1_in[0] a_1923_31743# 0.39fF
C6191 a_34226_20536# a_34226_19532# 1.00fF
C6192 a_31214_67174# vcm 0.62fF
C6193 a_18546_71232# a_39154_71190# 0.35fF
C6194 a_28202_71190# a_29206_71190# 0.97fF
C6195 VDD a_12431_69367# 0.49fF
C6196 a_13091_28327# a_15435_29111# 0.41fF
C6197 ANTENNA__1395__A1.DIODE a_13459_28111# 0.67fF
C6198 VDD a_6141_44629# 0.36fF
C6199 pmat.col_n[29] ANTENNA__1395__B1.DIODE 0.48fF
C6200 cgen.dlycontrol2_in[4] cgen.dlycontrol2_in[3] 1.41fF
C6201 VDD a_4979_38127# 1.24fF
C6202 VDD a_3199_53877# 0.51fF
C6203 a_32218_8488# a_33222_8488# 0.97fF
C6204 a_18546_8486# a_47186_8894# 0.35fF
C6205 a_18546_65208# a_44174_65166# 0.35fF
C6206 nmat.col_n[3] nmat.col_n[7] 0.98fF
C6207 pmat.sample pmat.row_n[10] 0.56fF
C6208 VDD a_28245_35877# 1.39fF
C6209 a_20170_17524# ctopn 3.57fF
C6210 VDD a_22178_13508# 0.52fF
C6211 a_40250_14512# a_40250_13508# 1.00fF
C6212 VDD a_21395_50857# 0.49fF
C6213 ANTENNA__1197__A.DIODE a_24407_31375# 0.32fF
C6214 _1194_.A2 a_21739_29415# 0.38fF
C6215 a_18546_67216# a_44174_67174# 0.35fF
C6216 a_44266_57134# a_44266_56130# 1.00fF
C6217 _1192_.A2 a_11927_27399# 0.63fF
C6218 a_48282_19532# a_49286_19532# 0.97fF
C6219 a_23182_19532# a_23182_18528# 1.00fF
C6220 a_36234_55126# m3_36136_55078# 2.45fF
C6221 m2_18936_24282# m2_18936_23278# 0.99fF
C6222 pmat.row_n[14] pmat.rowon_n[14] 20.33fF
C6223 VDD a_12987_26159# 1.22fF
C6224 a_7521_47081# a_10515_15055# 0.85fF
C6225 a_4075_68583# a_4025_54965# 0.72fF
C6226 VDD a_31214_15516# 0.52fF
C6227 pmat.rowoff_n[7] a_2467_35925# 0.54fF
C6228 a_18546_14510# a_22086_14918# 0.35fF
C6229 pmat.col[10] vcm 5.88fF
C6230 a_18546_7482# a_44174_7890# 0.35fF
C6231 a_5363_33551# a_5535_29980# 0.60fF
C6232 a_47278_10496# a_48282_10496# 0.97fF
C6233 cgen.dlycontrol3_in[3] a_14379_6567# 0.76fF
C6234 VDD a_50290_12504# 0.54fF
C6235 VDD nmat.col[16] 4.30fF
C6236 VDD m2_28976_7214# 0.91fF
C6237 a_6283_31591# a_7717_14735# 0.69fF
C6238 VDD a_7407_17455# 0.39fF
C6239 a_22178_65166# vcm 0.62fF
C6240 a_29206_21540# vcm 0.65fF
C6241 VDD a_2603_22357# 0.48fF
C6242 pmat.row_n[13] pmat.rowoff_n[12] 0.70fF
C6243 VDD a_27198_60146# 0.52fF
C6244 a_11067_27239# a_28915_50959# 0.36fF
C6245 a_24591_28327# pmat.col[19] 0.36fF
C6246 a_18563_27791# a_21365_27247# 1.22fF
C6247 a_44266_58138# vcm 0.62fF
C6248 a_1923_61759# a_2163_65469# 0.73fF
C6249 VDD a_12076_62839# 0.30fF
C6250 a_19166_67174# m2_17932_66994# 0.96fF
C6251 a_18546_23546# ctopn 1.49fF
C6252 a_21174_17524# a_21174_16520# 1.00fF
C6253 m2_17932_59966# vcm 0.44fF
C6254 m2_31988_54946# m3_32120_55078# 2.79fF
C6255 _1192_.A2 _1184_.A2 4.54fF
C6256 a_2389_45859# a_2983_48071# 0.77fF
C6257 a_18546_19530# a_33130_19938# 0.35fF
C6258 a_23182_14512# ctopn 3.58fF
C6259 a_18162_60186# vcm 6.95fF
C6260 a_27198_12504# a_28202_12504# 0.97fF
C6261 a_18546_12502# a_37146_12910# 0.35fF
C6262 a_3351_27249# a_5899_21807# 0.43fF
C6263 _1187_.A2 pmat.col[7] 0.44fF
C6264 VDD a_13837_39069# 1.36fF
C6265 a_3339_59879# a_7658_71543# 0.73fF
C6266 a_40250_22544# a_41254_22544# 0.97fF
C6267 VDD a_22085_42902# 1.44fF
C6268 a_30663_50087# a_44774_40821# 0.45fF
C6269 VDD a_33222_16520# 0.52fF
C6270 _1154_.X vcm 1.47fF
C6271 VDD a_23090_55126# 0.42fF
C6272 a_24591_28327# nmat.col[21] 0.51fF
C6273 VDD a_43170_7890# 0.34fF
C6274 VDD a_1823_58237# 1.50fF
C6275 VDD a_20170_57134# 0.52fF
C6276 VDD a_12531_34743# 0.64fF
C6277 a_24591_28327# ANTENNA__1195__A1.DIODE 1.44fF
C6278 ANTENNA__1184__B1.DIODE a_16311_28327# 0.41fF
C6279 ANTENNA__1395__A2.DIODE a_13459_28111# 0.44fF
C6280 a_11067_27239# ANTENNA__1395__B1.DIODE 2.90fF
C6281 a_36234_69182# vcm 0.62fF
C6282 a_18546_23546# a_42166_23954# 0.35fF
C6283 VDD a_43191_49551# 0.41fF
C6284 cgen.dlycontrol3_in[2] a_31793_41570# 0.38fF
C6285 a_18546_9490# a_46182_9898# 0.35fF
C6286 a_41237_28585# inn_analog 0.37fF
C6287 a_45270_59142# vcm 0.62fF
C6288 a_28202_63158# pmat.col[9] 0.31fF
C6289 a_10873_38517# a_10953_34951# 0.37fF
C6290 _1154_.X _1194_.B1 1.30fF
C6291 VDD a_1687_13621# 0.58fF
C6292 a_1923_69823# a_2163_69821# 0.35fF
C6293 a_46274_62154# pmat.col[27] 0.31fF
C6294 a_40250_56130# ctopp 3.40fF
C6295 VDD a_49286_56130# 0.55fF
C6296 a_19166_71190# a_20170_71190# 0.97fF
C6297 a_41731_49525# a_40837_46261# 0.42fF
C6298 _1192_.A2 a_9411_2215# 0.34fF
C6299 cgen.enable_dlycontrol_in nmat.sw 1.90fF
C6300 a_22178_61150# vcm 0.62fF
C6301 ANTENNA__1187__B1.DIODE pmat.col[20] 0.38fF
C6302 a_32218_21540# ctopn 3.58fF
C6303 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm 140.26fF
C6304 a_1899_35051# a_2791_57703# 2.23fF
C6305 nmat.sample_n a_7717_14735# 2.64fF
C6306 VDD a_22733_47381# 0.40fF
C6307 VDD a_31214_22544# 0.52fF
C6308 a_43262_66170# ctopp 3.58fF
C6309 m2_46044_72014# m3_46176_72146# 2.79fF
C6310 a_18162_72234# ctopp 0.30fF
C6311 a_35244_32411# a_40951_31599# 0.33fF
C6312 a_49286_11500# a_50290_11500# 0.97fF
C6313 VDD a_28431_34735# 0.44fF
C6314 a_2791_57703# a_2419_53351# 0.64fF
C6315 VDD _1224_.X 23.50fF
C6316 a_36234_63158# ctopp 3.58fF
C6317 a_2407_49289# a_4075_68583# 0.40fF
C6318 VDD a_45270_63158# 0.52fF
C6319 a_7479_53909# a_7645_53909# 0.75fF
C6320 a_28202_17524# vcm 0.65fF
C6321 a_36234_56130# a_36234_55126# 1.00fF
C6322 a_4339_27804# a_9777_26935# 1.00fF
C6323 a_18546_61192# a_44174_61150# 0.35fF
C6324 nmat.col_n[21] nmat.col[26] 0.36fF
C6325 a_2727_58470# a_3508_69135# 0.39fF
C6326 a_29206_8488# vcm 0.64fF
C6327 VDD a_82787_13077# 0.31fF
C6328 a_30571_50959# a_38851_28327# 0.46fF
C6329 nmat.rowon_n[4] ctopn 1.40fF
C6330 VDD a_33283_42333# 1.16fF
C6331 VDD a_5547_14735# 0.52fF
C6332 a_6369_39465# a_2411_33749# 0.33fF
C6333 pmat.col[2] vcm 5.88fF
C6334 a_2199_13887# a_2439_13889# 0.69fF
C6335 pmat.col_n[28] m2_47048_54946# 0.47fF
C6336 a_45270_19532# vcm 0.65fF
C6337 VDD nmat.rowon_n[2] 6.55fF
C6338 _1179_.X ANTENNA__1195__A1.DIODE 2.08fF
C6339 ANTENNA__1196__A2.DIODE a_13459_28111# 0.36fF
C6340 a_43262_18528# a_43262_17524# 1.00fF
C6341 a_16800_47213# a_16083_50069# 0.88fF
C6342 pmat.rowoff_n[12] a_18546_68220# 4.09fF
C6343 a_14641_57167# pmat.rowoff_n[11] 0.86fF
C6344 a_1769_13103# a_1739_47893# 0.38fF
C6345 a_44266_10496# vcm 0.65fF
C6346 a_18546_13506# a_38150_13914# 0.35fF
C6347 a_10055_31591# _1194_.A2 0.40fF
C6348 a_10515_15055# a_13091_52047# 0.40fF
C6349 cgen.enable_dlycontrol_in a_11149_36924# 2.20fF
C6350 a_10873_39605# a_24833_40719# 0.62fF
C6351 a_3339_59879# a_11797_60431# 0.48fF
C6352 a_43262_63158# a_43262_62154# 1.00fF
C6353 VDD m2_51064_61974# 1.00fF
C6354 a_18546_60188# a_19074_60146# 0.35fF
C6355 pmat.col_n[1] ANTENNA__1395__A2.DIODE 1.04fF
C6356 a_41254_67174# ctopp 3.58fF
C6357 a_18546_18526# a_34134_18934# 0.35fF
C6358 a_5351_19913# a_3688_17179# 0.44fF
C6359 VDD a_50290_67174# 0.54fF
C6360 nmat.col_n[0] nmat.col[1] 6.69fF
C6361 _1192_.B1 a_15667_27239# 0.55fF
C6362 a_49286_22544# a_49286_21540# 1.00fF
C6363 a_24186_12504# vcm 0.65fF
C6364 a_29206_64162# ctopp 3.58fF
C6365 VDD a_39246_14512# 0.52fF
C6366 a_48282_14512# a_49286_14512# 0.97fF
C6367 VDD a_38242_64162# 0.52fF
C6368 nmat.col_n[31] nmat.col_n[24] 0.77fF
C6369 a_34226_55126# pmat.col[15] 0.38fF
C6370 a_47278_64162# a_48282_64162# 0.97fF
C6371 a_18823_50247# a_21279_48999# 0.71fF
C6372 a_42258_13508# a_42258_12504# 1.00fF
C6373 a_18162_20536# ctopn 1.49fF
C6374 VDD config_1_in[2] 1.26fF
C6375 VDD a_17996_44007# 1.31fF
C6376 a_12447_16143# a_14887_46377# 0.95fF
C6377 nmat.rowon_n[2] nmat.rowoff_n[2] 20.31fF
C6378 VDD m2_26968_24282# 0.62fF
C6379 a_22199_30287# nmat.col[12] 1.98fF
C6380 a_1591_31599# a_1923_53055# 1.32fF
C6381 pmat.row_n[8] a_18546_64204# 0.35fF
C6382 a_12069_38517# cgen.dlycontrol2_in[2] 1.24fF
C6383 VDD nmat.col_n[15] 5.32fF
C6384 VDD a_18777_51183# 0.53fF
C6385 a_12345_36924# a_16381_35286# 0.62fF
C6386 a_11317_36924# a_19086_34343# 0.45fF
C6387 a_24833_34191# a_28247_34191# 1.11fF
C6388 a_18546_69224# vcm 0.40fF
C6389 a_12987_26159# a_12449_22895# 0.32fF
C6390 a_31214_17524# ctopn 3.58fF
C6391 a_46274_11500# vcm 0.65fF
C6392 VDD a_22178_62154# 0.52fF
C6393 a_10147_29415# a_35520_30083# 0.70fF
C6394 cgen.enable_dlycontrol_in a_12116_40871# 0.61fF
C6395 a_32218_8488# ctopn 3.40fF
C6396 pmat.row_n[10] a_18546_66212# 0.35fF
C6397 a_26194_56130# a_27198_56130# 0.97fF
C6398 a_18546_56172# a_35138_56130# 0.35fF
C6399 VDD a_34134_24958# 0.39fF
C6400 m2_47048_24282# m2_48052_24282# 0.96fF
C6401 a_29937_31055# a_46027_44905# 0.57fF
C6402 a_37291_29397# nmat.col[29] 1.40fF
C6403 a_15667_27239# a_10441_21263# 0.30fF
C6404 a_48282_19532# ctopn 3.58fF
C6405 a_32218_65166# ctopp 3.58fF
C6406 VDD a_3983_41941# 0.44fF
C6407 a_11091_26311# a_8568_26703# 0.89fF
C6408 VDD a_41254_65166# 0.52fF
C6409 a_20475_49783# a_20619_49551# 0.38fF
C6410 VDD a_48282_21540# 0.52fF
C6411 a_49286_65166# a_49286_64162# 1.00fF
C6412 a_47278_10496# ctopn 3.58fF
C6413 VDD comp_latch 17.05fF
C6414 a_18546_68220# a_43170_68178# 0.35fF
C6415 a_50290_68178# vcm 0.62fF
C6416 ANTENNA__1187__B1.DIODE a_27763_27221# 2.53fF
C6417 VDD a_21174_70186# 0.52fF
C6418 ANTENNA__1190__A1.DIODE a_41731_49525# 0.30fF
C6419 VDD a_18546_17522# 32.63fF
C6420 VDD a_19675_51157# 0.31fF
C6421 VDD a_12225_74575# 0.46fF
C6422 a_38242_16520# a_38242_15516# 1.00fF
C6423 a_31214_62154# a_32218_62154# 0.97fF
C6424 _1196_.B1 ANTENNA__1395__B1.DIODE 0.68fF
C6425 nmat.col_n[7] vcm 2.82fF
C6426 a_44266_63158# pmat.col[25] 0.31fF
C6427 a_29206_66170# a_30210_66170# 0.97fF
C6428 a_18546_60188# a_48190_60146# 0.35fF
C6429 pmat.row_n[3] pmat.rowon_n[3] 20.76fF
C6430 nmat.sw a_2411_33749# 1.12fF
C6431 a_27198_12504# ctopn 3.58fF
C6432 VDD a_4123_32661# 0.36fF
C6433 VDD a_19166_8488# 0.60fF
C6434 a_12237_36596# a_22537_36911# 0.83fF
C6435 a_23182_56130# vcm 0.62fF
C6436 VDD a_25209_36965# 1.33fF
C6437 ANTENNA__1196__A2.DIODE a_9528_20407# 0.48fF
C6438 VDD a_9183_72007# 0.36fF
C6439 a_2727_58470# pmat.rowoff_n[7] 0.50fF
C6440 nmat.col[9] nmat.col_n[9] 1.05fF
C6441 a_22178_63158# a_23182_63158# 0.97fF
C6442 a_18546_63200# a_27106_63158# 0.35fF
C6443 VDD m2_46044_72014# 1.00fF
C6444 a_46274_69182# ctopp 3.58fF
C6445 a_26194_66170# vcm 0.62fF
C6446 m2_36004_72014# m2_37008_72014# 0.96fF
C6447 a_10515_15055# a_9135_60967# 0.46fF
C6448 a_33423_47695# a_7415_29397# 0.31fF
C6449 VDD cgen.dlycontrol4_in[2] 8.55fF
C6450 ANTENNA__1197__B.DIODE ANTENNA__1183__B1.DIODE 4.03fF
C6451 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 1.46fF
C6452 pmat.col[5] m2_23956_54946# 0.39fF
C6453 a_49286_11500# ctopn 3.57fF
C6454 VDD a_15660_31029# 0.36fF
C6455 a_2695_76757# a_2999_76922# 0.62fF
C6456 VDD a_3413_6037# 0.34fF
C6457 pmat.col_n[6] _1187_.A2 0.33fF
C6458 a_13275_48783# a_40949_48437# 0.38fF
C6459 nmat.col_n[31] ctopn 2.16fF
C6460 pmat.rowon_n[8] a_6283_31591# 1.06fF
C6461 m2_51064_23278# vcm 0.51fF
C6462 VDD a_19505_38779# 1.08fF
C6463 a_32218_61150# ctopp 3.58fF
C6464 a_30210_70186# a_31214_70186# 0.97fF
C6465 VDD a_18162_9492# 2.74fF
C6466 VDD a_41254_61150# 0.52fF
C6467 VDD a_33309_41479# 1.09fF
C6468 a_24374_29941# ANTENNA__1183__B1.DIODE 0.61fF
C6469 VDD a_35230_20536# 0.52fF
C6470 a_15667_27239# a_43720_32143# 1.13fF
C6471 nmat.col[4] ctopn 1.97fF
C6472 a_22178_10496# a_22178_9492# 1.00fF
C6473 a_24186_67174# vcm 0.62fF
C6474 a_18546_71232# a_32126_71190# 0.35fF
C6475 a_33222_23548# m2_32992_24282# 0.99fF
C6476 a_12069_38517# a_11339_39319# 0.36fF
C6477 a_18546_72236# a_49194_72194# 0.35fF
C6478 a_13432_62581# a_5462_62215# 0.41fF
C6479 VDD a_47278_17524# 0.52fF
C6480 VDD m2_22952_54946# 0.62fF
C6481 VDD a_38569_46831# 0.57fF
C6482 a_18546_8486# a_40158_8894# 0.35fF
C6483 a_23182_60146# a_23182_59142# 1.00fF
C6484 pmat.row_n[3] pmat.rowoff_n[2] 1.15fF
C6485 a_18546_65208# a_37146_65166# 0.35fF
C6486 pmat.row_n[4] nmat.sample 0.34fF
C6487 a_1591_67503# a_2163_67645# 0.63fF
C6488 VDD a_31263_32117# 0.42fF
C6489 VDD a_48282_8488# 0.55fF
C6490 nmat.col_n[0] vcm 2.80fF
C6491 pmat.col_n[9] ctopp 2.02fF
C6492 a_12069_36341# a_12309_36483# 0.73fF
C6493 a_18546_21538# a_51202_21946# 0.35fF
C6494 VDD a_4601_35727# 0.41fF
C6495 m2_51064_64986# m2_51064_63982# 0.99fF
C6496 a_2411_33749# a_1858_25615# 0.50fF
C6497 VDD a_35138_72194# 0.33fF
C6498 a_41254_62154# a_41254_61150# 1.00fF
C6499 VDD a_5579_12394# 1.81fF
C6500 a_10441_21263# a_14943_26703# 0.40fF
C6501 a_50290_67174# m2_51064_66994# 0.96fF
C6502 VDD a_9557_17705# 0.42fF
C6503 a_4068_25615# a_7140_27805# 0.58fF
C6504 a_27198_67174# a_28202_67174# 0.97fF
C6505 a_18546_67216# a_37146_67174# 0.35fF
C6506 pmat.row_n[0] a_18162_56170# 25.57fF
C6507 a_11067_16359# a_5682_56311# 0.74fF
C6508 nmat.rowon_n[12] a_12079_9615# 0.85fF
C6509 a_24186_66170# a_24186_65166# 1.00fF
C6510 VDD a_24186_15516# 0.52fF
C6511 ANTENNA__1190__A2.DIODE nmat.col_n[19] 7.95fF
C6512 a_11041_40948# a_12197_41570# 1.69fF
C6513 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[31] 0.35fF
C6514 a_41254_15516# a_41254_14512# 1.00fF
C6515 pmat.en_bit_n[2] a_7717_14735# 1.21fF
C6516 pmat.col_n[22] pmat.col[22] 0.74fF
C6517 a_18546_7482# a_37146_7890# 0.35fF
C6518 ANTENNA__1197__A.DIODE ANTENNA__1187__B1.DIODE 0.97fF
C6519 pmat.row_n[0] nmat.rowon_n[15] 20.50fF
C6520 a_43262_69182# a_43262_68178# 1.00fF
C6521 a_21174_68178# a_22178_68178# 0.97fF
C6522 VDD a_31399_30511# 0.50fF
C6523 _1154_.X nmat.col_n[7] 1.08fF
C6524 pmat.rowon_n[8] nmat.col[7] 1.02fF
C6525 VDD pmat.row_n[14] 15.58fF
C6526 VDD a_43262_12504# 0.52fF
C6527 VDD nmat.col[28] 7.29fF
C6528 ANTENNA__1187__B1.DIODE clk_comp 1.55fF
C6529 VDD a_1823_76181# 1.43fF
C6530 a_22178_21540# vcm 0.65fF
C6531 pmat.col_n[11] ANTENNA__1187__B1.DIODE 0.33fF
C6532 pmat.col_n[10] a_11067_27239# 0.37fF
C6533 VDD a_14839_66103# 0.98fF
C6534 VDD a_2511_25615# 0.47fF
C6535 VDD a_20170_60146# 0.52fF
C6536 a_50290_71190# vcm 0.60fF
C6537 pmat.row_n[5] a_18546_61192# 0.35fF
C6538 a_7415_29397# a_6830_22895# 0.47fF
C6539 a_37238_58138# vcm 0.62fF
C6540 nmat.rowoff_n[11] a_18546_12502# 4.09fF
C6541 cgen.dlycontrol4_in[4] a_1895_26372# 0.34fF
C6542 a_25575_31055# a_6664_26159# 0.82fF
C6543 m2_51064_19262# m2_51064_18258# 0.99fF
C6544 a_18546_19530# a_26102_19938# 0.35fF
C6545 VDD a_20475_49783# 5.10fF
C6546 a_18546_12502# a_30118_12910# 0.35fF
C6547 a_1586_18231# a_1757_23445# 0.33fF
C6548 VDD a_26194_16520# 0.52fF
C6549 VDD m2_50060_24282# 0.50fF
C6550 a_18241_31698# a_23933_32143# 0.69fF
C6551 a_1769_47919# a_1957_43567# 1.29fF
C6552 VDD a_29635_31029# 0.58fF
C6553 VDD a_36142_7890# 0.33fF
C6554 a_45270_11500# a_45270_10496# 1.00fF
C6555 VDD a_47591_35407# 0.43fF
C6556 nmat.en_C0_n nmat.col_n[1] 0.30fF
C6557 a_29206_69182# vcm 0.62fF
C6558 VDD a_11693_70767# 0.49fF
C6559 _1154_.A a_13275_48783# 0.43fF
C6560 a_11067_64015# pmat.rowon_n[0] 0.63fF
C6561 a_2419_69455# nmat.rowon_n[7] 0.47fF
C6562 a_18546_23546# a_35138_23954# 0.35fF
C6563 a_26194_23548# a_27198_23548# 0.97fF
C6564 a_15667_27239# a_30663_50087# 0.82fF
C6565 m2_31988_24282# vcm 0.42fF
C6566 m2_17932_20266# m3_18064_20398# 2.76fF
C6567 VDD m2_17932_64986# 1.00fF
C6568 VDD a_25802_48169# 1.75fF
C6569 a_2411_43301# a_6559_33767# 0.72fF
C6570 a_18546_9490# a_39154_9898# 0.35fF
C6571 a_28202_9492# a_29206_9492# 0.97fF
C6572 pmat.row_n[2] a_18546_10494# 0.35fF
C6573 ANTENNA__1190__A1.DIODE vcm 1.66fF
C6574 a_38242_59142# vcm 0.62fF
C6575 a_35230_12504# a_35230_11500# 1.00fF
C6576 _1192_.B1 a_44870_48437# 0.59fF
C6577 VDD a_25319_42359# 0.60fF
C6578 a_11067_27239# _1192_.B1 1.04fF
C6579 a_17842_27497# a_18200_27497# 0.43fF
C6580 pmat.row_n[1] pmat.rowoff_n[2] 1.83fF
C6581 a_18546_17522# a_20078_17930# 0.35fF
C6582 a_18162_17524# nmat.rowon_n[6] 1.33fF
C6583 a_12197_41570# a_14589_40726# 3.01fF
C6584 a_33222_56130# ctopp 3.40fF
C6585 pmat.rowoff_n[12] a_14641_57711# 0.95fF
C6586 VDD a_33011_29941# 0.41fF
C6587 a_2648_29397# a_5173_9839# 0.55fF
C6588 VDD a_42258_56130# 0.55fF
C6589 a_44266_20536# a_45270_20536# 0.97fF
C6590 a_10239_14183# nmat.col[10] 0.31fF
C6591 a_12809_69679# a_13203_70767# 0.37fF
C6592 VDD a_2944_52789# 0.38fF
C6593 a_18546_15514# ctopn 1.59fF
C6594 _1192_.B1 a_35312_31599# 0.36fF
C6595 VDD a_18546_11498# 32.64fF
C6596 a_13459_28111# a_2007_25597# 1.54fF
C6597 a_2215_47375# a_2411_43301# 0.85fF
C6598 a_1923_61759# a_2215_47375# 0.50fF
C6599 VDD m3_18064_69134# 0.32fF
C6600 pmat.rowon_n[0] a_3576_17143# 1.58fF
C6601 a_25190_21540# ctopn 3.58fF
C6602 a_24591_28327# a_39939_29967# 0.62fF
C6603 a_18546_15514# a_20078_15922# 0.35fF
C6604 _1187_.A2 nmat.en_bit_n[1] 1.18fF
C6605 a_23395_53135# a_11067_27239# 0.35fF
C6606 a_43262_9492# a_43262_8488# 1.00fF
C6607 a_18546_65208# a_18162_65206# 2.62fF
C6608 VDD a_24186_22544# 0.52fF
C6609 a_36234_66170# ctopp 3.58fF
C6610 VDD a_45270_66170# 0.52fF
C6611 _1196_.B1 a_44533_33749# 1.28fF
C6612 a_25190_21540# a_26194_21540# 0.97fF
C6613 VDD pmat.col_n[2] 5.30fF
C6614 a_29206_63158# ctopp 3.58fF
C6615 VDD a_38242_63158# 0.52fF
C6616 a_21174_17524# vcm 0.65fF
C6617 a_30431_37683# ndecision_finish 0.94fF
C6618 m2_27972_24282# m3_28104_24414# 2.79fF
C6619 a_18546_67216# a_18162_67214# 2.62fF
C6620 nmat.col[24] m2_43032_24282# 0.39fF
C6621 a_18546_61192# a_37146_61150# 0.35fF
C6622 VDD a_14371_25071# 0.81fF
C6623 a_6664_26159# a_2683_22089# 0.40fF
C6624 a_20170_62154# pmat.col[1] 0.31fF
C6625 m2_43032_54946# m2_44036_54946# 0.96fF
C6626 a_26194_71190# a_26194_70186# 1.00fF
C6627 a_22178_8488# vcm 0.64fF
C6628 a_6467_29415# a_6821_18543# 0.40fF
C6629 a_40250_58138# a_41254_58138# 0.97fF
C6630 a_1781_9308# a_18241_31698# 1.84fF
C6631 VDD a_12228_40693# 3.43fF
C6632 a_11067_27239# a_10441_21263# 1.00fF
C6633 VDD a_3609_65015# 0.66fF
C6634 pmat.col_n[24] m2_43032_54946# 0.37fF
C6635 nmat.sample_n a_7415_29397# 1.63fF
C6636 VDD a_22307_27791# 1.25fF
C6637 a_38242_19532# vcm 0.65fF
C6638 VDD a_10339_21263# 0.40fF
C6639 nmat.rowon_n[7] a_10515_15055# 1.48fF
C6640 a_13091_28327# a_16311_28327# 2.45fF
C6641 m2_51064_72014# vcm 0.34fF
C6642 VDD a_31263_28309# 1.54fF
C6643 pmat.sample_n a_14839_66103# 0.81fF
C6644 a_38557_48469# a_33423_47695# 0.62fF
C6645 a_37238_10496# vcm 0.65fF
C6646 a_24186_13508# a_25190_13508# 0.97fF
C6647 a_18546_13506# a_31122_13914# 0.35fF
C6648 VDD a_3175_72641# 0.50fF
C6649 a_2727_58470# a_1591_61519# 0.91fF
C6650 a_2263_43719# a_31675_47695# 0.35fF
C6651 a_20170_16520# a_20170_15516# 1.00fF
C6652 pmat.rowoff_n[4] pmat.row_n[5] 0.36fF
C6653 a_36234_71190# m2_36004_72014# 1.00fF
C6654 VDD cgen.dlycontrol3_in[2] 6.36fF
C6655 a_40250_61150# a_40250_60146# 1.00fF
C6656 a_34226_67174# ctopp 3.58fF
C6657 a_48282_19532# a_48282_18528# 1.00fF
C6658 a_22178_18528# a_23182_18528# 0.97fF
C6659 a_18546_18526# a_27106_18934# 0.35fF
C6660 ANTENNA__1395__B1.DIODE a_45019_38645# 0.59fF
C6661 VDD a_43262_67174# 0.52fF
C6662 a_16083_50069# a_18547_51565# 1.91fF
C6663 a_22178_64162# ctopp 3.58fF
C6664 VDD a_32218_14512# 0.52fF
C6665 m2_51064_11230# vcm 0.51fF
C6666 m2_20944_7214# m3_21076_7346# 2.79fF
C6667 VDD a_31214_64162# 0.52fF
C6668 nmat.en_bit_n[0] a_12851_28853# 0.50fF
C6669 VDD a_17996_40743# 1.25fF
C6670 a_18546_17522# a_49194_17930# 0.35fF
C6671 VDD a_19965_39867# 1.28fF
C6672 a_18546_57176# a_45178_57134# 0.35fF
C6673 ANTENNA__1196__A2.DIODE a_12079_9615# 0.39fF
C6674 a_41254_59142# a_41254_58138# 1.00fF
C6675 a_19541_28879# a_11784_47099# 0.60fF
C6676 a_12585_39355# a_14600_37607# 0.51fF
C6677 ANTENNA__1197__B.DIODE a_21739_29415# 1.59fF
C6678 VDD m3_18064_16382# 0.33fF
C6679 a_24833_40719# a_12116_40871# 0.52fF
C6680 cgen.dlycontrol4_in[2] a_11113_40835# 0.96fF
C6681 pmat.en_bit_n[0] ANTENNA__1395__A2.DIODE 0.80fF
C6682 a_18546_15514# a_49194_15922# 0.35fF
C6683 a_33222_15516# a_34226_15516# 0.97fF
C6684 a_38851_28327# a_44444_32233# 0.31fF
C6685 pmat.rowon_n[2] pmat.row_n[2] 20.04fF
C6686 VDD m2_46044_54946# 0.62fF
C6687 a_32218_69182# a_33222_69182# 0.97fF
C6688 VDD a_38905_28853# 1.85fF
C6689 VDD a_5935_6575# 0.40fF
C6690 VDD a_47592_35643# 0.32fF
C6691 a_24186_17524# ctopn 3.58fF
C6692 VDD dummypin[9] 1.11fF
C6693 a_39246_11500# vcm 0.65fF
C6694 _1154_.X ANTENNA__1190__A1.DIODE 3.06fF
C6695 a_2419_53351# a_3345_62839# 0.96fF
C6696 a_18162_22544# ctopn 1.47fF
C6697 a_11317_36924# clk_dig 1.84fF
C6698 a_46274_17524# a_46274_16520# 1.00fF
C6699 m2_27972_54946# vcm 0.42fF
C6700 a_25190_8488# ctopn 3.40fF
C6701 a_18546_56172# a_28110_56130# 0.35fF
C6702 a_18546_9490# a_21082_9898# 0.35fF
C6703 VDD a_27106_24958# 0.44fF
C6704 m2_40020_24282# m2_41024_24282# 0.96fF
C6705 pmat.col[6] vcm 5.88fF
C6706 pmat.row_n[7] pmat.rowon_n[3] 4.46fF
C6707 a_41254_19532# ctopn 3.58fF
C6708 a_25190_65166# ctopp 3.58fF
C6709 VDD a_37739_43177# 0.64fF
C6710 nmat.en_bit_n[1] pmat.col[1] 0.66fF
C6711 m2_51064_8218# m2_51064_7214# 0.99fF
C6712 VDD a_34226_65166# 0.52fF
C6713 cgen.dlycontrol3_in[4] cgen.dlycontrol4_in[1] 0.37fF
C6714 _1184_.A2 a_9777_26935# 1.04fF
C6715 VDD nmat.col[0] 12.13fF
C6716 VDD a_41254_21540# 0.52fF
C6717 a_41254_59142# a_42258_59142# 0.97fF
C6718 a_16311_28327# a_17139_30503# 1.30fF
C6719 pmat.col_n[16] pmat.en_bit_n[2] 0.34fF
C6720 a_40250_10496# ctopn 3.58fF
C6721 a_18546_68220# a_36142_68178# 0.35fF
C6722 VDD ANTENNA__1183__B1.DIODE 22.36fF
C6723 a_47278_58138# ctopp 3.58fF
C6724 a_43262_68178# vcm 0.62fF
C6725 VDD a_3583_11775# 0.48fF
C6726 VDD nmat.col[25] 4.32fF
C6727 a_30210_23548# a_30210_22544# 1.00fF
C6728 VDD a_11807_51157# 0.56fF
C6729 VDD a_1823_74557# 1.84fF
C6730 nmat.col[10] ctopn 1.97fF
C6731 pmat.rowoff_n[7] config_1_in[15] 0.87fF
C6732 VDD a_30999_48071# 0.89fF
C6733 a_29206_60146# a_30210_60146# 0.97fF
C6734 a_18546_60188# a_41162_60146# 0.35fF
C6735 a_18546_66212# ctopp 1.59fF
C6736 pmat.row_n[7] a_2648_29397# 0.42fF
C6737 pmat.row_n[5] nmat.rowon_n[10] 20.11fF
C6738 a_38851_28327# a_32687_46607# 2.97fF
C6739 pmat.sample pmat.rowon_n[7] 0.41fF
C6740 m2_38012_54946# m3_38144_55078# 2.79fF
C6741 VDD m2_31988_72014# 1.12fF
C6742 a_37238_68178# a_37238_67174# 1.00fF
C6743 _1196_.B1 _1192_.B1 0.72fF
C6744 a_48282_23548# vcm 0.65fF
C6745 a_18546_61192# a_18162_61190# 2.62fF
C6746 a_39246_69182# ctopp 3.58fF
C6747 a_31675_47695# a_40105_47375# 1.63fF
C6748 a_50290_9492# vcm 0.65fF
C6749 VDD a_48282_69182# 0.52fF
C6750 pmat.en_bit_n[2] ANTENNA__1195__A1.DIODE 0.54fF
C6751 m2_28976_72014# m2_29980_72014# 0.96fF
C6752 VDD a_20811_39095# 0.60fF
C6753 a_6292_65479# a_5081_53135# 0.31fF
C6754 a_6927_30503# nmat.sw 0.52fF
C6755 a_30278_30511# a_29163_29423# 0.49fF
C6756 VDD a_2559_46261# 0.43fF
C6757 a_20170_19532# vcm 0.65fF
C6758 a_9963_13967# nmat.rowoff_n[1] 0.44fF
C6759 a_48282_59142# ctopp 3.58fF
C6760 a_42258_11500# ctopn 3.58fF
C6761 _1196_.B1 a_23395_53135# 0.92fF
C6762 VDD a_24565_34789# 1.33fF
C6763 a_8491_47911# a_5682_56311# 0.59fF
C6764 VDD a_10471_12791# 0.57fF
C6765 a_5579_12394# a_4895_12559# 0.48fF
C6766 nmat.col_n[7] nmat.col_n[0] 0.53fF
C6767 ANTENNA__1196__A2.DIODE a_32405_32463# 1.64fF
C6768 a_35230_16520# a_36234_16520# 0.97fF
C6769 a_2835_13077# a_12815_8213# 0.34fF
C6770 a_9135_62613# a_9301_62613# 0.69fF
C6771 a_6835_51183# a_5682_56311# 0.82fF
C6772 a_25190_67174# a_25190_66170# 1.00fF
C6773 VDD a_2411_16101# 4.49fF
C6774 VDD a_2743_38279# 0.40fF
C6775 a_25190_61150# ctopp 3.58fF
C6776 pmat.sw clk_ena 0.45fF
C6777 VDD a_6872_8725# 0.50fF
C6778 VDD a_34226_61150# 0.52fF
C6779 VDD a_22725_40229# 1.56fF
C6780 inp_analog m2_50060_54946# 0.73fF
C6781 a_46274_13508# vcm 0.65fF
C6782 VDD a_1717_13647# 5.58fF
C6783 a_12447_16143# a_12263_50959# 0.70fF
C6784 a_5320_27023# a_6323_26409# 0.32fF
C6785 a_1586_50247# a_2935_38279# 0.60fF
C6786 VDD a_7797_63151# 1.36fF
C6787 a_18546_55168# a_35138_55126# 0.39fF
C6788 VDD config_2_in[0] 0.76fF
C6789 a_28704_29568# a_6664_26159# 0.32fF
C6790 a_44266_18528# vcm 0.65fF
C6791 a_21371_50087# a_21279_48999# 0.43fF
C6792 a_25695_28111# nmat.col[15] 1.53fF
C6793 VDD a_28202_20536# 0.52fF
C6794 _1154_.A a_25695_28111# 0.86fF
C6795 a_24186_17524# a_25190_17524# 0.97fF
C6796 a_18243_28327# a_27763_27221# 3.11fF
C6797 a_7521_47081# a_7373_49007# 0.42fF
C6798 pmat.row_n[5] nmat.rowoff_n[14] 0.50fF
C6799 a_22178_57134# a_23182_57134# 0.97fF
C6800 pmat.col[25] m2_44036_54946# 0.39fF
C6801 VDD a_2787_55535# 0.42fF
C6802 a_27198_20536# a_27198_19532# 1.00fF
C6803 a_8305_20871# clk_dig 0.39fF
C6804 a_21174_71190# a_22178_71190# 0.97fF
C6805 a_18546_71232# a_25098_71190# 0.35fF
C6806 VDD a_4995_52815# 0.62fF
C6807 a_2419_69455# a_3345_62839# 2.16fF
C6808 pmat.col_n[24] pmat.col[25] 6.04fF
C6809 VDD a_40250_17524# 0.52fF
C6810 VDD a_37795_29111# 0.35fF
C6811 a_25190_8488# a_26194_8488# 0.97fF
C6812 a_18546_8486# a_33130_8894# 0.35fF
C6813 pmat.rowon_n[8] a_5363_33551# 0.84fF
C6814 a_18546_65208# a_30118_65166# 0.35fF
C6815 a_2835_13077# a_8656_12675# 0.60fF
C6816 m2_51064_72014# m3_51196_72146# 2.79fF
C6817 a_44266_70186# a_44266_69182# 1.00fF
C6818 VDD a_41254_8488# 0.55fF
C6819 a_21365_27247# nmat.col_n[7] 1.98fF
C6820 a_18546_21538# a_44174_21946# 0.35fF
C6821 a_2419_53351# a_3615_71631# 0.58fF
C6822 nmat.col[31] a_28812_29575# 0.53fF
C6823 a_33222_14512# a_33222_13508# 1.00fF
C6824 a_2407_49289# a_5651_66975# 0.34fF
C6825 a_11339_39319# a_17536_38567# 0.60fF
C6826 a_18546_67216# a_30118_67174# 0.35fF
C6827 a_37238_57134# a_37238_56130# 1.00fF
C6828 VDD result_out[1] 0.75fF
C6829 a_41254_19532# a_42258_19532# 0.97fF
C6830 nmat.rowon_n[7] ANTENNA__1184__B1.DIODE 1.18fF
C6831 ANTENNA__1195__A1.DIODE a_28336_29967# 0.81fF
C6832 pmat.col_n[4] vcm 2.80fF
C6833 a_9963_28111# nmat.col_n[12] 0.32fF
C6834 a_4351_55527# a_4075_50087# 1.26fF
C6835 a_18546_7482# a_30118_7890# 0.35fF
C6836 a_30663_50087# a_35312_31599# 2.06fF
C6837 nmat.rowon_n[7] a_10515_61839# 1.93fF
C6838 VDD a_10851_30485# 0.52fF
C6839 a_40250_10496# a_41254_10496# 0.97fF
C6840 VDD result_out[10] 0.62fF
C6841 VDD a_36234_12504# 0.52fF
C6842 VDD pmat.col[30] 4.31fF
C6843 a_18546_58180# ctopp 1.59fF
C6844 nmat.sw a_10873_40693# 3.17fF
C6845 a_49286_13508# ctopn 3.57fF
C6846 a_44266_57134# vcm 0.62fF
C6847 a_43262_71190# vcm 0.60fF
C6848 a_47278_18528# ctopn 3.58fF
C6849 a_21739_29415# a_22459_28879# 2.07fF
C6850 a_30210_58138# vcm 0.62fF
C6851 a_37238_56130# m2_37008_54946# 0.99fF
C6852 a_28915_50959# a_22199_30287# 0.53fF
C6853 pmat.en_bit_n[0] a_29455_31293# 0.50fF
C6854 nmat.col_n[26] nmat.col_n[29] 10.31fF
C6855 VDD a_13795_10687# 0.36fF
C6856 VDD a_15747_50069# 0.41fF
C6857 a_18546_12502# a_23090_12910# 0.35fF
C6858 VDD m3_43164_7346# 0.38fF
C6859 a_33222_22544# a_34226_22544# 0.97fF
C6860 VDD a_28245_44581# 1.17fF
C6861 VDD a_18162_16520# 2.74fF
C6862 m2_51064_69002# m3_51196_69134# 2.76fF
C6863 VDD a_38913_31055# 1.12fF
C6864 pmat.rowoff_n[15] a_18162_23548# 1.33fF
C6865 VDD a_29114_7890# 0.33fF
C6866 nmat.col_n[17] a_36234_24552# 0.32fF
C6867 a_16311_28327# a_9411_2215# 3.26fF
C6868 a_20475_49783# a_22499_49783# 2.50fF
C6869 a_12175_27221# nmat.col_n[1] 0.33fF
C6870 a_22178_69182# vcm 0.62fF
C6871 VDD pmat.rowon_n[15] 3.84fF
C6872 a_46705_38671# a_46947_39215# 0.30fF
C6873 a_18546_23546# a_28110_23954# 0.35fF
C6874 a_28336_29967# a_32865_30199# 0.37fF
C6875 cgen.dlycontrol4_in[4] cgen.dlycontrol4_in[2] 0.42fF
C6876 a_47278_63158# a_48282_63158# 0.97fF
C6877 cgen.dlycontrol3_in[2] a_11113_40835# 8.19fF
C6878 a_18546_9490# a_32126_9898# 0.35fF
C6879 nmat.col_n[12] a_9583_10121# 0.43fF
C6880 a_1957_43567# a_11455_50237# 0.34fF
C6881 a_31214_59142# vcm 0.62fF
C6882 VDD a_2263_43719# 11.21fF
C6883 a_32687_46607# a_37827_30793# 0.36fF
C6884 ANTENNA__1190__A1.DIODE a_40837_46261# 0.61fF
C6885 a_13091_52047# a_13091_28327# 0.45fF
C6886 ANTENNA__1197__A.DIODE a_18243_28327# 1.61fF
C6887 pmat.row_n[5] vcm 1.19fF
C6888 m2_17932_14242# vcm 0.44fF
C6889 a_26194_56130# ctopp 3.40fF
C6890 VDD a_12461_29673# 2.00fF
C6891 pmat.rowoff_n[15] nmat.sw 1.11fF
C6892 a_10953_34951# a_11409_34789# 0.46fF
C6893 VDD a_35230_56130# 0.54fF
C6894 a_1674_68047# a_2695_76757# 0.30fF
C6895 a_26194_8488# m2_25964_7214# 1.00fF
C6896 VDD a_9675_10396# 2.52fF
C6897 m2_17932_18258# a_19166_18528# 0.96fF
C6898 VDD m3_28104_72146# 0.33fF
C6899 a_18546_62196# a_49194_62154# 0.35fF
C6900 a_6853_14967# a_6835_14735# 0.31fF
C6901 _1196_.B1 pmat.col[14] 0.56fF
C6902 a_18546_66212# a_45178_66170# 0.35fF
C6903 a_11067_16359# a_1957_43567# 3.63fF
C6904 a_29206_66170# ctopp 3.58fF
C6905 VDD a_38242_66170# 0.52fF
C6906 pmat.row_n[5] _1194_.B1 1.36fF
C6907 a_4955_40277# a_6127_40516# 0.36fF
C6908 a_42258_11500# a_43262_11500# 0.97fF
C6909 VDD a_40399_36911# 0.47fF
C6910 a_22178_63158# ctopp 3.58fF
C6911 VDD a_6559_53903# 0.50fF
C6912 VDD a_31214_63158# 0.52fF
C6913 pmat.row_n[6] a_18162_62194# 25.57fF
C6914 a_44266_64162# a_44266_63158# 1.00fF
C6915 a_4523_21276# a_14371_25071# 0.42fF
C6916 a_24407_31375# nmat.col_n[29] 0.56fF
C6917 ANTENNA__1197__A.DIODE a_28704_29568# 0.79fF
C6918 a_47278_10496# a_47278_9492# 1.00fF
C6919 a_18546_61192# a_30118_61150# 0.35fF
C6920 a_6664_26159# ANTENNA__1190__A2.DIODE 0.87fF
C6921 a_44266_58138# a_44266_57134# 1.00fF
C6922 a_9963_13967# a_14457_15823# 0.43fF
C6923 a_11041_40948# a_12585_40443# 0.34fF
C6924 a_10873_40693# a_12116_40871# 5.15fF
C6925 VDD a_2163_65469# 0.49fF
C6926 pmat.col_n[20] m2_39016_54946# 0.37fF
C6927 VDD nmat.col[31] 7.93fF
C6928 VDD a_21739_29415# 11.74fF
C6929 a_26891_28327# nmat.en_bit_n[2] 0.37fF
C6930 a_31214_19532# vcm 0.65fF
C6931 a_48282_60146# a_48282_59142# 1.00fF
C6932 a_36234_18528# a_36234_17524# 1.00fF
C6933 m2_51064_65990# m3_51196_66122# 2.76fF
C6934 VDD a_20310_28029# 0.86fF
C6935 pmat.rowoff_n[7] a_4976_16091# 1.45fF
C6936 a_30210_10496# vcm 0.65fF
C6937 a_18546_13506# a_24094_13914# 0.35fF
C6938 nmat.rowon_n[12] ctopn 1.40fF
C6939 a_36234_63158# a_36234_62154# 1.00fF
C6940 VDD a_21215_48071# 0.94fF
C6941 a_27198_67174# ctopp 3.58fF
C6942 VDD a_28079_38825# 0.61fF
C6943 a_18546_18526# a_19074_18934# 0.35fF
C6944 a_18546_70228# a_47186_70186# 0.35fF
C6945 a_7730_69109# a_7674_69135# 0.92fF
C6946 VDD a_36234_67174# 0.52fF
C6947 VDD a_33765_38053# 1.14fF
C6948 m2_17932_67998# m2_17932_66994# 0.99fF
C6949 a_49286_66170# a_49286_65166# 1.00fF
C6950 a_42258_22544# a_42258_21540# 1.00fF
C6951 a_8583_29199# a_22307_27791# 0.70fF
C6952 VDD a_40315_42089# 0.67fF
C6953 VDD a_25190_14512# 0.52fF
C6954 ANTENNA__1190__A1.DIODE a_21365_27247# 0.63fF
C6955 a_13091_52047# a_17139_30503# 0.50fF
C6956 a_41254_14512# a_42258_14512# 0.97fF
C6957 a_46274_62154# vcm 0.62fF
C6958 VDD a_24186_64162# 0.52fF
C6959 a_21371_50087# a_29076_48695# 0.67fF
C6960 VDD a_6127_40516# 0.37fF
C6961 a_18546_17522# a_42166_17930# 0.35fF
C6962 a_40250_64162# a_41254_64162# 0.97fF
C6963 a_13459_28111# inn_analog 0.37fF
C6964 a_46274_68178# a_47278_68178# 0.97fF
C6965 a_19166_68178# a_19166_67174# 1.00fF
C6966 a_18546_57176# a_38150_57134# 0.35fF
C6967 VDD a_4587_53505# 0.69fF
C6968 cgen.dlycontrol4_in[2] a_3325_36495# 0.57fF
C6969 a_3339_59879# a_12815_74581# 0.36fF
C6970 a_13091_28327# nmat.col_n[26] 0.79fF
C6971 a_2935_38279# cgen.dlycontrol3_in[1] 0.96fF
C6972 a_45270_8488# m2_45040_7214# 1.00fF
C6973 VDD a_4298_69367# 0.49fF
C6974 a_35230_13508# a_35230_12504# 1.00fF
C6975 a_12585_39355# a_13357_37429# 0.99fF
C6976 a_11067_30287# a_14917_23983# 0.45fF
C6977 a_18546_15514# a_42166_15922# 0.35fF
C6978 VDD a_40105_47375# 2.89fF
C6979 VDD a_51202_55126# 0.49fF
C6980 nmat.sw a_12934_35823# 0.30fF
C6981 cgen.enable_dlycontrol_in clk_dig 0.94fF
C6982 pmat.col_n[12] ctopp 2.02fF
C6983 pmat.rowon_n[3] a_6553_53047# 0.85fF
C6984 a_9963_13967# a_4259_31375# 2.09fF
C6985 VDD a_19689_35877# 1.19fF
C6986 a_45270_70186# vcm 0.62fF
C6987 a_33957_48437# a_33467_46261# 0.81fF
C6988 VDD a_38150_72194# 0.32fF
C6989 a_32218_11500# vcm 0.65fF
C6990 VDD a_18546_13506# 32.63fF
C6991 ANTENNA__1187__B1.DIODE a_33467_46261# 0.65fF
C6992 a_11067_16359# cgen.enable_dlycontrol_in 1.06fF
C6993 VDD m2_51064_16250# 1.15fF
C6994 a_7693_22365# a_5899_21807# 0.53fF
C6995 ANTENNA__1187__B1.DIODE ANTENNA__1184__B1.DIODE 10.32fF
C6996 a_24867_53135# ANTENNA__1197__B.DIODE 0.91fF
C6997 a_18546_56172# a_21082_56130# 0.35fF
C6998 a_7026_24527# a_9528_20407# 0.35fF
C6999 pmat.row_n[4] pmat.row_n[3] 0.70fF
C7000 a_18563_27791# nmat.col_n[13] 0.76fF
C7001 a_10873_38517# a_11297_36091# 1.12fF
C7002 VDD a_7067_53511# 0.40fF
C7003 a_1823_68565# a_2215_47375# 2.15fF
C7004 a_20438_35431# a_12069_36341# 0.56fF
C7005 a_34226_19532# ctopn 3.58fF
C7006 VDD a_17625_42902# 1.03fF
C7007 VDD a_27198_65166# 0.52fF
C7008 pmat.en_bit_n[0] a_2007_25597# 0.44fF
C7009 VDD a_9741_28585# 0.84fF
C7010 VDD a_34226_21540# 0.52fF
C7011 a_5363_33551# a_9307_31068# 1.32fF
C7012 a_42258_65166# a_42258_64162# 1.00fF
C7013 m2_51064_62978# m3_51196_63110# 2.76fF
C7014 a_33222_10496# ctopn 3.58fF
C7015 a_18546_68220# a_29114_68178# 0.35fF
C7016 ANTENNA__1190__A2.DIODE a_8197_20871# 0.33fF
C7017 _1184_.A2 a_10071_17999# 0.49fF
C7018 a_40250_58138# ctopp 3.58fF
C7019 a_36234_68178# vcm 0.62fF
C7020 pmat.rowon_n[8] a_5266_17143# 1.09fF
C7021 a_42258_63158# pmat.col[23] 0.31fF
C7022 VDD a_49286_58138# 0.52fF
C7023 a_4075_50087# a_3615_71631# 0.30fF
C7024 a_19166_15516# vcm 0.65fF
C7025 a_24186_62154# a_25190_62154# 0.97fF
C7026 a_31214_16520# a_31214_15516# 1.00fF
C7027 a_9319_15279# a_9485_15279# 0.66fF
C7028 a_18162_65206# vcm 6.95fF
C7029 VDD a_12328_48168# 0.38fF
C7030 nmat.col[12] vcm 5.78fF
C7031 _1154_.A _1224_.X 1.00fF
C7032 a_22178_66170# a_23182_66170# 0.97fF
C7033 cgen.dlycontrol4_in[0] a_1586_18231# 0.72fF
C7034 a_18546_60188# a_34134_60146# 0.35fF
C7035 a_4991_69831# a_11067_16359# 0.55fF
C7036 a_32405_32463# a_2007_25597# 1.35fF
C7037 a_16478_29423# a_15667_28111# 0.74fF
C7038 a_2411_43301# a_1591_43029# 0.34fF
C7039 pmat.row_n[13] vcm 1.26fF
C7040 a_6664_26159# a_15667_28111# 0.71fF
C7041 _1194_.A2 a_12175_27221# 0.42fF
C7042 pmat.row_n[11] clk_dig 0.32fF
C7043 a_12245_21807# a_12247_20175# 0.50fF
C7044 a_19166_17524# a_19166_16520# 1.00fF
C7045 VDD m2_17932_72014# 1.44fF
C7046 _1179_.X _1192_.A2 0.61fF
C7047 a_4075_68583# a_1769_47919# 0.50fF
C7048 a_41254_23548# vcm 0.65fF
C7049 a_32218_69182# ctopp 3.58fF
C7050 a_13091_28327# a_24407_31375# 1.62fF
C7051 a_43262_9492# vcm 0.65fF
C7052 VDD a_41254_69182# 0.52fF
C7053 m2_21948_72014# m2_22952_72014# 0.96fF
C7054 VDD a_2867_43541# 0.42fF
C7055 a_10515_13967# a_13091_18535# 4.12fF
C7056 a_3339_70759# a_4075_50087# 2.07fF
C7057 a_18241_31698# a_31263_32117# 1.40fF
C7058 a_43262_65166# a_44266_65166# 0.97fF
C7059 a_41254_59142# ctopp 3.58fF
C7060 VDD a_17047_27497# 0.42fF
C7061 a_35230_11500# ctopn 3.58fF
C7062 a_1586_18231# rst_n 1.14fF
C7063 VDD a_50290_59142# 0.56fF
C7064 a_11057_35836# a_11255_35862# 0.30fF
C7065 a_6283_31591# a_11067_30287# 4.00fF
C7066 a_33467_46261# a_33839_46805# 1.73fF
C7067 a_1739_47893# a_1769_14735# 0.57fF
C7068 a_9411_2215# a_10071_17999# 0.99fF
C7069 a_48282_63158# pmat.col[29] 0.31fF
C7070 a_18546_16518# a_46182_16926# 0.35fF
C7071 m2_41024_24282# vcm 0.42fF
C7072 a_7644_16341# a_3571_13627# 0.64fF
C7073 nmat.col_n[3] nmat.col_n[13] 0.40fF
C7074 a_23182_70186# a_24186_70186# 0.97fF
C7075 VDD a_27198_61150# 0.52fF
C7076 a_39246_13508# vcm 0.65fF
C7077 VDD a_33223_42359# 0.57fF
C7078 VDD a_10055_31591# 12.04fF
C7079 pmat.en_bit_n[0] a_31339_31787# 0.70fF
C7080 a_37238_18528# vcm 0.65fF
C7081 VDD a_21174_20536# 0.52fF
C7082 a_16311_28327# nmat.col[24] 0.86fF
C7083 m2_51064_59966# m3_51196_60098# 2.76fF
C7084 a_18546_57176# a_20078_57134# 0.35fF
C7085 pmat.row_n[11] vcm 1.16fF
C7086 a_18162_61190# vcm 6.95fF
C7087 a_49286_13508# a_50290_13508# 0.97fF
C7088 nmat.col[15] nmat.col_n[15] 0.64fF
C7089 a_1923_61759# a_9135_62613# 0.72fF
C7090 ANTENNA__1196__A2.DIODE a_40951_31599# 1.02fF
C7091 a_17139_30503# a_44757_37289# 0.59fF
C7092 a_48282_15516# vcm 0.65fF
C7093 VDD a_33222_17524# 0.52fF
C7094 a_18546_8486# a_26102_8894# 0.35fF
C7095 a_1769_47919# a_6927_30503# 1.15fF
C7096 a_18546_65208# a_23090_65166# 0.35fF
C7097 a_47278_18528# a_48282_18528# 0.97fF
C7098 VDD a_34226_8488# 0.55fF
C7099 VDD a_1591_31599# 4.50fF
C7100 a_8443_20719# nmat.col_n[3] 0.66fF
C7101 pmat.row_n[4] a_10839_11989# 0.32fF
C7102 a_18546_21538# a_37146_21946# 0.35fF
C7103 VDD a_22541_36603# 1.32fF
C7104 VDD pmat.col_n[5] 5.54fF
C7105 a_34226_62154# a_34226_61150# 1.00fF
C7106 a_44266_23548# ctopn 3.40fF
C7107 VDD a_50290_19532# 0.54fF
C7108 a_46274_9492# ctopn 3.57fF
C7109 m2_32992_24282# m3_33124_24414# 2.79fF
C7110 a_20170_67174# a_21174_67174# 0.97fF
C7111 a_18546_67216# a_23090_67174# 0.35fF
C7112 nmat.rowon_n[1] vcm 0.56fF
C7113 a_24407_31375# a_17139_30503# 0.37fF
C7114 nmat.col_n[21] nmat.col[22] 6.76fF
C7115 a_44266_60146# vcm 0.62fF
C7116 VDD a_49286_10496# 0.52fF
C7117 a_34226_15516# a_34226_14512# 1.00fF
C7118 VDD a_7027_29673# 0.39fF
C7119 a_18546_7482# a_23090_7890# 0.35fF
C7120 VDD a_3183_19258# 0.65fF
C7121 a_36234_69182# a_36234_68178# 1.00fF
C7122 VDD m2_17932_17254# 1.01fF
C7123 _1154_.X nmat.col[12] 0.37fF
C7124 a_44266_21540# a_44266_20536# 1.00fF
C7125 a_18546_68220# vcm 0.40fF
C7126 a_4259_31375# a_1923_31743# 0.66fF
C7127 VDD a_29206_12504# 0.52fF
C7128 a_50290_16520# vcm 0.65fF
C7129 a_10781_42869# a_10979_43222# 0.30fF
C7130 VDD a_13688_47893# 0.84fF
C7131 a_42258_13508# ctopn 3.58fF
C7132 VDD a_8569_60405# 0.63fF
C7133 _1192_.A2 pmat.col[0] 0.42fF
C7134 a_37238_57134# vcm 0.62fF
C7135 a_36234_71190# vcm 0.60fF
C7136 a_40250_18528# ctopn 3.58fF
C7137 VDD a_30857_41245# 1.34fF
C7138 a_23182_58138# vcm 0.62fF
C7139 pmat.row_n[0] a_13091_7655# 1.38fF
C7140 m2_25964_7214# m3_26096_7346# 2.79fF
C7141 VDD a_20605_40719# 1.17fF
C7142 m2_51064_56954# m3_51196_57086# 2.76fF
C7143 a_1674_57711# a_1591_56623# 0.40fF
C7144 a_8491_47911# a_1957_43567# 2.03fF
C7145 a_13327_70741# a_12809_69679# 0.31fF
C7146 a_23395_53135# pmat.col[12] 0.38fF
C7147 ANTENNA__1187__B1.DIODE a_13641_23439# 0.65fF
C7148 a_18546_69224# a_51202_69182# 0.35fF
C7149 VDD a_22086_7890# 0.33fF
C7150 a_38242_11500# a_38242_10496# 1.00fF
C7151 a_1586_18231# a_1591_20181# 0.81fF
C7152 VDD a_10591_35561# 0.60fF
C7153 a_44774_48695# a_21279_48999# 0.38fF
C7154 VDD a_18162_62194# 2.73fF
C7155 m2_37008_54946# vcm 0.42fF
C7156 a_21174_9492# a_22178_9492# 0.97fF
C7157 a_18546_9490# a_25098_9898# 0.35fF
C7158 a_48282_22544# vcm 0.65fF
C7159 a_43262_61150# a_44266_61150# 0.97fF
C7160 a_46274_68178# ctopp 3.58fF
C7161 a_11067_64015# a_6283_31591# 0.37fF
C7162 a_24186_59142# vcm 0.62fF
C7163 VDD a_5535_57993# 2.56fF
C7164 a_28202_12504# a_28202_11500# 1.00fF
C7165 VDD a_10949_42364# 2.32fF
C7166 a_1957_43567# a_11823_46973# 0.35fF
C7167 a_30663_50087# a_45019_38645# 1.23fF
C7168 a_24407_31375# a_26891_28327# 0.50fF
C7169 a_12520_51451# a_12559_51325# 0.79fF
C7170 VDD a_2237_29423# 0.39fF
C7171 VDD a_28202_56130# 0.55fF
C7172 a_37238_20536# a_38242_20536# 0.97fF
C7173 a_4075_31591# a_6007_33767# 0.38fF
C7174 _1519_.A vcm 5.56fF
C7175 VDD m2_44036_7214# 1.04fF
C7176 a_5687_71829# a_4025_54965# 0.32fF
C7177 a_18546_62196# a_42166_62154# 0.35fF
C7178 a_50290_67174# a_50290_66170# 1.00fF
C7179 a_18546_66212# a_38150_66170# 0.35fF
C7180 a_36234_9492# a_36234_8488# 1.00fF
C7181 pmat.row_n[9] pmat.rowon_n[9] 20.51fF
C7182 a_22178_66170# ctopp 3.58fF
C7183 m2_17932_72014# m3_18064_72146# 2.79fF
C7184 VDD a_31214_66170# 0.52fF
C7185 a_23395_53135# a_22199_30287# 0.31fF
C7186 nmat.col_n[30] nmat.col[18] 2.77fF
C7187 VDD a_24186_63158# 0.52fF
C7188 a_8583_29199# a_12461_29673# 0.39fF
C7189 a_29455_31293# a_10147_29415# 0.43fF
C7190 a_22628_30485# a_22186_30485# 0.65fF
C7191 a_49286_17524# a_50290_17524# 0.97fF
C7192 _1192_.B1 a_14947_26159# 0.41fF
C7193 m2_43032_54946# m3_43164_55078# 2.79fF
C7194 nmat.col[29] nmat.col_n[31] 0.77fF
C7195 a_13275_48783# a_40349_40726# 0.31fF
C7196 a_47278_57134# a_48282_57134# 0.97fF
C7197 a_18546_61192# a_23090_61150# 0.35fF
C7198 a_46274_71190# a_47278_71190# 0.97fF
C7199 a_12263_50959# a_19541_28879# 0.43fF
C7200 _1196_.B1 a_10883_3303# 0.95fF
C7201 VDD a_29827_39095# 0.63fF
C7202 a_33222_58138# a_34226_58138# 0.97fF
C7203 VDD a_30819_40191# 2.33fF
C7204 a_24186_19532# vcm 0.65fF
C7205 pmat.rowon_n[1] ctopp 1.56fF
C7206 ANTENNA__1187__B1.DIODE nmat.col_n[29] 1.95fF
C7207 cgen.dlycontrol3_in[4] nmat.sw 0.39fF
C7208 VDD a_11133_34427# 1.06fF
C7209 a_23182_10496# vcm 0.65fF
C7210 cgen.dlycontrol3_in[0] cgen.dlycontrol2_in[4] 4.00fF
C7211 a_2419_69455# a_3199_40455# 0.51fF
C7212 VDD a_36265_48981# 0.39fF
C7213 a_9135_60967# a_7939_31591# 1.30fF
C7214 a_33222_61150# a_33222_60146# 1.00fF
C7215 VDD a_10097_22895# 0.52fF
C7216 a_20170_67174# ctopp 3.57fF
C7217 VDD a_24867_53135# 9.32fF
C7218 a_41254_19532# a_41254_18528# 1.00fF
C7219 a_18546_70228# a_40158_70186# 0.35fF
C7220 pmat.row_n[13] a_18546_69224# 0.35fF
C7221 VDD a_29206_67174# 0.52fF
C7222 pmat.row_n[2] vcm 1.19fF
C7223 VDD a_29735_40183# 0.64fF
C7224 a_13357_37429# a_21219_36885# 0.77fF
C7225 a_19166_57134# vcm 0.61fF
C7226 VDD a_13443_38007# 0.61fF
C7227 pmat.sw a_13459_28111# 0.70fF
C7228 a_39246_62154# vcm 0.62fF
C7229 a_18546_17522# a_35138_17930# 0.35fF
C7230 pmat.row_n[1] a_18546_57176# 0.35fF
C7231 a_18546_57176# a_31122_57134# 0.35fF
C7232 a_14287_69455# pmat.rowoff_n[11] 1.48fF
C7233 VDD a_6559_33767# 6.72fF
C7234 a_34226_59142# a_34226_58138# 1.00fF
C7235 a_24407_31375# a_9411_2215# 0.31fF
C7236 a_8491_47911# a_4991_69831# 1.75fF
C7237 a_3746_58487# a_8079_46519# 0.38fF
C7238 cgen.start_conv_in a_14497_42658# 0.50fF
C7239 a_26194_15516# a_27198_15516# 0.97fF
C7240 a_18546_15514# a_35138_15922# 0.35fF
C7241 a_6835_51183# a_5211_57172# 0.84fF
C7242 VDD a_10772_77563# 0.57fF
C7243 a_25190_69182# a_26194_69182# 0.97fF
C7244 nmat.col_n[4] vcm 2.80fF
C7245 nmat.col[12] nmat.col_n[7] 4.29fF
C7246 nmat.col_n[17] ctopn 2.01fF
C7247 VDD a_11057_35836# 2.09fF
C7248 a_38242_70186# vcm 0.62fF
C7249 a_25190_11500# vcm 0.65fF
C7250 VDD a_2215_47375# 7.57fF
C7251 nmat.col_n[13] vcm 2.80fF
C7252 a_39246_17524# a_39246_16520# 1.00fF
C7253 m2_17932_55950# vcm 0.44fF
C7254 VDD a_12245_21807# 0.43fF
C7255 ANTENNA__1395__B1.DIODE nmat.col_n[3] 0.54fF
C7256 a_45270_12504# a_46274_12504# 0.97fF
C7257 _1187_.A2 nmat.col_n[31] 0.42fF
C7258 pmat.col_n[7] vcm 2.80fF
C7259 a_27198_19532# ctopn 3.58fF
C7260 VDD a_20170_65166# 0.52fF
C7261 a_15667_27239# nmat.col[21] 1.10fF
C7262 _1154_.X _1519_.A 11.06fF
C7263 a_2407_49289# a_5687_71829# 0.55fF
C7264 VDD a_27198_21540# 0.52fF
C7265 a_34226_59142# a_35230_59142# 0.97fF
C7266 a_18546_59184# a_51202_59142# 0.35fF
C7267 ANTENNA__1195__A1.DIODE a_15667_27239# 0.65fF
C7268 a_26194_10496# ctopn 3.58fF
C7269 a_18546_68220# a_22086_68178# 0.35fF
C7270 a_47278_57134# ctopp 3.57fF
C7271 a_2149_45717# a_6051_74183# 0.70fF
C7272 a_46274_71190# ctopp 3.40fF
C7273 a_33222_58138# ctopp 3.58fF
C7274 pmat.col[11] m2_29980_54946# 0.39fF
C7275 a_29206_68178# vcm 0.62fF
C7276 VDD a_3838_70455# 0.76fF
C7277 a_2215_47375# a_4719_30287# 0.48fF
C7278 _1196_.B1 cgen.dlycontrol1_in[3] 0.81fF
C7279 VDD a_42258_58138# 0.52fF
C7280 a_23182_23548# a_23182_22544# 1.00fF
C7281 VDD a_8385_51727# 0.91fF
C7282 _1194_.B1 nmat.rowoff_n[6] 0.36fF
C7283 VDD a_8197_76757# 0.67fF
C7284 a_38242_62154# pmat.col[19] 0.31fF
C7285 a_18546_66212# a_20078_66170# 0.35fF
C7286 a_18162_21540# vcm 6.95fF
C7287 a_18546_60188# a_27106_60146# 0.35fF
C7288 a_22178_60146# a_23182_60146# 0.97fF
C7289 ANTENNA__1197__A.DIODE _1194_.A2 0.90fF
C7290 VDD a_4508_65845# 0.81fF
C7291 a_2952_25045# a_4339_27804# 1.64fF
C7292 a_10515_15055# a_2046_30184# 1.11fF
C7293 a_2407_49289# a_4583_68021# 0.59fF
C7294 m2_17932_54946# m3_18064_55078# 2.79fF
C7295 a_30210_68178# a_30210_67174# 1.00fF
C7296 a_14641_57711# a_11067_16359# 0.60fF
C7297 a_34226_23548# vcm 0.65fF
C7298 a_25190_69182# ctopp 3.58fF
C7299 m2_18936_55950# m2_18936_54946# 0.99fF
C7300 a_36234_9492# vcm 0.65fF
C7301 VDD a_34226_69182# 0.52fF
C7302 VDD a_2972_9991# 1.72fF
C7303 VDD a_38851_28327# 13.26fF
C7304 cgen.dlycontrol2_in[4] a_12969_40175# 1.16fF
C7305 VDD a_32827_46805# 0.70fF
C7306 a_34226_59142# ctopp 3.58fF
C7307 VDD a_4443_27247# 0.40fF
C7308 a_28202_11500# ctopn 3.58fF
C7309 VDD a_43262_59142# 0.52fF
C7310 cgen.dlycontrol1_in[4] cgen.dlycontrol1_in[1] 0.82fF
C7311 a_18546_10494# a_20078_10902# 0.35fF
C7312 VDD a_25667_35253# 0.41fF
C7313 ANTENNA__1187__B1.DIODE a_13091_28327# 1.36fF
C7314 VDD a_8919_71615# 0.35fF
C7315 a_10515_15055# ANTENNA__1190__A2.DIODE 0.97fF
C7316 a_18546_16518# a_39154_16926# 0.35fF
C7317 a_28202_16520# a_29206_16520# 0.97fF
C7318 VDD a_18947_49811# 0.48fF
C7319 pmat.row_n[2] a_11067_49871# 0.46fF
C7320 VDD pmat.col[9] 4.83fF
C7321 VDD a_4298_67191# 0.31fF
C7322 VDD a_20170_61150# 0.52fF
C7323 a_32218_13508# vcm 0.65fF
C7324 a_9963_28111# a_14943_26703# 0.37fF
C7325 VDD a_18235_42359# 0.62fF
C7326 m2_48052_7214# m2_49056_7214# 0.96fF
C7327 nmat.col[10] nmat.rowoff_n[1] 0.32fF
C7328 a_30210_18528# vcm 0.65fF
C7329 VDD a_5179_20175# 0.44fF
C7330 a_5462_62215# a_10190_60663# 0.34fF
C7331 VDD a_25325_29125# 0.87fF
C7332 a_6292_65479# a_12225_74575# 0.35fF
C7333 a_4259_73807# a_4697_74005# 1.05fF
C7334 a_2648_29397# a_3576_17143# 0.41fF
C7335 VDD m3_43164_72146# 0.41fF
C7336 nmat.en_bit_n[1] nmat.col_n[15] 0.33fF
C7337 a_41254_15516# vcm 0.65fF
C7338 VDD a_26194_17524# 0.52fF
C7339 a_5363_33551# a_11067_30287# 3.46fF
C7340 pmat.rowoff_n[15] pmat.rowoff_n[4] 1.80fF
C7341 VDD m2_51064_57958# 1.02fF
C7342 pmat.row_n[12] a_14287_69455# 0.41fF
C7343 a_37238_70186# a_37238_69182# 1.00fF
C7344 VDD a_27198_8488# 0.55fF
C7345 a_20170_11500# a_20170_10496# 1.00fF
C7346 a_18546_21538# a_30118_21946# 0.35fF
C7347 VDD a_11113_36483# 2.03fF
C7348 a_26194_14512# a_26194_13508# 1.00fF
C7349 VDD a_47449_52271# 0.48fF
C7350 a_37238_23548# ctopn 3.40fF
C7351 VDD a_43262_19532# 0.52fF
C7352 a_4339_27804# a_2683_22089# 0.85fF
C7353 a_39246_9492# ctopn 3.57fF
C7354 pmat.rowoff_n[15] nmat.col_n[3] 0.57fF
C7355 a_30210_57134# a_30210_56130# 1.00fF
C7356 a_8568_26703# nmat.col[1] 3.15fF
C7357 a_34226_19532# a_35230_19532# 0.97fF
C7358 a_3866_57399# a_4985_51433# 0.67fF
C7359 a_18546_8486# vcm 0.39fF
C7360 a_37238_60146# vcm 0.62fF
C7361 VDD a_42258_10496# 0.52fF
C7362 a_15667_27239# a_7415_29397# 0.68fF
C7363 a_1781_9308# a_22365_32149# 0.60fF
C7364 a_22199_30287# a_30663_50087# 0.71fF
C7365 VDD a_6981_28879# 0.51fF
C7366 a_6787_47607# a_8491_47911# 0.53fF
C7367 a_18546_58180# a_49194_58138# 0.35fF
C7368 a_33222_10496# a_34226_10496# 0.97fF
C7369 a_18546_10494# a_49194_10902# 0.35fF
C7370 ANTENNA__1187__B1.DIODE a_17139_30503# 0.93fF
C7371 VDD a_22178_12504# 0.52fF
C7372 a_49286_62154# ctopp 3.57fF
C7373 VDD a_2879_57487# 7.96fF
C7374 a_43262_16520# vcm 0.65fF
C7375 a_12447_16143# a_9528_20407# 0.98fF
C7376 VDD a_36209_49257# 0.50fF
C7377 a_44266_56130# a_45270_56130# 0.97fF
C7378 a_11067_16359# a_6927_30503# 0.46fF
C7379 VDD a_38711_37683# 2.03fF
C7380 a_35230_13508# ctopn 3.58fF
C7381 a_30210_57134# vcm 0.62fF
C7382 VDD a_40591_38007# 0.70fF
C7383 a_29206_71190# vcm 0.60fF
C7384 a_3325_20175# clk_dig 0.89fF
C7385 a_33222_18528# ctopn 3.58fF
C7386 a_18162_64202# ctopp 1.49fF
C7387 pmat.sw a_19541_28879# 1.47fF
C7388 VDD a_12235_39913# 0.67fF
C7389 ANTENNA__1190__A2.DIODE nmat.col[19] 4.62fF
C7390 a_48282_70186# ctopp 3.57fF
C7391 a_1858_25615# nmat.sample 0.47fF
C7392 a_44266_15516# ctopn 3.58fF
C7393 a_10515_15055# nmat.col_n[1] 0.69fF
C7394 a_18823_50247# a_25850_48981# 0.52fF
C7395 VDD a_44266_11500# 0.52fF
C7396 a_26194_22544# a_27198_22544# 0.97fF
C7397 a_11067_30287# nmat.col_n[12] 1.36fF
C7398 VDD a_11619_16367# 0.48fF
C7399 VDD nmat.en_C0_n 0.37fF
C7400 ANTENNA__1197__B.DIODE nmat.en_bit_n[0] 0.40fF
C7401 a_49286_62154# a_50290_62154# 0.97fF
C7402 VDD a_5173_45993# 0.76fF
C7403 a_47278_66170# a_48282_66170# 0.97fF
C7404 a_1674_68047# a_2419_53351# 0.61fF
C7405 a_18546_69224# a_44174_69182# 0.35fF
C7406 VDD a_18162_7484# 29.42fF
C7407 a_12449_22895# a_12245_21807# 0.38fF
C7408 pmat.col_n[15] ctopp 2.04fF
C7409 VDD a_26515_35831# 0.60fF
C7410 VDD a_41162_72194# 0.32fF
C7411 a_23021_29199# nmat.col_n[7] 0.53fF
C7412 VDD a_22475_50095# 0.49fF
C7413 VDD a_4413_62037# 0.33fF
C7414 cgen.dlycontrol3_in[0] a_11041_39860# 1.62fF
C7415 a_40250_63158# a_41254_63158# 0.97fF
C7416 a_18546_16518# a_21082_16926# 0.35fF
C7417 a_41254_22544# vcm 0.65fF
C7418 a_39246_68178# ctopp 3.58fF
C7419 VDD a_48282_68178# 0.52fF
C7420 VDD a_20164_27791# 0.48fF
C7421 nmat.col_n[20] m2_39016_24282# 0.37fF
C7422 nmat.sw a_13091_18535# 2.91fF
C7423 a_4985_51433# a_6175_60039# 2.20fF
C7424 cgen.dlycontrol2_in[2] a_11497_38543# 2.30fF
C7425 VDD a_27329_42902# 1.05fF
C7426 a_24374_29941# nmat.en_bit_n[0] 0.34fF
C7427 VDD a_37827_30793# 0.98fF
C7428 VDD a_21174_56130# 0.55fF
C7429 a_18546_20534# a_50198_20942# 0.35fF
C7430 a_46274_16520# ctopn 3.58fF
C7431 VDD a_7730_69109# 0.79fF
C7432 VDD a_7370_27791# 0.59fF
C7433 a_13327_70741# a_3615_71631# 1.18fF
C7434 VDD nmat.col_n[19] 9.18fF
C7435 VDD m2_29980_7214# 0.93fF
C7436 ANTENNA__1184__B1.DIODE a_11948_49783# 2.32fF
C7437 VDD pmat.col[28] 4.45fF
C7438 a_18546_62196# a_35138_62154# 0.35fF
C7439 a_18546_66212# a_31122_66170# 0.35fF
C7440 a_18546_60188# ctopp 1.59fF
C7441 a_4075_31591# a_6467_29415# 0.68fF
C7442 a_48282_70186# a_49286_70186# 0.97fF
C7443 VDD a_24186_66170# 0.52fF
C7444 ANTENNA__1184__B1.DIODE a_30571_50959# 0.60fF
C7445 a_35230_11500# a_36234_11500# 0.97fF
C7446 a_10883_3303# a_8861_24527# 0.42fF
C7447 a_11067_64015# a_5363_33551# 2.27fF
C7448 a_37238_64162# a_37238_63158# 1.00fF
C7449 pmat.en_bit_n[0] clk_ena 2.15fF
C7450 a_5651_66975# a_1586_63927# 0.77fF
C7451 a_40250_10496# a_40250_9492# 1.00fF
C7452 a_37238_58138# a_37238_57134# 1.00fF
C7453 a_19166_60146# vcm 0.61fF
C7454 a_1591_31599# cgen.dlycontrol4_in[4] 0.68fF
C7455 a_9441_20189# a_12311_19783# 0.33fF
C7456 VDD a_11317_40188# 2.77fF
C7457 a_49286_14512# vcm 0.65fF
C7458 a_12447_16143# a_19541_28879# 0.32fF
C7459 a_10781_42364# a_12116_40871# 4.54fF
C7460 a_48282_64162# vcm 0.62fF
C7461 a_41254_60146# a_41254_59142# 1.00fF
C7462 pmat.row_n[14] nmat.en_bit_n[1] 0.37fF
C7463 a_29206_18528# a_29206_17524# 1.00fF
C7464 ANTENNA__1184__B1.DIODE ANTENNA__1190__A2.DIODE 0.58fF
C7465 VDD a_3484_58229# 0.34fF
C7466 pmat.rowoff_n[12] a_10883_3303# 1.37fF
C7467 m3_34128_24414# ctopn 0.39fF
C7468 a_1591_20181# a_1757_20181# 0.42fF
C7469 VDD a_17113_34789# 1.29fF
C7470 a_45019_38645# a_45861_29967# 0.44fF
C7471 m2_51064_62978# m2_51064_61974# 0.99fF
C7472 _1194_.B1 ANTENNA__1395__B1.DIODE 1.66fF
C7473 a_24591_28327# a_16311_28327# 0.42fF
C7474 ANTENNA__1187__B1.DIODE _1184_.A2 4.16fF
C7475 a_2791_57703# a_2727_58470# 1.99fF
C7476 a_44266_22544# ctopn 3.57fF
C7477 VDD a_49286_18528# 0.52fF
C7478 a_29206_63158# a_29206_62154# 1.00fF
C7479 a_22178_71190# m2_21948_72014# 1.00fF
C7480 VDD a_4075_49007# 0.51fF
C7481 a_45270_67174# a_46274_67174# 0.97fF
C7482 nmat.col[8] m2_26968_24282# 0.40fF
C7483 VDD a_1757_23445# 0.63fF
C7484 a_18546_70228# a_33130_70186# 0.35fF
C7485 VDD a_22178_67174# 0.52fF
C7486 nmat.col[10] a_14457_15823# 0.96fF
C7487 VDD a_11773_39087# 1.04fF
C7488 a_11921_37462# a_12513_36924# 0.38fF
C7489 a_6651_51733# a_6817_51733# 0.72fF
C7490 a_42258_66170# a_42258_65166# 1.00fF
C7491 a_35230_22544# a_35230_21540# 1.00fF
C7492 VDD a_10985_42044# 1.25fF
C7493 VDD a_2199_13887# 7.10fF
C7494 a_18546_14510# a_51202_14918# 0.35fF
C7495 a_34226_14512# a_35230_14512# 0.97fF
C7496 a_32218_62154# vcm 0.62fF
C7497 a_1781_9308# a_1923_31743# 1.28fF
C7498 a_20616_27791# a_22459_28879# 1.03fF
C7499 _1187_.A2 nmat.col[10] 4.38fF
C7500 a_33222_64162# a_34226_64162# 0.97fF
C7501 a_18546_64204# a_49194_64162# 0.35fF
C7502 a_18546_17522# a_28110_17930# 0.35fF
C7503 a_1858_25615# a_5535_29980# 1.38fF
C7504 a_18243_28327# a_10223_26703# 0.53fF
C7505 a_15667_27239# nmat.col_n[28] 0.39fF
C7506 VDD a_83677_3855# 0.35fF
C7507 a_39246_68178# a_40250_68178# 0.97fF
C7508 a_18546_57176# a_24094_57134# 0.35fF
C7509 a_12585_39355# a_11497_38543# 1.41fF
C7510 VDD a_19746_27791# 0.39fF
C7511 a_19409_40719# a_20221_40835# 0.45fF
C7512 VDD a_2315_44124# 4.02fF
C7513 a_28202_13508# a_28202_12504# 1.00fF
C7514 a_12513_39100# a_12197_38306# 1.02fF
C7515 a_1674_57711# a_6175_60039# 0.99fF
C7516 pmat.row_n[9] a_11435_58791# 0.73fF
C7517 a_18546_15514# a_28110_15922# 0.35fF
C7518 ANTENNA_fanout52_A.DIODE a_30571_50959# 1.20fF
C7519 a_47278_60146# ctopp 3.58fF
C7520 nmat.col_n[8] ctopn 2.02fF
C7521 VDD a_24833_34191# 1.91fF
C7522 a_31214_70186# vcm 0.62fF
C7523 VDD pmat.col_n[8] 5.38fF
C7524 ANTENNA__1187__B1.DIODE a_9411_2215# 0.89fF
C7525 m2_39016_24282# m3_39148_24414# 2.79fF
C7526 nmat.col_n[10] nmat.col[11] 6.61fF
C7527 a_10883_3303# nmat.sw 3.85fF
C7528 _1154_.X a_28915_50959# 0.82fF
C7529 a_2419_69455# a_2411_43301# 0.49fF
C7530 a_35186_47375# a_41926_46983# 0.45fF
C7531 a_5351_19913# a_11337_25071# 0.38fF
C7532 VDD a_35752_43781# 1.23fF
C7533 VDD a_7295_14441# 0.58fF
C7534 a_2439_13889# a_2400_13763# 0.75fF
C7535 _1179_.X a_16311_28327# 1.91fF
C7536 a_18546_59184# a_44174_59142# 0.35fF
C7537 a_35230_65166# a_35230_64162# 1.00fF
C7538 a_10873_40693# a_11071_41046# 0.30fF
C7539 a_18162_10496# ctopn 1.49fF
C7540 a_40250_57134# ctopp 3.57fF
C7541 a_39246_71190# ctopp 3.40fF
C7542 VDD a_49286_57134# 0.52fF
C7543 a_26194_58138# ctopp 3.58fF
C7544 a_22178_68178# vcm 0.62fF
C7545 VDD a_48282_71190# 0.55fF
C7546 VDD a_35230_58138# 0.52fF
C7547 a_10515_15055# _1194_.A2 0.73fF
C7548 a_1923_61759# a_2467_63125# 0.55fF
C7549 a_44266_23548# a_45270_23548# 0.97fF
C7550 cgen.enable_dlycontrol_in a_11317_36924# 0.72fF
C7551 a_19166_60146# m2_17932_59966# 0.96fF
C7552 a_29627_43983# a_30140_43781# 0.32fF
C7553 VDD a_2695_76757# 0.49fF
C7554 a_24186_16520# a_24186_15516# 1.00fF
C7555 pmat.row_n[8] vcm 1.25fF
C7556 a_41254_71190# m2_41024_72014# 1.00fF
C7557 pmat.row_n[7] cgen.dlycontrol4_in[1] 2.25fF
C7558 VDD m2_17932_60970# 1.00fF
C7559 a_46274_9492# a_47278_9492# 0.97fF
C7560 pmat.rowon_n[8] a_10515_13967# 0.99fF
C7561 _1154_.X ANTENNA__1395__B1.DIODE 0.82fF
C7562 a_19166_70186# a_19166_69182# 1.00fF
C7563 VDD a_8789_60431# 0.39fF
C7564 a_2263_43719# a_11711_50959# 0.43fF
C7565 pmat.rowoff_n[15] vcm 0.81fF
C7566 m2_30984_7214# m3_31116_7346# 2.79fF
C7567 a_18546_24550# a_49194_24958# 0.35fF
C7568 inn_analog nmat.col_n[24] 0.57fF
C7569 VDD a_27895_41001# 0.62fF
C7570 VDD a_37813_39867# 1.58fF
C7571 nmat.col[5] vcm 5.76fF
C7572 a_27198_23548# vcm 0.65fF
C7573 nmat.col[20] nmat.col_n[19] 6.61fF
C7574 a_38851_28327# a_43533_30761# 0.63fF
C7575 a_25695_28111# a_35244_32411# 0.53fF
C7576 a_29206_9492# vcm 0.65fF
C7577 VDD a_27198_69182# 0.52fF
C7578 a_18546_12502# a_18162_12504# 2.61fF
C7579 a_24591_28327# a_25315_28335# 0.75fF
C7580 a_18546_22542# a_46182_22950# 0.35fF
C7581 VDD config_1_in[0] 1.30fF
C7582 a_19166_20536# ctopn 3.43fF
C7583 VDD a_19417_43990# 1.01fF
C7584 a_2021_26677# a_2411_33749# 2.44fF
C7585 a_6283_31591# a_6007_33767# 0.39fF
C7586 a_1781_9308# a_35244_32411# 0.47fF
C7587 VDD m2_27972_24282# 0.62fF
C7588 a_45270_20536# vcm 0.65fF
C7589 a_7658_71543# a_3615_71631# 0.49fF
C7590 nmat.sw a_10873_36341# 1.43fF
C7591 a_36234_65166# a_37238_65166# 0.97fF
C7592 a_27198_59142# ctopp 3.58fF
C7593 VDD nmat.col_n[16] 5.05fF
C7594 a_21174_11500# ctopn 3.58fF
C7595 VDD a_20616_27791# 3.10fF
C7596 nmat.col[16] a_35230_24552# 0.38fF
C7597 VDD a_19579_52789# 0.46fF
C7598 VDD a_36234_59142# 0.52fF
C7599 a_43262_21540# a_44266_21540# 0.97fF
C7600 a_18162_69222# vcm 6.95fF
C7601 a_10441_21263# nmat.col_n[3] 1.60fF
C7602 a_4128_64391# a_6559_33767# 0.35fF
C7603 a_11435_58791# a_19541_28879# 6.08fF
C7604 a_18546_16518# a_32126_16926# 0.35fF
C7605 m2_51064_22274# m3_51196_22406# 2.76fF
C7606 a_1591_31599# config_2_in[11] 0.92fF
C7607 pmat.row_n[10] a_18162_66210# 25.57fF
C7608 nmat.rowon_n[14] a_1586_8439# 1.08fF
C7609 a_44266_71190# a_44266_70186# 1.00fF
C7610 a_10883_3303# a_1858_25615# 0.88fF
C7611 a_25190_13508# vcm 0.65fF
C7612 a_24374_29941# a_16478_29423# 0.81fF
C7613 nmat.col[26] nmat.col_n[24] 0.61fF
C7614 a_9963_13967# nmat.rowon_n[2] 0.68fF
C7615 m2_41024_7214# m2_42028_7214# 0.96fF
C7616 a_19166_68178# m2_17932_67998# 0.96fF
C7617 cgen.dlycontrol3_in[4] a_12237_38772# 0.50fF
C7618 pmat.col_n[26] _1192_.A2 0.45fF
C7619 pmat.row_n[15] a_3351_27249# 0.71fF
C7620 a_23182_18528# vcm 0.65fF
C7621 nmat.sw cgen.dlycontrol1_in[3] 0.58fF
C7622 a_39079_40947# a_39413_40956# 0.34fF
C7623 m2_51064_67998# vcm 0.51fF
C7624 a_21739_29415# a_11711_50959# 1.50fF
C7625 a_9581_56079# a_12003_52815# 0.42fF
C7626 m2_51064_18258# m2_51064_17254# 0.99fF
C7627 a_42258_13508# a_43262_13508# 0.97fF
C7628 a_6283_31591# a_32771_31599# 0.36fF
C7629 a_34226_15516# vcm 0.65fF
C7630 a_10873_39605# cgen.dlycontrol2_in[3] 2.49fF
C7631 VDD a_21647_51183# 0.48fF
C7632 _1196_.B1 ANTENNA__1195__A1.DIODE 3.83fF
C7633 nmat.col_n[21] ctopn 2.04fF
C7634 VDD a_13643_29415# 8.07fF
C7635 a_33222_63158# pmat.col[14] 0.31fF
C7636 a_25879_31591# nmat.col_n[26] 1.16fF
C7637 m2_22952_72014# m3_23084_72146# 2.79fF
C7638 a_40250_18528# a_41254_18528# 0.97fF
C7639 VDD a_5391_32900# 0.42fF
C7640 _1187_.A2 _1183_.A2 5.59fF
C7641 a_11149_36924# a_10873_36341# 1.92fF
C7642 a_18546_21538# a_23090_21946# 0.35fF
C7643 VDD a_9375_72007# 0.53fF
C7644 a_27198_62154# a_27198_61150# 1.00fF
C7645 a_18162_63198# ctopp 1.49fF
C7646 a_30210_23548# ctopn 3.40fF
C7647 VDD a_36234_19532# 0.52fF
C7648 m2_48052_54946# m3_48184_55078# 2.79fF
C7649 a_32218_9492# ctopn 3.57fF
C7650 VDD m2_47048_72014# 1.40fF
C7651 cgen.dlycontrol3_in[3] cgen.dlycontrol2_in[4] 1.15fF
C7652 nmat.col_n[13] m2_31988_24282# 0.38fF
C7653 pmat.col_n[31] a_50290_56130# 0.33fF
C7654 a_30210_60146# vcm 0.62fF
C7655 VDD a_35230_10496# 0.52fF
C7656 VDD a_40591_39095# 0.70fF
C7657 a_19584_52423# a_20475_49783# 0.42fF
C7658 a_10515_15055# pmat.rowoff_n[9] 1.03fF
C7659 a_48282_20536# ctopn 3.58fF
C7660 VDD a_1591_43029# 0.41fF
C7661 a_11041_40948# a_10873_40693# 1.32fF
C7662 a_27198_15516# a_27198_14512# 1.00fF
C7663 VDD a_40467_46261# 0.35fF
C7664 VDD a_16083_50069# 2.68fF
C7665 a_18243_28327# a_13091_28327# 5.88fF
C7666 VDD a_34134_55126# 0.38fF
C7667 a_18546_58180# a_42166_58138# 0.35fF
C7668 VDD nmat.en_bit_n[0] 3.68fF
C7669 a_29206_69182# a_29206_68178# 1.00fF
C7670 a_2999_76922# a_2861_76757# 0.71fF
C7671 a_18546_10494# a_42166_10902# 0.35fF
C7672 a_37238_21540# a_37238_20536# 1.00fF
C7673 inn_analog ctopn 3.40fF
C7674 a_42258_62154# ctopp 3.58fF
C7675 VDD comp.adc_comp_circuit_0.adc_comp_buffer_1.in 0.44fF
C7676 a_36234_16520# vcm 0.65fF
C7677 a_12197_43746# cgen.dlycontrol4_in[1] 0.38fF
C7678 m2_17932_22274# vcm 0.44fF
C7679 a_14641_57711# pmat.rowoff_n[5] 0.59fF
C7680 VDD a_20627_38825# 0.64fF
C7681 a_28202_13508# ctopn 3.58fF
C7682 VDD a_19166_9492# 0.56fF
C7683 a_14712_37429# a_16981_37462# 1.10fF
C7684 a_23182_57134# vcm 0.62fF
C7685 VDD a_26501_37462# 1.14fF
C7686 a_2411_43301# cgen.dlycontrol4_in[3] 0.34fF
C7687 a_22178_71190# vcm 0.60fF
C7688 a_26194_18528# ctopn 3.58fF
C7689 a_9963_13967# comp_latch 0.38fF
C7690 _1187_.A2 a_34204_27765# 0.95fF
C7691 a_19166_64162# a_19166_63158# 1.00fF
C7692 a_41254_70186# ctopp 3.57fF
C7693 VDD a_2124_55107# 0.57fF
C7694 a_37238_15516# ctopn 3.58fF
C7695 VDD a_50290_70186# 0.54fF
C7696 VDD a_37238_11500# 0.52fF
C7697 a_48282_23548# a_48282_22544# 1.00fF
C7698 pmat.col_n[23] a_16311_28327# 0.82fF
C7699 a_40837_46261# a_44389_40553# 0.38fF
C7700 VDD a_12175_27221# 1.03fF
C7701 VDD m2_23956_54946# 0.62fF
C7702 a_5179_31591# a_7939_31591# 2.44fF
C7703 a_24407_31375# a_25879_31591# 2.54fF
C7704 a_47278_60146# a_48282_60146# 0.97fF
C7705 a_3576_17143# a_5266_17143# 0.57fF
C7706 a_2835_13077# a_10839_11989# 0.46fF
C7707 a_18546_69224# a_37146_69182# 0.35fF
C7708 VDD a_30278_30511# 2.31fF
C7709 VDD pmat.rowoff_n[6] 2.34fF
C7710 nmat.col[18] vcm 14.43fF
C7711 a_12513_36924# a_14589_35286# 3.32fF
C7712 nmat.col[26] ctopn 1.98fF
C7713 a_31214_11500# a_31214_10496# 1.00fF
C7714 VDD a_5271_35407# 0.78fF
C7715 a_1769_13103# config_2_in[13] 0.33fF
C7716 VDD a_7165_13353# 0.33fF
C7717 VDD a_9135_62613# 0.47fF
C7718 a_34226_22544# vcm 0.65fF
C7719 a_36234_61150# a_37238_61150# 0.97fF
C7720 a_32218_68178# ctopp 3.58fF
C7721 ANTENNA__1395__B1.DIODE nmat.col_n[7] 0.39fF
C7722 VDD a_41254_68178# 0.52fF
C7723 a_21174_12504# a_21174_11500# 1.00fF
C7724 pmat.col_n[10] vcm 2.80fF
C7725 a_10873_40693# a_12197_41570# 2.77fF
C7726 a_48282_63158# vcm 0.62fF
C7727 a_16311_28327# nmat.col[7] 1.60fF
C7728 pmat.row_n[7] _1196_.B1 0.30fF
C7729 _1194_.A2 ANTENNA__1184__B1.DIODE 0.68fF
C7730 ANTENNA__1395__A1.DIODE _1187_.A2 2.02fF
C7731 ANTENNA__1197__A.DIODE ANTENNA__1197__B.DIODE 1.55fF
C7732 a_18243_28327# a_17139_30503# 1.12fF
C7733 pmat.rowoff_n[7] a_2283_39189# 0.42fF
C7734 VDD a_9581_56079# 2.30fF
C7735 a_30210_20536# a_31214_20536# 0.97fF
C7736 a_18546_20534# a_43170_20942# 0.35fF
C7737 a_39246_16520# ctopn 3.58fF
C7738 VDD a_14641_57167# 1.06fF
C7739 m2_51064_19262# a_50290_19532# 0.96fF
C7740 pmat.col[25] ctopp 1.97fF
C7741 VDD a_5497_73719# 1.27fF
C7742 a_18546_62196# a_28110_62154# 0.35fF
C7743 a_18546_66212# a_24094_66170# 0.35fF
C7744 a_43262_67174# a_43262_66170# 1.00fF
C7745 a_29206_9492# a_29206_8488# 1.00fF
C7746 VDD a_46274_23548# 0.55fF
C7747 VDD a_48282_9492# 0.52fF
C7748 a_11921_37462# a_12309_36483# 0.40fF
C7749 a_18546_11498# a_46182_11906# 0.35fF
C7750 VDD a_46229_37583# 1.09fF
C7751 pmat.rowon_n[11] a_10239_14183# 0.35fF
C7752 pmat.row_n[5] a_18162_61190# 25.57fF
C7753 a_42258_56130# m2_42028_54946# 0.99fF
C7754 ANTENNA__1197__A.DIODE a_31675_47695# 0.38fF
C7755 a_9785_28879# a_7415_29397# 0.31fF
C7756 a_42258_17524# a_43262_17524# 0.97fF
C7757 pmat.sample_n a_16083_50069# 0.44fF
C7758 a_40250_57134# a_41254_57134# 0.97fF
C7759 ANTENNA__1395__B1.DIODE a_40837_46261# 1.70fF
C7760 a_45270_20536# a_45270_19532# 1.00fF
C7761 a_39246_71190# a_40250_71190# 0.97fF
C7762 a_13091_28327# a_12851_28853# 1.27fF
C7763 a_2007_25597# a_5351_19913# 0.41fF
C7764 VDD a_46705_38671# 0.65fF
C7765 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col[26] 1.01fF
C7766 a_26194_58138# a_27198_58138# 0.97fF
C7767 VDD a_10781_42869# 7.26fF
C7768 a_42258_14512# vcm 0.65fF
C7769 a_41254_64162# vcm 0.62fF
C7770 pmat.row_n[7] a_3659_39733# 0.34fF
C7771 VDD pmat.col[20] 4.44fF
C7772 a_43262_8488# a_44266_8488# 0.97fF
C7773 VDD a_10953_34951# 1.18fF
C7774 VDD a_13102_71311# 1.18fF
C7775 a_6283_31591# cgen.dlycontrol3_in[3] 1.39fF
C7776 VDD a_44266_13508# 0.52fF
C7777 pmat.col_n[10] pmat.col[10] 0.74fF
C7778 a_37238_22544# ctopn 3.57fF
C7779 VDD a_42258_18528# 0.52fF
C7780 m2_32992_24282# vcm 0.42fF
C7781 a_26194_61150# a_26194_60146# 1.00fF
C7782 a_34226_19532# a_34226_18528# 1.00fF
C7783 a_18546_70228# a_26102_70186# 0.35fF
C7784 VDD a_9643_66389# 1.09fF
C7785 _1184_.A2 a_83196_3561# 0.32fF
C7786 a_10071_17999# a_4976_16091# 0.34fF
C7787 a_1781_9308# a_7619_30485# 0.94fF
C7788 a_2683_22089# a_2191_25045# 0.38fF
C7789 a_9777_26935# a_9217_23983# 0.52fF
C7790 a_18546_14510# a_44174_14918# 0.35fF
C7791 a_25190_62154# vcm 0.62fF
C7792 a_13091_52047# a_33423_47695# 0.74fF
C7793 a_2315_44124# a_3417_47919# 0.51fF
C7794 a_6927_30503# a_9595_30511# 0.62fF
C7795 a_18546_64204# a_42166_64162# 0.35fF
C7796 a_2835_13077# a_9583_10121# 0.48fF
C7797 VDD a_20439_27247# 0.75fF
C7798 a_4991_69831# a_1957_43567# 0.35fF
C7799 a_20534_35431# cgen.dlycontrol1_in[0] 1.07fF
C7800 a_27198_59142# a_27198_58138# 1.00fF
C7801 VDD a_4659_53738# 1.25fF
C7802 a_31214_8488# m2_30984_7214# 1.00fF
C7803 a_2149_45717# pmat.rowon_n[3] 1.57fF
C7804 nmat.col_n[10] ctopn 2.02fF
C7805 a_50290_13508# m2_51064_13238# 0.96fF
C7806 a_50290_60146# m2_51064_59966# 0.96fF
C7807 a_44266_65166# vcm 0.62fF
C7808 _1187_.A2 ANTENNA__1395__A2.DIODE 0.64fF
C7809 a_40250_60146# ctopp 3.58fF
C7810 clk_ena ctopn 0.89fF
C7811 a_18546_69224# a_18162_69222# 2.62fF
C7812 VDD a_10764_32117# 0.65fF
C7813 VDD a_49286_60146# 0.52fF
C7814 VDD a_14113_36604# 1.28fF
C7815 a_24186_70186# vcm 0.62fF
C7816 a_11019_71543# a_11115_71285# 1.97fF
C7817 a_1899_35051# a_1823_68565# 2.49fF
C7818 a_13479_26935# a_14365_22351# 0.55fF
C7819 a_32218_17524# a_32218_16520# 1.00fF
C7820 a_30663_50087# a_41731_49525# 3.39fF
C7821 a_45270_14512# ctopn 3.58fF
C7822 a_38242_12504# a_39246_12504# 0.97fF
C7823 pmat.sample pmat.row_n[14] 0.52fF
C7824 a_2411_16101# a_3688_17179# 0.36fF
C7825 a_10515_61839# pmat.rowoff_n[9] 0.47fF
C7826 VDD a_22357_43493# 1.27fF
C7827 VDD a_9319_15279# 0.44fF
C7828 VDD a_16478_29423# 3.55fF
C7829 a_35230_55126# ctopp 1.70fF
C7830 a_18546_59184# pmat.rowoff_n[3] 4.09fF
C7831 a_27198_59142# a_28202_59142# 0.97fF
C7832 a_18546_59184# a_37146_59142# 0.35fF
C7833 pmat.row_n[7] a_18546_63200# 0.35fF
C7834 pmat.rowon_n[7] a_18162_63198# 1.19fF
C7835 cgen.dlycontrol2_in[3] cgen.dlycontrol2_in[2] 1.29fF
C7836 a_1858_25615# a_7717_14735# 0.35fF
C7837 m2_17932_71010# vcm 0.42fF
C7838 a_33222_57134# ctopp 3.57fF
C7839 a_4075_68583# a_3923_68021# 0.58fF
C7840 a_11837_68591# pmat.rowoff_n[12] 0.48fF
C7841 VDD a_6664_26159# 5.39fF
C7842 a_32218_71190# ctopp 3.40fF
C7843 VDD a_42258_57134# 0.52fF
C7844 VDD a_35382_34191# 0.53fF
C7845 a_26891_28327# a_28704_29568# 0.37fF
C7846 a_33467_46261# a_32687_46607# 1.28fF
C7847 a_24867_53135# pmat.col[7] 0.36fF
C7848 ANTENNA__1190__A1.DIODE a_28915_50959# 1.70fF
C7849 VDD a_41254_71190# 0.55fF
C7850 a_20170_24552# m2_20944_24282# 0.96fF
C7851 VDD a_28202_58138# 0.52fF
C7852 VDD a_1739_47893# 5.74fF
C7853 VDD a_3891_60431# 0.39fF
C7854 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top a_52398_39208# 0.73fF
C7855 cgen.dlycontrol4_in[2] a_1923_31743# 0.31fF
C7856 VDD a_18235_41271# 0.62fF
C7857 pmat.row_n[4] a_3576_17143# 1.65fF
C7858 m2_17932_10226# vcm 0.44fF
C7859 a_18546_24550# a_42166_24958# 0.35fF
C7860 a_50290_68178# m2_51064_67998# 0.96fF
C7861 a_28704_29568# a_40969_30287# 0.32fF
C7862 VDD a_19509_39638# 1.08fF
C7863 pmat.rowon_n[11] ctopn 0.60fF
C7864 a_23182_68178# a_23182_67174# 1.00fF
C7865 a_50290_8488# m2_50060_7214# 1.00fF
C7866 a_22178_9492# vcm 0.65fF
C7867 VDD a_20170_69182# 0.52fF
C7868 a_44266_61150# vcm 0.62fF
C7869 _1154_.X _1192_.B1 0.82fF
C7870 a_41254_23548# m2_41024_24282# 0.99fF
C7871 a_12585_39355# a_14712_37429# 1.44fF
C7872 _1194_.B1 a_46027_44905# 0.66fF
C7873 ANTENNA__1190__A1.DIODE ANTENNA__1395__B1.DIODE 14.72fF
C7874 a_24591_28327# a_24407_31375# 0.52fF
C7875 a_18546_22542# a_39154_22950# 0.35fF
C7876 VDD a_10651_44211# 1.00fF
C7877 VDD a_27763_27221# 1.08fF
C7878 _1224_.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.34fF
C7879 VDD m2_47048_54946# 0.62fF
C7880 a_17139_30503# a_30571_50959# 1.25fF
C7881 a_38242_20536# vcm 0.65fF
C7882 a_20170_59142# ctopp 3.57fF
C7883 VDD a_29206_59142# 0.52fF
C7884 a_18243_28327# a_9411_2215# 0.46fF
C7885 pmat.col_n[18] ctopp 2.02fF
C7886 a_21371_50087# a_25695_28111# 0.87fF
C7887 VDD a_44174_72194# 0.32fF
C7888 _1154_.A a_24867_53135# 0.34fF
C7889 a_50290_17524# vcm 0.65fF
C7890 a_19166_22544# ctopn 3.24fF
C7891 cgen.dlycontrol4_in[4] a_11317_40188# 1.65fF
C7892 a_21174_16520# a_22178_16520# 0.97fF
C7893 a_18546_16518# a_25098_16926# 0.35fF
C7894 m2_28976_54946# vcm 0.42fF
C7895 a_4955_40277# cgen.dlycontrol4_in[0] 0.30fF
C7896 a_19166_9492# a_20170_9492# 0.97fF
C7897 VDD a_12061_26703# 2.17fF
C7898 VDD a_1643_61493# 0.38fF
C7899 a_2327_11477# a_2493_11477# 0.72fF
C7900 VDD a_37960_42693# 1.12fF
C7901 _1187_.A2 a_41926_46983# 0.41fF
C7902 ANTENNA__1395__A2.DIODE pmat.col[1] 1.05fF
C7903 m2_33996_7214# m2_35000_7214# 0.96fF
C7904 a_17139_30503# ANTENNA__1190__A2.DIODE 3.74fF
C7905 pmat.row_n[5] pmat.row_n[2] 0.47fF
C7906 a_10239_14183# a_12447_16143# 0.35fF
C7907 VDD a_5417_11445# 0.55fF
C7908 a_18546_72236# a_21082_72194# 0.35fF
C7909 VDD nmat.col[27] 4.36fF
C7910 a_17139_30503# a_44811_36469# 1.02fF
C7911 a_27198_15516# vcm 0.65fF
C7912 VDD a_12520_51451# 0.55fF
C7913 cgen.dlycontrol2_in[1] a_26583_34343# 1.20fF
C7914 VDD a_8197_20871# 1.14fF
C7915 a_18162_66210# ctopp 1.49fF
C7916 a_30210_70186# a_30210_69182# 1.00fF
C7917 VDD a_14071_8511# 0.35fF
C7918 pmat.row_n[0] vcm 1.14fF
C7919 m2_17932_65990# m2_17932_64986# 0.99fF
C7920 a_46274_12504# vcm 0.65fF
C7921 pmat.en_bit_n[0] a_15753_28879# 0.78fF
C7922 a_23182_23548# ctopn 3.40fF
C7923 pmat.col[14] vcm 5.88fF
C7924 VDD a_29206_19532# 0.52fF
C7925 cgen.enable_dlycontrol_in a_12069_38517# 1.40fF
C7926 a_25190_9492# ctopn 3.57fF
C7927 VDD m2_32992_72014# 0.98fF
C7928 a_23182_57134# a_23182_56130# 1.00fF
C7929 _1192_.B1 pmat.col[2] 0.52fF
C7930 _1179_.X a_24407_31375# 0.80fF
C7931 _1192_.A2 a_15667_27239# 0.45fF
C7932 a_27198_19532# a_28202_19532# 0.97fF
C7933 a_23182_60146# vcm 0.62fF
C7934 VDD a_28202_10496# 0.52fF
C7935 a_3746_58487# cgen.dlycontrol4_in[5] 1.32fF
C7936 pmat.rowon_n[3] a_14195_7351# 1.92fF
C7937 cgen.dlycontrol2_in[3] a_11339_39319# 3.92fF
C7938 VDD a_25117_39141# 1.33fF
C7939 a_34705_51959# a_25695_28111# 0.68fF
C7940 a_41254_20536# ctopn 3.58fF
C7941 VDD cgen.dlycontrol4_in[0] 7.23fF
C7942 a_18546_59184# a_18162_59182# 2.62fF
C7943 pmat.col[10] m2_28976_54946# 0.39fF
C7944 a_18546_58180# a_35138_58138# 0.35fF
C7945 a_18546_10494# a_35138_10902# 0.35fF
C7946 a_26194_10496# a_27198_10496# 0.97fF
C7947 VDD a_11711_12565# 0.44fF
C7948 a_35230_62154# ctopp 3.58fF
C7949 VDD a_44266_62154# 0.52fF
C7950 VDD m2_51064_12234# 1.02fF
C7951 a_29206_16520# vcm 0.65fF
C7952 a_30571_50959# a_26891_28327# 0.78fF
C7953 pmat.row_n[11] nmat.rowon_n[1] 0.40fF
C7954 a_18823_50247# a_20475_49783# 0.52fF
C7955 pmat.sw a_10147_29415# 0.85fF
C7956 VDD a_16219_49007# 0.46fF
C7957 a_37238_56130# a_38242_56130# 0.97fF
C7958 VDD a_6639_23413# 0.43fF
C7959 VDD a_5659_38127# 0.36fF
C7960 a_21174_13508# ctopn 3.58fF
C7961 ANTENNA__1196__A2.DIODE pmat.col[1] 0.37fF
C7962 VDD a_20535_40183# 0.65fF
C7963 a_13597_37571# a_16981_37462# 0.65fF
C7964 VDD a_11261_37981# 1.34fF
C7965 _1194_.A2 nmat.col_n[29] 10.81fF
C7966 a_18162_18528# ctopn 1.49fF
C7967 VDD a_14149_39747# 1.40fF
C7968 VDD rst_n 1.52fF
C7969 a_2983_48071# a_4313_44111# 0.49fF
C7970 a_11435_58791# a_4703_24527# 0.40fF
C7971 a_6007_33767# nmat.col_n[12] 1.45fF
C7972 a_34226_70186# ctopp 3.57fF
C7973 VDD ANTENNA__1197__A.DIODE 14.23fF
C7974 a_30210_15516# ctopn 3.58fF
C7975 VDD a_43262_70186# 0.52fF
C7976 VDD a_30210_11500# 0.52fF
C7977 a_18546_22542# a_21082_22950# 0.35fF
C7978 _1184_.A2 a_2046_30184# 0.90fF
C7979 a_24591_28327# a_17842_27497# 1.11fF
C7980 a_49286_16520# a_49286_15516# 1.00fF
C7981 a_42258_62154# a_43262_62154# 0.97fF
C7982 pmat.rowon_n[8] nmat.sw 0.60fF
C7983 pmat.rowoff_n[7] cgen.dlycontrol4_in[1] 2.38fF
C7984 a_40250_66170# a_41254_66170# 0.97fF
C7985 VDD clk_comp 2.49fF
C7986 a_20170_20536# vcm 0.65fF
C7987 a_49286_12504# ctopn 3.57fF
C7988 a_18546_69224# a_30118_69182# 0.35fF
C7989 a_3351_27249# a_4068_25615# 0.72fF
C7990 a_45270_56130# vcm 0.62fF
C7991 VDD pmat.col_n[11] 5.13fF
C7992 a_10147_29415# a_27001_30511# 0.31fF
C7993 cgen.dlycontrol4_in[4] a_19417_43990# 0.77fF
C7994 a_18546_63200# a_49194_63158# 0.35fF
C7995 a_33222_63158# a_34226_63158# 0.97fF
C7996 m2_44036_24282# m3_44168_24414# 2.79fF
C7997 a_27198_22544# vcm 0.65fF
C7998 a_25190_68178# ctopp 3.58fF
C7999 _1194_.B1 a_30663_50087# 0.74fF
C8000 VDD config_2_in[15] 0.89fF
C8001 a_7415_29397# a_8861_24527# 0.37fF
C8002 a_48282_66170# vcm 0.62fF
C8003 VDD a_34226_68178# 0.52fF
C8004 pmat.col[13] m2_31988_54946# 0.40fF
C8005 a_17163_50857# a_10883_3303# 0.33fF
C8006 pmat.rowoff_n[4] a_10883_3303# 0.32fF
C8007 VDD a_46013_42997# 0.64fF
C8008 a_41254_63158# vcm 0.62fF
C8009 _1184_.A2 ANTENNA__1190__A2.DIODE 2.49fF
C8010 ANTENNA__1190__B1.DIODE nmat.rowoff_n[1] 0.38fF
C8011 ANTENNA__1195__A1.DIODE pmat.col[12] 0.46fF
C8012 a_14287_69455# pmat.rowoff_n[13] 0.53fF
C8013 a_18546_20534# a_36142_20942# 0.35fF
C8014 a_32218_16520# ctopn 3.58fF
C8015 VDD result_out[8] 0.78fF
C8016 a_11948_49783# a_9411_2215# 2.84fF
C8017 pmat.rowoff_n[12] pmat.row_n[7] 0.40fF
C8018 a_10883_3303# nmat.col_n[3] 4.45fF
C8019 a_18546_62196# a_21082_62154# 0.35fF
C8020 a_18162_58178# ctopp 1.49fF
C8021 VDD a_39647_48767# 0.34fF
C8022 a_20616_27791# nmat.col_n[2] 0.60fF
C8023 VDD a_39246_23548# 0.55fF
C8024 a_41254_70186# a_42258_70186# 0.97fF
C8025 a_25879_31591# a_26479_32117# 2.80fF
C8026 VDD a_10921_64786# 2.51fF
C8027 VDD a_41254_9492# 0.52fF
C8028 a_24407_31375# pmat.col[0] 0.76fF
C8029 a_28202_11500# a_29206_11500# 0.97fF
C8030 a_18546_11498# a_39154_11906# 0.35fF
C8031 a_2021_11043# a_8481_10396# 0.31fF
C8032 nmat.sample vcm 15.34fF
C8033 VDD a_22393_37692# 1.36fF
C8034 a_10239_14183# a_11435_58791# 2.51fF
C8035 pmat.row_n[10] a_18162_18528# 25.57fF
C8036 m2_36004_7214# m3_36136_7346# 2.79fF
C8037 a_1769_13103# config_1_in[15] 0.49fF
C8038 a_30210_64162# a_30210_63158# 1.00fF
C8039 pmat.row_n[13] pmat.row_n[2] 10.90fF
C8040 a_33222_10496# a_33222_9492# 1.00fF
C8041 a_1899_35051# a_4955_40277# 0.39fF
C8042 a_18546_19530# a_18162_19532# 2.61fF
C8043 a_46274_67174# vcm 0.62fF
C8044 a_30210_58138# a_30210_57134# 1.00fF
C8045 VDD a_11051_8903# 0.70fF
C8046 VDD a_19439_50095# 0.32fF
C8047 a_7693_22365# a_7644_16341# 1.56fF
C8048 inn_analog ctopp 0.99fF
C8049 a_13091_7655# a_12981_8213# 0.38fF
C8050 VDD a_26331_44535# 0.63fF
C8051 a_35230_14512# vcm 0.65fF
C8052 VDD a_19166_16520# 0.58fF
C8053 a_5351_19913# a_7026_24527# 1.33fF
C8054 a_6787_47607# a_4991_69831# 2.84fF
C8055 a_34226_64162# vcm 0.62fF
C8056 VDD m2_37008_24282# 0.61fF
C8057 a_34226_60146# a_34226_59142# 1.00fF
C8058 a_9411_2215# ANTENNA__1190__A2.DIODE 2.37fF
C8059 a_22178_18528# a_22178_17524# 1.00fF
C8060 a_2046_30184# a_7939_31591# 0.93fF
C8061 a_12069_38517# a_12228_39605# 0.37fF
C8062 _1192_.B1 a_40837_46261# 1.15fF
C8063 a_11927_27399# nmat.col_n[1] 0.36fF
C8064 a_12061_26703# a_12449_22895# 0.34fF
C8065 a_19166_9492# m2_17932_9222# 0.96fF
C8066 VDD a_1591_69679# 1.12fF
C8067 VDD a_37238_13508# 0.52fF
C8068 pmat.col_n[19] _1196_.B1 0.48fF
C8069 a_3615_71631# a_4075_31591# 0.86fF
C8070 a_5363_70543# a_10055_31591# 0.71fF
C8071 a_30210_22544# ctopn 3.57fF
C8072 ANTENNA__1195__A1.DIODE a_22199_30287# 0.57fF
C8073 VDD a_35230_18528# 0.52fF
C8074 a_22178_63158# a_22178_62154# 1.00fF
C8075 a_38242_67174# a_39246_67174# 0.97fF
C8076 a_4955_40277# a_6554_43255# 0.48fF
C8077 a_5351_19913# a_7533_19087# 0.48fF
C8078 a_6664_26159# a_7840_27247# 0.60fF
C8079 a_5651_66975# a_12107_62037# 0.77fF
C8080 a_35230_66170# a_35230_65166# 1.00fF
C8081 a_28202_22544# a_28202_21540# 1.00fF
C8082 VDD a_13561_42333# 1.32fF
C8083 VDD a_46274_15516# 0.52fF
C8084 a_18546_14510# a_37146_14918# 0.35fF
C8085 a_27198_14512# a_28202_14512# 0.97fF
C8086 pmat.row_n[15] a_10814_29111# 0.34fF
C8087 a_25695_28111# a_37820_30485# 0.32fF
C8088 VDD a_1591_20181# 0.39fF
C8089 a_26194_64162# a_27198_64162# 0.97fF
C8090 a_18546_64204# a_35138_64162# 0.35fF
C8091 a_32218_68178# a_33222_68178# 0.97fF
C8092 a_21174_13508# a_21174_12504# 1.00fF
C8093 a_18546_21538# ctopn 1.59fF
C8094 VDD a_1899_35051# 11.36fF
C8095 a_37238_65166# vcm 0.62fF
C8096 a_44266_21540# vcm 0.65fF
C8097 a_33222_60146# ctopp 3.58fF
C8098 m2_27972_72014# m3_28104_72146# 2.79fF
C8099 VDD a_45119_32661# 0.45fF
C8100 VDD a_42258_60146# 0.52fF
C8101 pmat.col_n[0] ctopp 1.81fF
C8102 cgen.dlycontrol2_in[0] a_11681_35823# 0.37fF
C8103 VDD a_2419_53351# 9.28fF
C8104 a_4128_64391# a_9581_56079# 1.41fF
C8105 VDD a_7645_53909# 0.69fF
C8106 a_9595_30511# a_9761_30511# 0.39fF
C8107 pmat.row_n[13] a_18162_21540# 25.57fF
C8108 m2_18936_24282# m3_19068_24414# 2.79fF
C8109 a_11883_62063# a_11797_60431# 1.70fF
C8110 ANTENNA__1197__A.DIODE pmat.rowoff_n[1] 1.91fF
C8111 a_18546_19530# a_48190_19938# 0.35fF
C8112 a_38242_14512# ctopn 3.58fF
C8113 _1224_.X a_21371_50087# 0.57fF
C8114 a_31339_31787# nmat.col[29] 0.48fF
C8115 pmat.rowon_n[10] pmat.row_n[7] 0.84fF
C8116 a_24407_31375# nmat.sample_n 1.64fF
C8117 VDD a_48282_16520# 0.52fF
C8118 a_18546_59184# a_30118_59142# 0.35fF
C8119 a_28202_65166# a_28202_64162# 1.00fF
C8120 a_26194_57134# ctopp 3.57fF
C8121 VDD a_20895_30199# 0.51fF
C8122 nmat.rowon_n[7] a_4976_16091# 1.35fF
C8123 VDD a_9655_6335# 0.39fF
C8124 ANTENNA__1196__A2.DIODE a_13275_48783# 0.60fF
C8125 a_25190_71190# ctopp 3.40fF
C8126 VDD a_35230_57134# 0.52fF
C8127 VDD a_34226_71190# 0.55fF
C8128 cgen.dlycontrol3_in[3] a_4128_46983# 1.05fF
C8129 VDD a_18546_12502# 32.63fF
C8130 VDD a_21174_58138# 0.52fF
C8131 a_37238_23548# a_38242_23548# 0.97fF
C8132 nmat.col_n[14] ctopn 2.02fF
C8133 a_39246_9492# a_40250_9492# 0.97fF
C8134 a_2407_49289# pmat.rowoff_n[7] 0.88fF
C8135 a_38851_28327# a_37291_29397# 1.65fF
C8136 a_9135_60967# pmat.rowon_n[3] 0.56fF
C8137 a_18546_18526# a_20078_18934# 0.35fF
C8138 a_16981_37462# a_19928_37253# 0.66fF
C8139 a_14712_37429# a_21219_36885# 0.47fF
C8140 a_46274_12504# a_46274_11500# 1.00fF
C8141 a_18546_11498# a_21082_11906# 0.35fF
C8142 VDD a_32035_38007# 0.66fF
C8143 _1194_.A2 a_17139_30503# 0.45fF
C8144 a_25190_56130# m2_24960_54946# 0.99fF
C8145 pmat.row_n[15] nmat.rowon_n[7] 1.74fF
C8146 a_18546_55168# a_46182_55126# 0.35fF
C8147 a_18546_24550# a_35138_24958# 0.39fF
C8148 nmat.col_n[31] nmat.col[28] 0.50fF
C8149 nmat.col_n[30] nmat.col[21] 2.97fF
C8150 a_1591_33775# a_1757_33775# 0.69fF
C8151 a_37238_61150# vcm 0.62fF
C8152 a_9411_2215# a_15667_28111# 0.62fF
C8153 a_12309_38659# a_10873_38517# 1.68fF
C8154 a_11067_27239# _1192_.A2 2.34fF
C8155 pmat.rowoff_n[8] pmat.row_n[9] 3.52fF
C8156 pmat.rowoff_n[12] config_2_in[1] 0.34fF
C8157 a_18546_22542# a_32126_22950# 0.35fF
C8158 a_47278_21540# ctopn 3.58fF
C8159 VDD a_45112_47607# 0.65fF
C8160 a_31214_20536# vcm 0.65fF
C8161 a_29206_65166# a_30210_65166# 0.97fF
C8162 VDD a_46274_22544# 0.52fF
C8163 VDD a_22178_59142# 0.52fF
C8164 a_19166_20536# m2_17932_20266# 0.96fF
C8165 a_12539_10389# a_12705_10389# 0.69fF
C8166 a_36234_21540# a_37238_21540# 0.97fF
C8167 VDD a_18235_35831# 0.63fF
C8168 pmat.sample a_2263_43719# 0.38fF
C8169 a_10441_21263# a_21365_27247# 0.47fF
C8170 VDD a_4535_50639# 0.58fF
C8171 VDD m2_17932_15246# 1.01fF
C8172 a_5899_21807# a_12247_20175# 0.56fF
C8173 ANTENNA__1187__B1.DIODE a_24591_28327# 0.53fF
C8174 ANTENNA__1184__B1.DIODE ANTENNA__1197__B.DIODE 0.87fF
C8175 a_24867_53135# nmat.en_bit_n[1] 1.40fF
C8176 ANTENNA__1190__A1.DIODE _1192_.B1 17.86fF
C8177 a_43262_17524# vcm 0.65fF
C8178 a_40837_46261# a_43720_32143# 0.92fF
C8179 a_2389_45859# a_4257_34319# 0.38fF
C8180 nmat.col_n[31] m2_50060_24282# 0.62fF
C8181 ANTENNA__1395__A1.DIODE a_25695_28111# 0.96fF
C8182 m2_31988_24282# m2_32992_24282# 0.96fF
C8183 a_37238_71190# a_37238_70186# 1.00fF
C8184 a_12309_38659# a_14773_38306# 0.83fF
C8185 a_44266_8488# vcm 0.64fF
C8186 pmat.col_n[13] vcm 2.80fF
C8187 pmat.rowon_n[9] ctopp 1.57fF
C8188 VDD a_19965_43131# 1.15fF
C8189 m2_26968_7214# m2_27972_7214# 0.96fF
C8190 a_7717_14735# a_18563_27791# 0.56fF
C8191 ANTENNA__1190__A1.DIODE a_23395_53135# 0.61fF
C8192 ANTENNA__1190__B1.DIODE _1187_.A2 2.75fF
C8193 a_35244_32411# ANTENNA__1183__B1.DIODE 0.39fF
C8194 a_10239_14183# a_6829_26703# 0.37fF
C8195 a_11067_16359# a_10883_3303# 0.57fF
C8196 clk_ena ctopp 1.19fF
C8197 VDD a_14833_56053# 0.43fF
C8198 VDD a_2419_69455# 7.56fF
C8199 a_11067_30287# a_8583_47381# 0.53fF
C8200 a_35230_13508# a_36234_13508# 0.97fF
C8201 ANTENNA__1183__B1.DIODE nmat.rowon_n[4] 0.87fF
C8202 ANTENNA__1184__B1.DIODE a_31675_47695# 0.32fF
C8203 a_12228_40693# a_11497_40719# 0.36fF
C8204 a_5363_33551# a_6467_29415# 1.36fF
C8205 a_19166_65166# vcm 0.61fF
C8206 cgen.dlycontrol2_in[1] a_11681_35823# 1.94fF
C8207 a_33222_18528# a_34226_18528# 0.97fF
C8208 a_18546_18526# a_49194_18934# 0.35fF
C8209 a_17139_30503# a_44444_32233# 0.77fF
C8210 a_2199_13887# a_3551_6202# 0.38fF
C8211 a_20170_62154# a_20170_61150# 1.00fF
C8212 a_39246_12504# vcm 0.65fF
C8213 a_44266_64162# ctopp 3.58fF
C8214 VDD a_2467_63125# 0.44fF
C8215 VDD a_22178_19532# 0.52fF
C8216 VDD m2_18936_72014# 1.34fF
C8217 a_4081_61127# a_2263_43719# 0.52fF
C8218 a_20170_14512# ctopn 3.57fF
C8219 VDD a_21174_10496# 0.52fF
C8220 VDD a_2847_38975# 0.65fF
C8221 a_34226_20536# ctopn 3.58fF
C8222 a_40250_63158# pmat.col[21] 0.31fF
C8223 a_44266_15516# a_45270_15516# 0.97fF
C8224 a_27498_32117# a_24374_29941# 0.33fF
C8225 VDD a_2195_51701# 0.38fF
C8226 VDD a_18200_27497# 0.46fF
C8227 VDD a_20078_55126# 0.38fF
C8228 a_18546_58180# a_28110_58138# 0.35fF
C8229 a_22178_69182# a_22178_68178# 1.00fF
C8230 a_43262_69182# a_44266_69182# 0.97fF
C8231 a_18546_10494# a_28110_10902# 0.35fF
C8232 _1179_.X ANTENNA__1187__B1.DIODE 1.27fF
C8233 ANTENNA_fanout52_A.DIODE ANTENNA__1197__B.DIODE 4.22fF
C8234 a_30210_21540# a_30210_20536# 1.00fF
C8235 VDD a_7067_34293# 0.47fF
C8236 VDD a_13203_70767# 0.39fF
C8237 a_46274_17524# ctopn 3.58fF
C8238 a_28202_62154# ctopp 3.58fF
C8239 VDD a_37238_62154# 0.52fF
C8240 a_22178_16520# vcm 0.65fF
C8241 a_10873_36341# clk_dig 0.62fF
C8242 a_47278_8488# ctopn 3.40fF
C8243 m2_42028_24282# vcm 0.42fF
C8244 a_18546_56172# a_50198_56130# 0.35fF
C8245 pmat.rowon_n[11] ctopp 1.57fF
C8246 VDD a_49194_24958# 0.45fF
C8247 a_4075_68583# a_5211_57172# 0.74fF
C8248 pmat.rowon_n[5] ctopp 1.57fF
C8249 VDD a_18162_67214# 2.73fF
C8250 VDD a_1949_9308# 0.58fF
C8251 a_11067_64015# a_10515_13967# 0.64fF
C8252 a_47278_65166# ctopp 3.58fF
C8253 _1194_.A2 _1184_.A2 6.96fF
C8254 VDD a_10515_15055# 12.73fF
C8255 a_18546_55168# a_29114_55126# 0.35fF
C8256 nmat.col[24] ANTENNA__1190__A2.DIODE 4.39fF
C8257 pmat.rowoff_n[7] a_18546_63200# 4.09fF
C8258 _1194_.B1 a_10883_3303# 0.66fF
C8259 a_1739_47893# cgen.dlycontrol4_in[4] 3.44fF
C8260 a_27198_70186# ctopp 3.57fF
C8261 a_2007_25597# a_2564_21959# 1.21fF
C8262 VDD a_36234_70186# 0.52fF
C8263 a_23182_15516# ctopn 3.58fF
C8264 a_19166_61150# vcm 0.61fF
C8265 VDD a_23182_11500# 0.52fF
C8266 a_24186_23548# m2_23956_24282# 0.99fF
C8267 nmat.col_n[6] nmat.col[6] 0.71fF
C8268 a_41254_23548# a_41254_22544# 1.00fF
C8269 a_2263_43719# a_18823_50247# 0.34fF
C8270 VDD a_14379_6567# 6.75fF
C8271 a_40250_60146# a_41254_60146# 0.97fF
C8272 a_42258_12504# ctopn 3.58fF
C8273 a_18546_69224# a_23090_69182# 0.35fF
C8274 a_8443_20719# a_12437_28585# 0.40fF
C8275 a_24186_11500# a_24186_10496# 1.00fF
C8276 a_38242_56130# vcm 0.62fF
C8277 pmat.rowoff_n[4] pmat.row_n[3] 2.26fF
C8278 pmat.rowon_n[0] a_1586_18231# 0.48fF
C8279 a_19439_30511# a_19605_30511# 0.39fF
C8280 a_37291_29397# a_37827_30793# 0.68fF
C8281 nmat.en_bit_n[1] pmat.col[9] 0.42fF
C8282 a_18546_63200# a_42166_63158# 0.35fF
C8283 a_48282_68178# a_48282_67174# 1.00fF
C8284 a_26891_28327# a_44444_32233# 1.20fF
C8285 a_29206_61150# a_30210_61150# 0.97fF
C8286 a_41254_66170# vcm 0.62fF
C8287 VDD a_27198_68178# 0.52fF
C8288 pmat.rowoff_n[7] a_2835_13077# 0.69fF
C8289 a_21739_29415# a_43267_47081# 0.34fF
C8290 pmat.col_n[26] pmat.col[26] 0.95fF
C8291 ANTENNA__1190__A1.DIODE a_43720_32143# 0.41fF
C8292 a_19166_11500# m2_17932_11230# 0.96fF
C8293 pmat.row_n[3] nmat.col_n[3] 0.30fF
C8294 a_34226_63158# vcm 0.62fF
C8295 _1194_.A2 a_9411_2215# 0.61fF
C8296 a_33684_32143# a_33869_31599# 0.57fF
C8297 pmat.row_n[15] a_14825_50095# 0.62fF
C8298 VDD a_7803_29673# 0.69fF
C8299 a_6292_65479# a_2879_57487# 0.48fF
C8300 _1196_.B1 _1192_.A2 4.21fF
C8301 VDD a_48190_55126# 0.43fF
C8302 a_4123_76181# a_2149_45717# 0.80fF
C8303 a_4991_69831# a_6927_30503# 0.38fF
C8304 a_36234_24552# m3_36136_24702# 2.45fF
C8305 a_18546_20534# a_29114_20942# 0.35fF
C8306 a_23182_20536# a_24186_20536# 0.97fF
C8307 a_18162_68218# vcm 6.95fF
C8308 a_25190_16520# ctopn 3.58fF
C8309 a_33839_46805# a_33423_47695# 0.42fF
C8310 a_25190_62154# pmat.col[6] 0.31fF
C8311 VDD a_4075_50087# 11.25fF
C8312 a_46274_16520# a_47278_16520# 0.97fF
C8313 a_36234_67174# a_36234_66170# 1.00fF
C8314 a_22178_9492# a_22178_8488# 1.00fF
C8315 pmat.rowon_n[11] a_3746_58487# 1.99fF
C8316 VDD a_32218_23548# 0.55fF
C8317 a_47278_61150# ctopp 3.58fF
C8318 pmat.rowon_n[7] a_12263_50959# 0.53fF
C8319 VDD a_34226_9492# 0.52fF
C8320 a_14773_38306# cgen.dlycontrol1_in[4] 0.41fF
C8321 a_18546_11498# a_32126_11906# 0.35fF
C8322 _1224_.X _1183_.A2 1.95fF
C8323 a_10055_31591# a_9963_13967# 0.33fF
C8324 pmat.en_bit_n[2] a_24407_31375# 0.34fF
C8325 VDD a_30463_41271# 0.61fF
C8326 VDD a_50290_20536# 0.54fF
C8327 VDD a_22269_40391# 1.04fF
C8328 nmat.col[21] m2_40020_24282# 0.41fF
C8329 a_35230_17524# a_36234_17524# 0.97fF
C8330 VDD a_28079_39913# 0.64fF
C8331 pmat.sw ctopp 0.32fF
C8332 a_33222_57134# a_34226_57134# 0.97fF
C8333 ANTENNA__1196__A2.DIODE a_1781_9308# 0.38fF
C8334 a_38242_20536# a_38242_19532# 1.00fF
C8335 a_4075_50087# a_4719_30287# 0.53fF
C8336 pmat.rowoff_n[15] a_1957_43567# 1.68fF
C8337 a_39246_67174# vcm 0.62fF
C8338 a_32218_71190# a_33222_71190# 0.97fF
C8339 a_18546_71232# a_47186_71190# 0.35fF
C8340 VDD cgen.dlycontrol4_in[3] 8.31fF
C8341 a_28202_14512# vcm 0.65fF
C8342 ANTENNA__1197__B.DIODE a_13641_23439# 0.40fF
C8343 a_27198_64162# vcm 0.62fF
C8344 a_36234_8488# a_37238_8488# 0.97fF
C8345 a_4351_55527# a_5784_52423# 1.40fF
C8346 VDD nmat.col[19] 9.84fF
C8347 a_26891_28327# a_32687_46607# 0.61fF
C8348 pmat.col_n[21] ctopp 2.02fF
C8349 a_4167_9615# a_3609_9295# 0.40fF
C8350 a_2972_9991# a_3663_9269# 0.68fF
C8351 a_21371_50087# a_20475_49783# 0.74fF
C8352 a_10883_3303# a_11067_49871# 0.45fF
C8353 VDD a_1770_35015# 0.57fF
C8354 nmat.rowon_n[7] a_2648_29397# 0.61fF
C8355 VDD a_47186_72194# 0.33fF
C8356 VDD a_30210_13508# 0.52fF
C8357 a_44266_14512# a_44266_13508# 1.00fF
C8358 VDD a_19166_62154# 0.56fF
C8359 a_23182_22544# ctopn 3.57fF
C8360 cgen.dlycontrol4_in[4] cgen.dlycontrol4_in[0] 6.63fF
C8361 a_18243_28327# a_25879_31591# 1.63fF
C8362 VDD a_28202_18528# 0.52fF
C8363 m2_38012_54946# vcm 0.42fF
C8364 a_48282_57134# a_48282_56130# 1.00fF
C8365 a_27198_19532# a_27198_18528# 1.00fF
C8366 VDD a_6087_67655# 0.54fF
C8367 a_45270_62154# pmat.col[26] 0.31fF
C8368 VDD a_39246_15516# 0.52fF
C8369 a_18546_14510# a_30118_14918# 0.35fF
C8370 a_24374_29941# a_13641_23439# 1.05fF
C8371 pmat.row_n[14] a_18162_22544# 25.57fF
C8372 a_18546_64204# a_28110_64162# 0.35fF
C8373 a_3267_74817# a_3228_74691# 0.72fF
C8374 a_6200_70919# a_3339_70759# 0.89fF
C8375 a_20170_59142# a_20170_58138# 1.00fF
C8376 a_2411_16101# a_1591_15829# 0.34fF
C8377 VDD a_18546_70228# 32.63fF
C8378 _1179_.X a_5179_31591# 1.01fF
C8379 pmat.row_n[9] ctopn 1.65fF
C8380 a_18546_72236# a_24094_72194# 0.35fF
C8381 a_14287_69455# pmat.row_n[6] 1.52fF
C8382 VDD m2_45040_7214# 0.91fF
C8383 a_6283_31591# a_26479_32117# 2.14fF
C8384 a_17902_43439# a_11021_43011# 1.10fF
C8385 a_2149_45717# a_5779_71285# 0.61fF
C8386 VDD a_7111_74575# 0.49fF
C8387 a_30210_65166# vcm 0.62fF
C8388 ANTENNA__1195__A1.DIODE a_34942_51701# 0.58fF
C8389 pmat.row_n[7] a_18162_15516# 25.57fF
C8390 a_37238_21540# vcm 0.65fF
C8391 a_26194_60146# ctopp 3.58fF
C8392 VDD a_35230_60146# 0.52fF
C8393 ANTENNA__1190__A1.DIODE a_30663_50087# 0.45fF
C8394 a_18546_21538# a_19074_21946# 0.35fF
C8395 VDD a_2944_72104# 0.54fF
C8396 cgen.start_conv_in clk_ena 1.30fF
C8397 nmat.col_n[3] a_10839_11989# 0.37fF
C8398 a_25190_17524# a_25190_16520# 1.00fF
C8399 nmat.col_n[28] nmat.col_n[30] 0.69fF
C8400 a_18546_19530# a_41162_19938# 0.35fF
C8401 m2_27972_54946# m2_28976_54946# 0.96fF
C8402 a_19166_71190# a_19166_70186# 1.00fF
C8403 a_12447_16143# a_7779_22583# 0.59fF
C8404 a_31214_14512# ctopn 3.58fF
C8405 _1179_.X a_25575_31055# 0.40fF
C8406 ANTENNA__1395__B1.DIODE a_22628_30485# 0.36fF
C8407 a_31214_12504# a_32218_12504# 0.97fF
C8408 a_18546_12502# a_45178_12910# 0.35fF
C8409 VDD a_29159_37607# 1.54fF
C8410 ANTENNA_fanout52_A.DIODE a_32162_34191# 0.59fF
C8411 a_6568_59887# a_5731_58951# 0.64fF
C8412 a_44266_22544# a_45270_22544# 0.97fF
C8413 VDD a_41254_16520# 0.52fF
C8414 a_18546_59184# a_23090_59142# 0.35fF
C8415 a_20170_59142# a_21174_59142# 0.97fF
C8416 VDD a_31122_55126# 0.42fF
C8417 ANTENNA__1187__B1.DIODE nmat.col[7] 0.63fF
C8418 VDD a_51202_7890# 0.40fF
C8419 _1224_.X ANTENNA__1395__A1.DIODE 2.12fF
C8420 pmat.rowon_n[0] cgen.dlycontrol2_in[0] 0.47fF
C8421 VDD a_28202_57134# 0.52fF
C8422 VDD a_1591_33775# 0.38fF
C8423 a_44266_69182# vcm 0.62fF
C8424 VDD a_27198_71190# 0.55fF
C8425 a_28629_48437# a_29076_48695# 0.39fF
C8426 a_4075_31591# a_2046_30184# 0.44fF
C8427 a_18546_23546# a_50198_23954# 0.35fF
C8428 a_10781_42869# a_13503_43421# 0.32fF
C8429 a_3367_14906# a_3063_14741# 0.36fF
C8430 a_27198_71190# m2_26968_72014# 1.00fF
C8431 VDD a_33467_46261# 4.29fF
C8432 VDD a_5899_21807# 3.53fF
C8433 VDD ANTENNA__1184__B1.DIODE 24.75fF
C8434 pmat.row_n[13] a_18162_69222# 25.57fF
C8435 VDD a_10047_8751# 1.03fF
C8436 VDD a_33765_40229# 1.34fF
C8437 VDD a_17021_38053# 1.22fF
C8438 a_18162_71230# vcm 6.95fF
C8439 VDD a_26331_42089# 0.62fF
C8440 VDD a_10515_61839# 23.70fF
C8441 a_18546_55168# a_39154_55126# 0.35fF
C8442 pmat.sample_n cgen.dlycontrol4_in[3] 0.35fF
C8443 a_18546_24550# a_28110_24958# 0.35fF
C8444 nmat.col[29] nmat.col[26] 2.63fF
C8445 _1187_.A2 nmat.col_n[21] 4.75fF
C8446 pmat.row_n[1] a_18162_57174# 25.57fF
C8447 a_48282_56130# ctopp 3.40fF
C8448 a_18243_28327# nmat.col_n[9] 0.32fF
C8449 a_30210_61150# vcm 0.62fF
C8450 a_10515_13967# a_3571_13627# 0.30fF
C8451 nmat.rowon_n[14] a_2835_13077# 0.76fF
C8452 a_6787_47607# a_6927_30503# 0.40fF
C8453 pmat.row_n[10] pmat.row_n[9] 15.62fF
C8454 a_18546_22542# a_25098_22950# 0.35fF
C8455 a_40250_21540# ctopn 3.58fF
C8456 a_10873_39605# a_21981_34191# 0.93fF
C8457 VDD m2_51064_55950# 1.06fF
C8458 pmat.rowoff_n[4] ANTENNA__1195__A1.DIODE 0.35fF
C8459 a_24186_20536# vcm 0.65fF
C8460 a_21739_29415# a_28131_50069# 1.40fF
C8461 VDD a_39246_22544# 0.52fF
C8462 VDD a_27498_32117# 0.65fF
C8463 a_1923_61759# a_2163_61761# 0.32fF
C8464 VDD a_6823_58951# 0.56fF
C8465 nmat.col[22] ctopn 1.97fF
C8466 VDD a_11297_36091# 6.06fF
C8467 pmat.rowon_n[8] pmat.rowoff_n[4] 0.70fF
C8468 VDD pmat.col_n[14] 5.21fF
C8469 a_44266_63158# ctopp 3.58fF
C8470 nmat.rowoff_n[11] nmat.rowoff_n[5] 0.38fF
C8471 a_12311_54135# a_12003_52815# 0.32fF
C8472 a_36234_17524# vcm 0.65fF
C8473 m2_49056_24282# m3_49188_24414# 2.79fF
C8474 m2_18936_55950# vcm 0.44fF
C8475 VDD a_13151_23957# 0.51fF
C8476 m2_24960_24282# m2_25964_24282# 0.96fF
C8477 a_37238_8488# vcm 0.64fF
C8478 nmat.col_n[14] nmat.col[14] 0.71fF
C8479 m2_19940_7214# m2_20944_7214# 0.96fF
C8480 a_5363_70543# a_13462_48071# 0.47fF
C8481 a_47278_18528# a_47278_17524# 1.00fF
C8482 a_16311_28327# a_15667_27239# 4.37fF
C8483 a_10239_14183# a_12079_9615# 0.83fF
C8484 VDD a_19439_30511# 0.41fF
C8485 m2_51064_60970# m2_51064_59966# 0.99fF
C8486 a_18546_13506# a_46182_13914# 0.35fF
C8487 a_6283_31591# a_5179_31591# 2.34fF
C8488 VDD ANTENNA_fanout52_A.DIODE 15.74fF
C8489 _1194_.B1 a_7717_14735# 0.61fF
C8490 a_47278_63158# a_47278_62154# 1.00fF
C8491 a_46274_71190# m2_46044_72014# 1.00fF
C8492 a_19166_21540# vcm 0.65fF
C8493 _1224_.X ANTENNA__1395__A2.DIODE 1.03fF
C8494 a_49286_67174# ctopp 3.57fF
C8495 a_16800_47213# a_6283_31591# 0.55fF
C8496 a_25879_31591# a_11948_49783# 1.36fF
C8497 a_18546_18526# a_42166_18934# 0.35fF
C8498 a_23182_70186# a_23182_69182# 1.00fF
C8499 a_11317_36924# a_12345_36924# 0.32fF
C8500 VDD a_30371_37737# 0.58fF
C8501 a_2411_16101# a_1591_18005# 0.33fF
C8502 nmat.rowon_n[12] comp_latch 2.06fF
C8503 a_32218_12504# vcm 0.65fF
C8504 a_37238_64162# ctopp 3.58fF
C8505 nmat.col_n[12] a_10814_29111# 0.34fF
C8506 VDD a_47278_14512# 0.52fF
C8507 _1194_.A2 nmat.col[24] 0.40fF
C8508 m2_41024_7214# m3_41156_7346# 2.79fF
C8509 VDD a_46274_64162# 0.52fF
C8510 a_17842_27497# a_28336_29967# 0.34fF
C8511 VDD a_19166_58138# 0.56fF
C8512 nmat.rowon_n[5] nmat.col[7] 0.37fF
C8513 a_5566_44905# a_4955_40277# 0.47fF
C8514 pmat.row_n[3] vcm 1.21fF
C8515 VDD a_4167_9615# 0.30fF
C8516 VDD a_47211_50069# 0.44fF
C8517 a_46274_13508# a_46274_12504# 1.00fF
C8518 a_27198_20536# ctopn 3.58fF
C8519 nmat.rowoff_n[14] a_18546_9490# 4.09fF
C8520 VDD a_35068_46805# 0.49fF
C8521 a_17842_27497# nmat.col[3] 1.67fF
C8522 VDD pmat.col[13] 5.17fF
C8523 a_41731_49525# nmat.col[21] 0.63fF
C8524 VDD a_6634_26133# 0.59fF
C8525 a_18546_58180# a_21082_58138# 0.35fF
C8526 ANTENNA__1195__A1.DIODE a_41731_49525# 3.15fF
C8527 VDD a_3431_57167# 0.35fF
C8528 _1192_.A2 a_45019_38645# 0.49fF
C8529 VDD a_22743_35561# 0.65fF
C8530 ANTENNA__1197__B.DIODE a_13091_28327# 1.00fF
C8531 a_39246_17524# ctopn 3.58fF
C8532 a_21174_62154# ctopp 3.58fF
C8533 VDD a_30210_62154# 0.52fF
C8534 a_40250_8488# ctopn 3.40fF
C8535 VDD a_21147_49525# 0.36fF
C8536 a_18546_56172# a_43170_56130# 0.35fF
C8537 a_30210_56130# a_31214_56130# 0.97fF
C8538 VDD a_42166_24958# 0.44fF
C8539 nmat.col[31] nmat.col_n[31] 1.41fF
C8540 a_21739_29415# nmat.col_n[31] 0.32fF
C8541 a_10055_31591# a_2935_38279# 1.72fF
C8542 a_40250_65166# ctopp 3.58fF
C8543 nmat.col[29] clk_ena 0.58fF
C8544 VDD a_49286_65166# 0.52fF
C8545 a_18546_55168# a_22086_55126# 0.35fF
C8546 a_18546_24550# a_18162_24552# 2.54fF
C8547 nmat.col_n[1] a_20170_24552# 0.31fF
C8548 VDD a_6821_18543# 1.39fF
C8549 ANTENNA__1395__B1.DIODE nmat.col_n[13] 1.96fF
C8550 a_18546_68220# a_51202_68178# 0.35fF
C8551 VDD a_25681_28879# 0.89fF
C8552 a_20170_70186# ctopp 3.56fF
C8553 a_20170_20536# a_20170_19532# 1.00fF
C8554 VDD a_29206_70186# 0.52fF
C8555 a_6283_31591# a_5935_46983# 0.40fF
C8556 nmat.sw a_11067_30287# 0.56fF
C8557 VDD a_2847_26133# 0.35fF
C8558 _1224_.X ANTENNA__1196__A2.DIODE 4.16fF
C8559 a_3339_70759# a_5784_52423# 1.56fF
C8560 a_35230_62154# a_36234_62154# 0.97fF
C8561 a_42258_16520# a_42258_15516# 1.00fF
C8562 VDD m2_17932_56954# 1.00fF
C8563 VDD a_5566_44905# 1.11fF
C8564 a_33222_66170# a_34226_66170# 0.97fF
C8565 a_1781_9308# a_4379_13818# 0.32fF
C8566 a_5535_57993# a_5528_57685# 0.54fF
C8567 a_9135_60967# a_9577_58229# 0.58fF
C8568 a_10883_3303# nmat.col_n[0] 3.78fF
C8569 m2_32992_72014# m3_33124_72146# 2.79fF
C8570 a_35230_12504# ctopn 3.58fF
C8571 a_16966_29673# nmat.col_n[3] 0.42fF
C8572 a_31214_56130# vcm 0.62fF
C8573 VDD a_12311_54135# 0.39fF
C8574 pmat.rowoff_n[7] a_1858_25615# 2.59fF
C8575 nmat.col[10] ANTENNA__1183__B1.DIODE 2.01fF
C8576 a_12345_39100# a_11681_35823# 1.07fF
C8577 a_26194_63158# a_27198_63158# 0.97fF
C8578 a_18546_63200# a_35138_63158# 0.35fF
C8579 ANTENNA__1197__A.DIODE a_41949_30761# 0.73fF
C8580 a_2411_43301# pmat.rowon_n[0] 0.36fF
C8581 a_25695_28111# a_2007_25597# 0.53fF
C8582 a_34226_66170# vcm 0.62fF
C8583 VDD a_20170_68178# 0.52fF
C8584 m2_44036_72014# m2_45040_72014# 0.96fF
C8585 a_1781_9308# a_2007_25597# 0.62fF
C8586 a_4719_30287# a_5566_44905# 0.33fF
C8587 a_27198_63158# vcm 0.62fF
C8588 VDD a_4339_27804# 3.99fF
C8589 _1179_.X a_18243_28327# 0.66fF
C8590 cgen.dlycontrol2_in[4] a_13909_39605# 2.32fF
C8591 VDD a_41162_55126# 0.42fF
C8592 VDD a_13641_23439# 5.15fF
C8593 VDD dummypin[14] 1.05fF
C8594 VDD pmat.col[23] 4.91fF
C8595 a_18546_20534# a_22086_20942# 0.35fF
C8596 ANTENNA__1197__B.DIODE a_17139_30503# 0.51fF
C8597 nmat.en_bit_n[1] a_13643_29415# 6.01fF
C8598 pmat.rowoff_n[12] nmat.rowon_n[14] 1.80fF
C8599 pmat.row_n[6] a_17139_30503# 0.33fF
C8600 a_5651_66975# a_1957_43567# 0.52fF
C8601 a_11435_58791# a_3746_58487# 0.82fF
C8602 VDD a_25190_23548# 0.55fF
C8603 pmat.col_n[9] pmat.col[9] 0.75fF
C8604 a_40250_61150# ctopp 3.58fF
C8605 a_34226_70186# a_35230_70186# 0.97fF
C8606 VDD a_27198_9492# 0.52fF
C8607 pmat.row_n[1] vcm 1.18fF
C8608 VDD a_49286_61150# 0.52fF
C8609 a_21174_11500# a_22178_11500# 0.97fF
C8610 a_18546_11498# a_25098_11906# 0.35fF
C8611 pmat.rowon_n[7] a_12447_16143# 1.54fF
C8612 a_19166_64162# ctopp 3.43fF
C8613 _1187_.A2 nmat.col_n[10] 0.39fF
C8614 a_15667_27239# pmat.col[26] 0.47fF
C8615 a_36234_24552# ctopn 0.65fF
C8616 VDD a_43262_20536# 0.52fF
C8617 a_23182_64162# a_23182_63158# 1.00fF
C8618 m2_51064_63982# vcm 0.51fF
C8619 pmat.col_n[0] pmat.col[1] 5.99fF
C8620 a_26194_10496# a_26194_9492# 1.00fF
C8621 _1187_.A2 clk_ena 0.32fF
C8622 a_17139_30503# a_31675_47695# 0.46fF
C8623 ANTENNA__1395__A1.DIODE nmat.col[28] 0.58fF
C8624 a_32218_67174# vcm 0.62fF
C8625 a_1923_69823# a_2163_74173# 0.56fF
C8626 a_2727_58470# a_1923_61759# 1.11fF
C8627 a_18546_71232# a_40158_71190# 0.35fF
C8628 a_18546_9490# vcm 0.40fF
C8629 VDD a_14287_69455# 3.26fF
C8630 a_14887_46377# a_1781_9308# 1.93fF
C8631 a_23182_58138# a_23182_57134# 1.00fF
C8632 a_21174_14512# vcm 0.65fF
C8633 a_24833_40719# a_10873_40693# 0.35fF
C8634 VDD a_10223_26703# 2.37fF
C8635 a_20170_64162# vcm 0.62fF
C8636 a_11067_30287# a_1858_25615# 1.75fF
C8637 a_18546_8486# a_48190_8894# 0.35fF
C8638 a_27198_60146# a_27198_59142# 1.00fF
C8639 a_18546_65208# a_45178_65166# 0.35fF
C8640 VDD a_26583_34343# 1.11fF
C8641 a_45270_62154# a_45270_61150# 1.00fF
C8642 VDD a_23182_13508# 0.52fF
C8643 cgen.dlycontrol3_in[0] a_10873_39605# 3.12fF
C8644 VDD a_21174_18528# 0.52fF
C8645 a_19166_16520# a_20170_16520# 0.97fF
C8646 a_18546_67216# a_45178_67174# 0.35fF
C8647 a_31214_67174# a_32218_67174# 0.97fF
C8648 a_7026_24527# a_6173_22895# 0.32fF
C8649 a_4128_64391# a_14379_6567# 1.21fF
C8650 pmat.rowoff_n[14] pmat.rowon_n[14] 20.86fF
C8651 a_17139_30503# a_19605_30511# 0.60fF
C8652 pmat.row_n[8] nmat.rowoff_n[6] 0.52fF
C8653 a_28202_66170# a_28202_65166# 1.00fF
C8654 a_21174_22544# a_21174_21540# 1.00fF
C8655 pmat.col_n[16] vcm 2.79fF
C8656 nmat.rowoff_n[6] a_12437_28879# 1.69fF
C8657 VDD a_30913_43131# 1.41fF
C8658 VDD a_32218_15516# 0.52fF
C8659 nmat.col_n[4] nmat.col[5] 6.69fF
C8660 nmat.col[23] nmat.col_n[22] 6.78fF
C8661 a_6787_47607# a_10864_68565# 0.46fF
C8662 a_45270_15516# a_45270_14512# 1.00fF
C8663 a_18546_14510# a_23090_14918# 0.35fF
C8664 pmat.col[19] vcm 5.88fF
C8665 _1154_.A ANTENNA__1197__A.DIODE 0.68fF
C8666 a_18546_7482# a_45178_7890# 0.35fF
C8667 a_18546_64204# a_21082_64162# 0.35fF
C8668 a_25190_68178# a_26194_68178# 0.97fF
C8669 a_47278_69182# a_47278_68178# 1.00fF
C8670 a_2835_13077# a_3571_13627# 1.44fF
C8671 VDD a_9139_68841# 0.79fF
C8672 a_1957_43567# cgen.dlycontrol3_in[4] 1.28fF
C8673 VDD nmat.col_n[29] 9.14fF
C8674 VDD m2_30984_7214# 1.28fF
C8675 a_2263_43719# a_26155_46831# 0.57fF
C8676 a_1586_33927# a_6007_42479# 0.34fF
C8677 VDD a_7092_74005# 1.09fF
C8678 a_3571_13627# a_4075_13653# 0.31fF
C8679 a_23182_65166# vcm 0.62fF
C8680 a_30210_21540# vcm 0.65fF
C8681 VDD a_3859_22655# 0.34fF
C8682 a_7644_16341# a_9485_15279# 0.53fF
C8683 VDD a_28202_60146# 0.52fF
C8684 a_11067_64015# nmat.sw 0.96fF
C8685 pmat.sw nmat.col[29] 0.63fF
C8686 a_50290_10496# m2_51064_10226# 0.96fF
C8687 a_45270_58138# vcm 0.62fF
C8688 nmat.col[21] vcm 8.60fF
C8689 a_47278_56130# m2_47048_54946# 0.99fF
C8690 VDD pmat.rowoff_n[10] 2.02fF
C8691 a_4396_66933# a_4298_67191# 0.89fF
C8692 a_9405_66627# a_9643_66389# 0.37fF
C8693 nmat.rowon_n[5] nmat.rowoff_n[5] 20.33fF
C8694 _1179_.X a_18547_51565# 0.36fF
C8695 a_18243_28327# pmat.col[0] 0.40fF
C8696 a_18546_19530# a_34134_19938# 0.35fF
C8697 m2_20944_54946# m2_21948_54946# 0.96fF
C8698 pmat.rowon_n[8] vcm 0.88fF
C8699 a_24186_14512# ctopn 3.58fF
C8700 a_13091_28327# a_22459_28879# 0.44fF
C8701 a_13459_28111# a_13479_26935# 1.13fF
C8702 a_18546_12502# a_38150_12910# 0.35fF
C8703 VDD a_13443_39095# 0.60fF
C8704 VDD a_11149_40188# 6.78fF
C8705 a_1957_43567# a_11547_48061# 0.36fF
C8706 VDD a_34226_16520# 0.52fF
C8707 VDD a_6817_51733# 0.65fF
C8708 a_21174_65166# a_21174_64162# 1.00fF
C8709 a_26891_28327# a_31675_47695# 1.59fF
C8710 VDD a_24094_55126# 0.42fF
C8711 VDD a_4951_31029# 0.47fF
C8712 _1183_.A2 ANTENNA__1183__B1.DIODE 8.64fF
C8713 VDD a_44174_7890# 0.33fF
C8714 VDD a_4720_58487# 0.32fF
C8715 a_49286_11500# a_49286_10496# 1.00fF
C8716 m3_36136_24702# ctopn 0.36fF
C8717 VDD a_21174_57134# 0.52fF
C8718 _1194_.B1 ANTENNA__1195__A1.DIODE 0.86fF
C8719 ANTENNA__1197__B.DIODE _1184_.A2 1.30fF
C8720 a_11067_27239# a_16311_28327# 2.81fF
C8721 a_37238_69182# vcm 0.62fF
C8722 VDD a_20170_71190# 0.56fF
C8723 _1184_.A2 a_10378_7637# 0.84fF
C8724 a_30210_23548# a_31214_23548# 0.97fF
C8725 a_18546_23546# a_43170_23954# 0.35fF
C8726 a_4523_21276# a_5899_21807# 0.59fF
C8727 m2_51064_17254# m2_51064_16250# 0.99fF
C8728 a_32218_9492# a_33222_9492# 0.97fF
C8729 a_18546_9490# a_47186_9898# 0.35fF
C8730 pmat.row_n[1] a_11067_49871# 0.48fF
C8731 a_1781_9308# a_7109_29423# 5.77fF
C8732 a_46274_59142# vcm 0.62fF
C8733 a_10239_14183# a_4703_24527# 0.92fF
C8734 VDD a_15093_39638# 1.15fF
C8735 a_39246_12504# a_39246_11500# 1.00fF
C8736 a_12658_42895# a_11297_36091# 2.21fF
C8737 VDD a_11921_41814# 2.12fF
C8738 VDD a_2400_13763# 0.40fF
C8739 VDD a_5065_63669# 0.35fF
C8740 nmat.rowon_n[14] a_1858_25615# 1.98fF
C8741 a_41254_56130# ctopp 3.40fF
C8742 _1184_.A2 a_31675_47695# 0.71fF
C8743 VDD a_50290_56130# 0.59fF
C8744 a_48282_20536# a_49286_20536# 0.97fF
C8745 a_36234_8488# m2_36004_7214# 1.00fF
C8746 a_23182_61150# vcm 0.62fF
C8747 pmat.row_n[5] nmat.sample 0.35fF
C8748 pmat.row_n[7] a_11067_16359# 0.36fF
C8749 a_33222_21540# ctopn 3.58fF
C8750 ANTENNA__1184__B1.DIODE a_8583_29199# 1.69fF
C8751 a_45119_32661# a_45277_32687# 0.34fF
C8752 ANTENNA__1395__B1.DIODE a_28915_50959# 1.43fF
C8753 a_47278_9492# a_47278_8488# 1.00fF
C8754 a_22178_65166# a_23182_65166# 0.97fF
C8755 a_44266_66170# ctopp 3.58fF
C8756 VDD a_32218_22544# 0.52fF
C8757 VDD a_20695_32447# 0.33fF
C8758 pmat.col_n[1] ctopp 2.01fF
C8759 nmat.col[11] ctopn 1.97fF
C8760 a_29206_21540# a_30210_21540# 0.97fF
C8761 a_37238_63158# ctopp 3.58fF
C8762 VDD a_46274_63158# 0.52fF
C8763 a_29206_17524# vcm 0.65fF
C8764 cgen.dlycontrol4_in[4] cgen.dlycontrol4_in[3] 0.99fF
C8765 pmat.rowon_n[0] pmat.rowoff_n[0] 20.79fF
C8766 pmat.row_n[12] pmat.rowoff_n[2] 1.09fF
C8767 a_2389_45859# a_4313_44111# 0.42fF
C8768 a_18546_61192# a_45178_61150# 0.35fF
C8769 a_30210_71190# a_30210_70186# 1.00fF
C8770 a_30210_8488# vcm 0.64fF
C8771 a_14691_27399# a_11927_27399# 0.49fF
C8772 a_44266_58138# a_45270_58138# 0.97fF
C8773 pmat.row_n[9] ctopp 1.65fF
C8774 VDD a_30543_40721# 1.93fF
C8775 pmat.row_n[14] ANTENNA__1196__A2.DIODE 0.99fF
C8776 a_12116_40871# a_21981_34191# 1.69fF
C8777 a_1923_53055# a_2715_51969# 0.96fF
C8778 VDD m2_51064_20266# 1.04fF
C8779 a_26479_32117# nmat.col_n[12] 0.35fF
C8780 a_46274_19532# vcm 0.65fF
C8781 a_6927_30503# a_12613_57141# 0.36fF
C8782 a_19166_10496# ctopn 3.43fF
C8783 VDD comp.adc_nor_latch_0.R 1.01fF
C8784 a_45270_10496# vcm 0.65fF
C8785 a_28202_13508# a_29206_13508# 0.97fF
C8786 a_18546_13506# a_39154_13914# 0.35fF
C8787 VDD a_13327_70741# 2.22fF
C8788 VDD a_13091_28327# 13.35fF
C8789 VDD a_2861_76757# 0.67fF
C8790 pmat.row_n[7] vcm 1.18fF
C8791 _1154_.X nmat.col[21] 0.36fF
C8792 a_44266_61150# a_44266_60146# 1.00fF
C8793 a_42258_67174# ctopp 3.58fF
C8794 a_6559_33767# a_9827_53379# 0.47fF
C8795 _1154_.X ANTENNA__1195__A1.DIODE 6.35fF
C8796 a_26194_18528# a_27198_18528# 0.97fF
C8797 a_18546_18526# a_35138_18934# 0.35fF
C8798 VDD a_12237_60431# 0.38fF
C8799 nmat.col_n[13] nmat.col[18] 1.86fF
C8800 a_25190_12504# vcm 0.65fF
C8801 a_30210_64162# ctopp 3.58fF
C8802 a_21739_29415# nmat.col[10] 0.39fF
C8803 VDD a_40250_14512# 0.52fF
C8804 VDD a_39246_64162# 0.52fF
C8805 pmat.en_bit_n[0] a_15101_29423# 0.57fF
C8806 VDD a_28975_40871# 0.42fF
C8807 nmat.col[28] m2_47048_24282# 0.39fF
C8808 VDD a_36227_38771# 1.43fF
C8809 pmat.rowon_n[13] ctopp 1.57fF
C8810 a_45270_59142# a_45270_58138# 1.00fF
C8811 a_38851_28327# a_35244_32411# 1.45fF
C8812 a_18547_51565# a_6283_31591# 0.57fF
C8813 a_12263_50959# a_13275_48783# 2.87fF
C8814 VDD a_7373_49007# 0.89fF
C8815 a_46274_23548# m2_46044_24282# 0.99fF
C8816 pmat.rowoff_n[7] config_2_in[9] 0.42fF
C8817 VDD config_1_in[8] 1.02fF
C8818 _1194_.B1 a_7415_29397# 0.93fF
C8819 a_37238_15516# a_38242_15516# 0.97fF
C8820 VDD m2_28976_24282# 0.62fF
C8821 pmat.rowoff_n[7] a_18162_15516# 1.33fF
C8822 a_36234_69182# a_37238_69182# 0.97fF
C8823 a_4583_68021# a_3923_68021# 0.47fF
C8824 VDD a_27155_31599# 1.96fF
C8825 VDD pmat.rowoff_n[3] 2.69fF
C8826 a_3615_71631# a_5363_33551# 1.56fF
C8827 pmat.col_n[24] ctopp 2.02fF
C8828 a_1586_18231# a_4976_16091# 0.43fF
C8829 pmat.row_n[15] a_2046_30184# 0.97fF
C8830 a_23182_21540# a_23182_20536# 1.00fF
C8831 a_19166_69182# vcm 0.61fF
C8832 a_5351_19913# a_9528_20407# 0.43fF
C8833 a_32218_17524# ctopn 3.58fF
C8834 VDD a_50198_72194# 0.32fF
C8835 a_47278_11500# vcm 0.65fF
C8836 pmat.col[21] vcm 5.88fF
C8837 VDD a_23182_62154# 0.52fF
C8838 a_28336_29967# a_28715_28879# 0.35fF
C8839 a_50290_17524# a_50290_16520# 1.00fF
C8840 a_33222_8488# ctopn 3.40fF
C8841 a_1591_31599# config_2_in[10] 0.73fF
C8842 a_18546_56172# a_36142_56130# 0.35fF
C8843 VDD a_35138_24958# 0.39fF
C8844 a_4719_30287# a_7373_49007# 0.76fF
C8845 m2_48052_24282# m2_49056_24282# 0.96fF
C8846 VDD a_1644_60949# 0.33fF
C8847 a_49286_19532# ctopn 3.57fF
C8848 a_33222_65166# ctopp 3.58fF
C8849 a_4523_21276# a_6821_18543# 1.37fF
C8850 VDD a_42258_65166# 0.52fF
C8851 VDD a_49286_21540# 0.52fF
C8852 a_45270_59142# a_46274_59142# 0.97fF
C8853 a_1858_25615# a_15435_29111# 0.31fF
C8854 m2_17932_66994# vcm 0.44fF
C8855 a_48282_10496# ctopn 3.58fF
C8856 a_18546_68220# a_44174_68178# 0.35fF
C8857 a_2149_45717# a_2407_49289# 1.17fF
C8858 a_2419_53351# a_5497_62839# 0.36fF
C8859 VDD a_22178_70186# 0.52fF
C8860 a_18546_72236# a_27106_72194# 0.35fF
C8861 VDD a_13145_26935# 0.99fF
C8862 a_34226_23548# a_34226_22544# 1.00fF
C8863 _1192_.B1 nmat.col_n[4] 0.40fF
C8864 _1224_.X pmat.col[25] 0.39fF
C8865 VDD nmat.rowon_n[6] 3.46fF
C8866 a_11435_58791# a_9427_50095# 0.41fF
C8867 VDD a_17139_30503# 16.71fF
C8868 nmat.rowoff_n[11] nmat.rowoff_n[10] 0.85fF
C8869 _1196_.B1 a_16311_28327# 0.70fF
C8870 VDD a_36178_48169# 0.45fF
C8871 a_12907_54997# a_13073_54997# 0.69fF
C8872 a_18546_60188# a_49194_60146# 0.35fF
C8873 a_33222_60146# a_34226_60146# 0.97fF
C8874 cgen.dlycontrol3_in[0] cgen.dlycontrol2_in[2] 0.86fF
C8875 a_28202_12504# ctopn 3.58fF
C8876 a_2952_25045# a_4068_25615# 0.66fF
C8877 a_11317_36924# a_10873_36341# 1.53fF
C8878 a_24186_56130# vcm 0.62fF
C8879 a_20170_21540# a_21174_21540# 0.97fF
C8880 VDD a_28061_36965# 1.36fF
C8881 VDD a_11115_71285# 1.74fF
C8882 a_19166_63158# ctopp 3.43fF
C8883 a_18546_63200# a_28110_63158# 0.35fF
C8884 VDD m2_48052_72014# 1.10fF
C8885 a_41254_68178# a_41254_67174# 1.00fF
C8886 cgen.dlycontrol3_in[4] a_12228_39605# 0.52fF
C8887 a_22178_61150# a_23182_61150# 0.97fF
C8888 a_47278_69182# ctopp 3.58fF
C8889 a_24407_31375# a_15667_27239# 5.45fF
C8890 pmat.row_n[13] nmat.sample 0.35fF
C8891 a_27198_66170# vcm 0.62fF
C8892 m2_37008_72014# m2_38012_72014# 0.96fF
C8893 nmat.rowon_n[7] pmat.row_n[4] 0.41fF
C8894 cgen.enable_dlycontrol_in nmat.sample 0.45fF
C8895 VDD a_1757_43029# 0.62fF
C8896 a_20170_63158# vcm 0.62fF
C8897 VDD a_40741_46565# 0.52fF
C8898 a_37471_32149# a_37637_32149# 0.46fF
C8899 a_13275_48783# clk_ena 0.51fF
C8900 nmat.sw cgen.dlycontrol1_in[1] 4.96fF
C8901 VDD a_34226_55126# 0.59fF
C8902 a_50290_11500# ctopn 3.43fF
C8903 _1224_.X ANTENNA__1190__B1.DIODE 1.17fF
C8904 pmat.col_n[7] a_23395_53135# 0.46fF
C8905 a_33467_46261# a_41663_47893# 0.32fF
C8906 a_18546_13506# a_21082_13914# 0.35fF
C8907 VDD a_5403_67655# 2.01fF
C8908 inp_analog _1192_.B1 0.37fF
C8909 a_5899_21807# a_3305_15823# 1.03fF
C8910 a_11337_25071# a_14371_25071# 0.78fF
C8911 a_39246_16520# a_40250_16520# 0.97fF
C8912 a_25879_31591# a_32687_46607# 0.98fF
C8913 a_29206_67174# a_29206_66170# 1.00fF
C8914 VDD a_45164_40847# 0.45fF
C8915 a_22153_37179# a_11317_36924# 1.94fF
C8916 VDD a_23700_38567# 1.18fF
C8917 a_33222_61150# ctopp 3.58fF
C8918 VDD a_42258_61150# 0.52fF
C8919 a_27603_34191# a_27687_34967# 0.70fF
C8920 VDD a_36617_42043# 1.42fF
C8921 a_1957_43567# a_14491_51969# 0.33fF
C8922 a_11435_58791# a_4383_7093# 0.37fF
C8923 a_29635_31029# a_29455_31293# 0.32fF
C8924 a_8583_29199# a_13641_23439# 1.05fF
C8925 VDD a_36234_20536# 0.52fF
C8926 VDD a_3295_40277# 0.33fF
C8927 a_28202_17524# a_29206_17524# 0.97fF
C8928 a_26194_57134# a_27198_57134# 0.97fF
C8929 a_14773_39394# a_23700_38567# 0.38fF
C8930 a_31214_20536# a_31214_19532# 1.00fF
C8931 pmat.sample_n pmat.rowoff_n[3] 0.42fF
C8932 a_25190_67174# vcm 0.62fF
C8933 a_18546_71232# a_33130_71190# 0.35fF
C8934 a_25190_71190# a_26194_71190# 0.97fF
C8935 a_11067_30287# a_26321_46831# 0.60fF
C8936 a_19166_59142# m2_17932_58962# 0.96fF
C8937 VDD a_48282_17524# 0.52fF
C8938 a_11113_39747# a_12116_39783# 2.20fF
C8939 a_11149_40188# a_11113_40835# 0.32fF
C8940 a_7717_14735# a_8507_20175# 0.58fF
C8941 VDD a_11927_27399# 4.70fF
C8942 _1194_.B1 a_9307_31068# 1.29fF
C8943 VDD m2_24960_54946# 0.62fF
C8944 VDD a_39647_47679# 0.49fF
C8945 a_21739_29415# _1183_.A2 0.88fF
C8946 a_18546_8486# a_41162_8894# 0.35fF
C8947 a_29206_8488# a_30210_8488# 0.97fF
C8948 a_1923_69823# a_2163_71997# 0.49fF
C8949 VDD a_7658_71543# 4.75fF
C8950 a_18546_65208# a_38150_65166# 0.35fF
C8951 pmat.row_n[11] nmat.sample 0.34fF
C8952 a_48282_70186# a_48282_69182# 1.00fF
C8953 VDD a_32957_30287# 0.60fF
C8954 VDD a_49286_8488# 0.55fF
C8955 VDD a_18162_59182# 2.73fF
C8956 nmat.col[9] vcm 5.76fF
C8957 pmat.row_n[12] a_19283_49783# 0.46fF
C8958 nmat.col_n[24] ctopn 2.03fF
C8959 VDD a_11681_35823# 3.23fF
C8960 m2_17932_63982# m2_17932_62978# 0.99fF
C8961 a_2411_33749# a_4831_34561# 0.56fF
C8962 VDD pmat.col_n[17] 5.05fF
C8963 a_10441_21263# a_8443_20719# 2.68fF
C8964 a_37238_14512# a_37238_13508# 1.00fF
C8965 VDD a_26891_28327# 11.49fF
C8966 nmat.col_n[28] vcm 5.63fF
C8967 VDD a_11145_17999# 0.38fF
C8968 a_4068_25615# a_2683_22089# 0.46fF
C8969 VDD m2_51064_69002# 1.16fF
C8970 nmat.col[30] nmat.col[26] 2.10fF
C8971 a_18546_67216# a_38150_67174# 0.35fF
C8972 a_41254_57134# a_41254_56130# 1.00fF
C8973 a_9135_60967# a_10878_58487# 0.35fF
C8974 a_45270_19532# a_46274_19532# 0.97fF
C8975 pmat.col[22] m2_41024_54946# 0.39fF
C8976 pmat.row_n[5] a_10883_3303# 0.37fF
C8977 ANTENNA__1190__A2.DIODE nmat.col[7] 0.74fF
C8978 VDD a_25190_15516# 0.52fF
C8979 VDD a_4379_28548# 0.69fF
C8980 a_18546_7482# a_38150_7890# 0.35fF
C8981 VDD a_40969_30287# 0.52fF
C8982 a_6607_75895# a_6051_74183# 0.32fF
C8983 cgen.dlycontrol1_in[1] a_1858_25615# 0.71fF
C8984 a_44266_10496# a_45270_10496# 0.97fF
C8985 VDD a_11835_56311# 0.40fF
C8986 VDD pmat.rowoff_n[14] 1.87fF
C8987 VDD a_44266_12504# 0.52fF
C8988 cgen.dlycontrol3_in[0] a_11339_39319# 0.44fF
C8989 VDD m2_51064_8218# 1.05fF
C8990 nmat.col_n[16] a_35230_24552# 0.31fF
C8991 a_17996_35303# clk_dig 0.48fF
C8992 VDD _1184_.A2 19.29fF
C8993 pmat.row_n[12] a_18546_20534# 0.35fF
C8994 VDD a_9183_76359# 0.38fF
C8995 a_23182_21540# vcm 0.65fF
C8996 pmat.row_n[9] pmat.rowon_n[7] 0.81fF
C8997 VDD a_21174_60146# 0.52fF
C8998 cgen.dlycontrol2_in[0] cgen.dlycontrol1_in[4] 1.25fF
C8999 VDD a_46815_37013# 0.32fF
C9000 a_38242_58138# vcm 0.62fF
C9001 m2_46044_7214# m3_46176_7346# 2.79fF
C9002 a_5535_29980# a_10287_29941# 0.52fF
C9003 VDD a_18162_19532# 2.74fF
C9004 m2_17932_18258# m2_17932_17254# 0.99fF
C9005 nmat.col[27] m2_46044_24282# 0.40fF
C9006 m2_23956_54946# m3_24088_55078# 2.79fF
C9007 pmat.row_n[2] pmat.row_n[0] 15.26fF
C9008 a_18546_19530# a_27106_19938# 0.35fF
C9009 VDD a_20659_49140# 0.46fF
C9010 a_24186_12504# a_25190_12504# 0.97fF
C9011 a_18546_12502# a_31122_12910# 0.35fF
C9012 VDD comp.adc_inverter_1.in 0.40fF
C9013 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[24] 4.91fF
C9014 a_37238_22544# a_38242_22544# 0.97fF
C9015 VDD a_27198_16520# 0.52fF
C9016 a_49286_62154# pmat.col[30] 0.31fF
C9017 VDD pmat.col[22] 4.41fF
C9018 VDD a_37146_7890# 0.33fF
C9019 VDD a_8697_57167# 0.40fF
C9020 VDD a_12568_35077# 1.01fF
C9021 a_30210_69182# vcm 0.62fF
C9022 a_33467_46261# a_40949_48437# 0.45fF
C9023 a_18546_23546# a_36142_23954# 0.35fF
C9024 a_18546_16518# vcm 0.40fF
C9025 a_10515_13967# a_6467_29415# 4.22fF
C9026 VDD a_9411_2215# 17.75fF
C9027 a_18546_9490# a_40158_9898# 0.35fF
C9028 nmat.col_n[20] vcm 2.80fF
C9029 a_1957_43567# a_10883_3303# 0.77fF
C9030 VDD a_11797_60431# 1.92fF
C9031 a_39246_59142# vcm 0.62fF
C9032 VDD a_77980_40594# 0.36fF
C9033 a_2021_11043# a_8111_11209# 0.70fF
C9034 _1179_.X _1194_.A2 1.55fF
C9035 VDD a_7419_14379# 0.54fF
C9036 ANTENNA__1395__A1.DIODE a_21739_29415# 0.98fF
C9037 a_13145_26935# a_12449_22895# 0.43fF
C9038 pmat.en_bit_n[2] a_28704_29568# 1.66fF
C9039 a_2315_44124# a_2935_38279# 0.78fF
C9040 a_6927_30503# a_9761_30511# 0.61fF
C9041 a_41254_62154# pmat.col[22] 0.31fF
C9042 a_34226_56130# ctopp 3.46fF
C9043 VDD a_35039_29941# 0.38fF
C9044 a_10515_13967# a_13091_52047# 0.48fF
C9045 VDD a_43262_56130# 0.55fF
C9046 nmat.col[15] nmat.col[19] 1.23fF
C9047 VDD a_2191_25045# 0.56fF
C9048 a_26194_21540# ctopn 3.58fF
C9049 pmat.row_n[11] a_13091_18535# 7.73fF
C9050 a_20170_8488# a_21174_8488# 0.97fF
C9051 a_18546_65208# a_20078_65166# 0.35fF
C9052 VDD a_25190_22544# 0.52fF
C9053 a_37238_66170# ctopp 3.58fF
C9054 m2_38012_72014# m3_38144_72146# 2.79fF
C9055 pmat.rowoff_n[4] a_11067_30287# 0.31fF
C9056 VDD a_7939_31591# 3.08fF
C9057 VDD a_46274_66170# 0.52fF
C9058 a_46274_11500# a_47278_11500# 0.97fF
C9059 VDD a_15049_36374# 2.10fF
C9060 a_2411_43301# cgen.dlycontrol2_in[4] 0.72fF
C9061 a_30210_63158# ctopp 3.58fF
C9062 a_7415_29397# nmat.col_n[7] 0.46fF
C9063 cgen.dlycontrol3_in[4] a_14600_37607# 1.68fF
C9064 VDD a_39246_63158# 0.52fF
C9065 a_22178_17524# vcm 0.65fF
C9066 a_2659_35015# a_3911_44431# 0.36fF
C9067 cgen.dlycontrol3_in[0] a_2051_44111# 0.67fF
C9068 a_48282_64162# a_48282_63158# 1.00fF
C9069 a_18546_67216# a_20078_67174# 0.35fF
C9070 a_18546_61192# a_38150_61150# 0.35fF
C9071 nmat.col[29] m2_48052_24282# 0.39fF
C9072 m2_44036_54946# m2_45040_54946# 0.96fF
C9073 a_23182_8488# vcm 0.64fF
C9074 a_48282_58138# a_48282_57134# 1.00fF
C9075 VDD a_20075_43447# 0.62fF
C9076 VDD a_27794_28879# 0.39fF
C9077 a_39246_19532# vcm 0.65fF
C9078 a_40250_18528# a_40250_17524# 1.00fF
C9079 a_1858_25615# a_19605_32149# 0.33fF
C9080 cgen.dlycontrol1_in[4] cgen.dlycontrol1_in[2] 0.55fF
C9081 a_38242_10496# vcm 0.65fF
C9082 a_18546_13506# a_32126_13914# 0.35fF
C9083 VDD a_3956_72373# 0.65fF
C9084 a_11317_40188# a_11497_40719# 0.49fF
C9085 a_4075_50087# a_7563_63303# 0.58fF
C9086 a_40250_63158# a_40250_62154# 1.00fF
C9087 VDD a_4167_48463# 0.45fF
C9088 _1196_.B1 a_6467_29415# 0.65fF
C9089 a_35230_67174# ctopp 3.58fF
C9090 a_36234_55126# vcm 0.58fF
C9091 a_18546_18526# a_28110_18934# 0.35fF
C9092 a_16311_28327# a_45019_38645# 0.34fF
C9093 VDD a_44266_67174# 0.52fF
C9094 _1192_.B1 ANTENNA__1395__B1.DIODE 2.15fF
C9095 VDD a_4843_54826# 3.84fF
C9096 a_13597_37571# a_13503_36893# 0.63fF
C9097 a_14600_37607# a_12345_36924# 0.49fF
C9098 VDD a_2467_35925# 0.87fF
C9099 a_46274_22544# a_46274_21540# 1.00fF
C9100 a_23182_64162# ctopp 3.58fF
C9101 VDD a_22817_41317# 1.66fF
C9102 VDD a_33222_14512# 0.52fF
C9103 a_30210_56130# m2_29980_54946# 0.99fF
C9104 a_45270_14512# a_46274_14512# 0.97fF
C9105 VDD a_32218_64162# 0.52fF
C9106 a_28704_29568# a_28336_29967# 0.93fF
C9107 a_44266_64162# a_45270_64162# 0.97fF
C9108 a_18546_17522# a_50198_17930# 0.35fF
C9109 VDD a_21087_39913# 0.65fF
C9110 nmat.col_n[8] m2_26968_24282# 0.38fF
C9111 pmat.row_n[10] ctopn 1.65fF
C9112 VDD vcm.sky130_fd_sc_hd__dlymetal6s6s_1_5.X 0.42fF
C9113 pmat.rowoff_n[15] a_9463_50877# 1.04fF
C9114 pmat.row_n[2] nmat.sample 0.35fF
C9115 cgen.dlycontrol3_in[3] a_10873_39605# 2.52fF
C9116 a_18546_57176# a_46182_57134# 0.35fF
C9117 pmat.row_n[15] _1194_.A2 0.59fF
C9118 a_13091_28327# a_8583_29199# 0.33fF
C9119 a_39246_13508# a_39246_12504# 1.00fF
C9120 _1187_.A2 a_13459_28111# 0.35fF
C9121 ANTENNA__1190__A1.DIODE ANTENNA__1195__A1.DIODE 0.31fF
C9122 ANTENNA__1395__A2.DIODE a_21739_29415# 0.95fF
C9123 VDD a_12292_44869# 1.01fF
C9124 VDD nmat.col[13] 7.99fF
C9125 a_18546_15514# a_50198_15922# 0.35fF
C9126 VDD m2_48052_54946# 0.62fF
C9127 VDD a_6743_47081# 0.52fF
C9128 a_3175_59585# a_3136_59459# 0.42fF
C9129 a_8491_47911# a_8907_48437# 0.42fF
C9130 VDD a_1643_31573# 0.36fF
C9131 VDD a_9459_5461# 0.51fF
C9132 a_14249_49525# a_12044_49641# 0.42fF
C9133 a_25190_17524# ctopn 3.58fF
C9134 a_40250_11500# vcm 0.65fF
C9135 _1154_.A a_33467_46261# 0.41fF
C9136 _1154_.A ANTENNA__1184__B1.DIODE 0.57fF
C9137 a_2791_57703# a_4025_54965# 0.51fF
C9138 _1194_.A2 pmat.col[0] 0.55fF
C9139 cgen.dlycontrol4_in[4] a_11149_40188# 0.32fF
C9140 a_26194_8488# ctopn 3.40fF
C9141 m2_29980_54946# vcm 0.42fF
C9142 vcm.sky130_fd_sc_hd__buf_4_2.X vcm.sky130_fd_sc_hd__buf_4_3.X 0.58fF
C9143 a_23182_56130# a_24186_56130# 0.97fF
C9144 a_18546_56172# a_29114_56130# 0.35fF
C9145 VDD a_28110_24958# 0.44fF
C9146 m2_41024_24282# m2_42028_24282# 0.96fF
C9147 VDD a_2163_61761# 0.48fF
C9148 nmat.col[2] m2_20944_24282# 0.39fF
C9149 nmat.col_n[25] m2_44036_24282# 0.32fF
C9150 pmat.col_n[19] vcm 2.80fF
C9151 a_42258_19532# ctopn 3.58fF
C9152 a_26194_65166# ctopp 3.58fF
C9153 VDD a_40315_43177# 0.68fF
C9154 ANTENNA__1196__A2.DIODE a_9675_10396# 0.31fF
C9155 VDD a_35230_65166# 0.52fF
C9156 a_11897_21263# a_10959_23983# 0.96fF
C9157 a_28704_29568# nmat.col_n[12] 0.38fF
C9158 VDD a_42258_21540# 0.52fF
C9159 nmat.sw a_6007_33767# 2.53fF
C9160 a_46274_65166# a_46274_64162# 1.00fF
C9161 pmat.row_n[0] a_18546_8486# 0.35fF
C9162 a_41254_10496# ctopn 3.58fF
C9163 a_18546_68220# a_37146_68178# 0.35fF
C9164 _1179_.X a_32687_46607# 0.36fF
C9165 pmat.row_n[15] a_2411_43301# 0.62fF
C9166 a_2791_57703# a_5730_54965# 0.36fF
C9167 a_2835_13077# a_14195_7351# 0.93fF
C9168 a_48282_58138# ctopp 3.58fF
C9169 a_44266_68178# vcm 0.62fF
C9170 a_19541_28879# a_24602_48169# 0.73fF
C9171 VDD a_5768_9527# 1.31fF
C9172 VDD nmat.col_n[27] 5.17fF
C9173 cgen.enable_dlycontrol_in a_10873_36341# 1.10fF
C9174 a_17139_30503# a_43533_30761# 1.58fF
C9175 VDD a_3228_74691# 0.71fF
C9176 a_28202_62154# a_29206_62154# 0.97fF
C9177 a_35230_16520# a_35230_15516# 1.00fF
C9178 VDD a_40047_47919# 0.37fF
C9179 a_26194_66170# a_27198_66170# 0.97fF
C9180 a_18546_60188# a_42166_60146# 0.35fF
C9181 a_19166_66170# ctopp 3.43fF
C9182 a_21174_12504# ctopn 3.58fF
C9183 VDD a_8243_7290# 1.07fF
C9184 VDD a_17675_37001# 1.08fF
C9185 a_6559_33767# a_9213_53903# 0.52fF
C9186 a_15101_29423# a_10147_29415# 0.90fF
C9187 pmat.col[17] vcm 5.88fF
C9188 a_4075_50087# a_7467_63303# 0.58fF
C9189 a_11067_64015# pmat.rowoff_n[4] 0.57fF
C9190 a_18546_63200# a_21082_63158# 0.35fF
C9191 VDD m2_33996_72014# 1.00fF
C9192 a_11927_27399# a_7840_27247# 0.78fF
C9193 a_49286_23548# vcm 0.65fF
C9194 a_18546_61192# a_20078_61150# 0.35fF
C9195 a_40250_69182# ctopp 3.58fF
C9196 ANTENNA__1196__A2.DIODE a_21739_29415# 0.32fF
C9197 pmat.col[8] ctopp 1.97fF
C9198 a_20170_66170# vcm 0.62fF
C9199 VDD a_49286_69182# 0.52fF
C9200 a_17139_30503# a_8583_29199# 0.34fF
C9201 m2_29980_72014# m2_30984_72014# 0.96fF
C9202 VDD a_23479_39095# 0.64fF
C9203 a_50290_59142# m2_51064_58962# 0.96fF
C9204 a_13183_72405# a_13349_72405# 0.53fF
C9205 pmat.col_n[14] m2_32992_54946# 0.37fF
C9206 VDD a_8051_46607# 0.40fF
C9207 nmat.col_n[5] vcm 2.80fF
C9208 a_47278_65166# a_48282_65166# 0.97fF
C9209 a_49286_59142# ctopp 3.57fF
C9210 a_1858_25615# a_5087_32687# 0.63fF
C9211 a_43262_11500# ctopn 3.58fF
C9212 _1154_.A ANTENNA_fanout52_A.DIODE 5.05fF
C9213 m3_50768_24414# ctopn 0.39fF
C9214 ANTENNA__1187__B1.DIODE a_15667_27239# 3.55fF
C9215 a_20170_10496# vcm 0.65fF
C9216 VDD a_11877_12565# 0.64fF
C9217 VDD m2_17932_11230# 1.12fF
C9218 a_4128_64391# a_7373_49007# 0.47fF
C9219 VDD a_18203_48981# 0.33fF
C9220 pmat.rowoff_n[7] nmat.rowoff_n[13] 0.55fF
C9221 pmat.rowoff_n[8] ctopp 0.60fF
C9222 a_26194_61150# ctopp 3.58fF
C9223 a_27198_70186# a_28202_70186# 0.97fF
C9224 VDD a_1895_8378# 0.43fF
C9225 VDD a_35230_61150# 0.52fF
C9226 a_13459_28111# pmat.col[1] 0.36fF
C9227 VDD a_25301_40229# 1.43fF
C9228 nmat.sw a_3351_27249# 0.84fF
C9229 a_47278_13508# vcm 0.65fF
C9230 a_19166_18528# ctopn 3.43fF
C9231 a_29163_29423# a_28336_29967# 1.55fF
C9232 nmat.col_n[12] a_12851_28853# 0.44fF
C9233 a_45270_18528# vcm 0.65fF
C9234 VDD a_29206_20536# 0.52fF
C9235 VDD a_10409_53903# 0.41fF
C9236 a_18546_71232# a_26102_71190# 0.35fF
C9237 a_16311_28327# nmat.sw 1.19fF
C9238 a_5784_52423# a_2411_43301# 0.82fF
C9239 a_29206_23548# m2_28976_24282# 0.99fF
C9240 a_19166_22544# a_20170_22544# 0.97fF
C9241 VDD a_41254_17524# 0.52fF
C9242 VDD nmat.col[24] 6.73fF
C9243 pmat.rowoff_n[7] vcm 0.83fF
C9244 a_9963_13967# a_8197_20871# 0.43fF
C9245 ANTENNA_fanout52_A.DIODE a_11711_50959# 0.33fF
C9246 VDD a_28455_47381# 0.43fF
C9247 a_18546_8486# a_34134_8894# 0.35fF
C9248 VDD a_5547_77295# 0.41fF
C9249 a_20170_60146# a_20170_59142# 1.00fF
C9250 a_18546_65208# a_31122_65166# 0.35fF
C9251 VDD a_42258_8488# 0.55fF
C9252 a_7779_22583# a_4703_24527# 0.42fF
C9253 a_9217_23983# nmat.col_n[1] 0.42fF
C9254 VDD a_2124_59067# 0.66fF
C9255 a_18546_21538# a_45178_21946# 0.35fF
C9256 pmat.row_n[5] pmat.row_n[3] 0.63fF
C9257 a_38242_62154# a_38242_61150# 1.00fF
C9258 a_12461_29673# a_13655_26703# 0.66fF
C9259 a_35312_31599# a_17842_27497# 0.31fF
C9260 a_30571_50959# a_43776_30287# 0.42fF
C9261 a_26891_28327# a_43533_30761# 1.01fF
C9262 nmat.col_n[21] comp_latch 1.55fF
C9263 a_18563_27791# a_24747_29967# 1.28fF
C9264 VDD nmat.rowon_n[13] 3.37fF
C9265 a_24186_67174# a_25190_67174# 0.97fF
C9266 a_18546_67216# a_31122_67174# 0.35fF
C9267 VDD a_18162_24552# 27.53fF
C9268 VDD config_2_in[13] 1.40fF
C9269 a_8583_29199# a_11927_27399# 0.42fF
C9270 a_28704_29568# nmat.col_n[18] 1.35fF
C9271 a_21174_66170# a_21174_65166# 1.00fF
C9272 a_26891_28327# a_22499_49783# 0.58fF
C9273 VDD a_11910_43047# 0.40fF
C9274 VDD a_6835_14735# 0.50fF
C9275 nmat.rowon_n[9] nmat.rowoff_n[9] 20.45fF
C9276 a_38242_15516# a_38242_14512# 1.00fF
C9277 a_13459_28111# nmat.col_n[11] 0.82fF
C9278 a_18546_7482# a_31122_7890# 0.35fF
C9279 a_40250_69182# a_40250_68178# 1.00fF
C9280 a_18546_68220# a_18162_68218# 2.62fF
C9281 VDD pmat.rowon_n[0] 16.52fF
C9282 a_48282_21540# a_48282_20536# 1.00fF
C9283 a_6283_31591# a_32687_46607# 1.70fF
C9284 VDD result_out[6] 0.70fF
C9285 VDD a_37238_12504# 0.52fF
C9286 _1184_.A2 a_4523_21276# 0.71fF
C9287 a_45019_38645# a_45915_29941# 0.75fF
C9288 a_19166_62154# a_20170_62154# 0.97fF
C9289 VDD a_40677_48437# 0.62fF
C9290 a_50290_13508# ctopn 3.43fF
C9291 nmat.rowon_n[14] nmat.rowoff_n[14] 20.71fF
C9292 a_2021_11043# a_9460_10615# 0.30fF
C9293 a_45270_57134# vcm 0.62fF
C9294 a_44266_71190# vcm 0.60fF
C9295 a_48282_18528# ctopn 3.58fF
C9296 a_24407_31375# a_9785_28879# 2.25fF
C9297 a_31214_58138# vcm 0.62fF
C9298 _1184_.A2 a_22499_49783# 0.32fF
C9299 a_28915_50959# a_30663_50087# 0.33fF
C9300 a_11892_21959# a_5899_21807# 0.61fF
C9301 ANTENNA__1190__B1.DIODE ANTENNA__1183__B1.DIODE 2.45fF
C9302 VDD vcm.sky130_fd_sc_hd__buf_4_0.X 0.82fF
C9303 a_1769_13103# config_1_in[13] 0.45fF
C9304 pmat.col_n[1] pmat.col[1] 0.68fF
C9305 a_7803_67655# a_7899_67477# 0.36fF
C9306 nmat.col_n[12] ANTENNA__1190__A2.DIODE 0.58fF
C9307 a_12069_38517# a_22153_37179# 1.54fF
C9308 pmat.col_n[9] ANTENNA__1197__A.DIODE 0.43fF
C9309 a_18546_12502# a_24094_12910# 0.35fF
C9310 VDD m3_47180_7346# 0.39fF
C9311 VDD a_30641_44743# 1.22fF
C9312 a_2411_43301# a_5639_49007# 0.34fF
C9313 VDD m2_38012_24282# 0.62fF
C9314 a_2648_29397# a_6559_8527# 0.38fF
C9315 a_23821_35279# a_29159_37607# 1.05fF
C9316 VDD nmat.col_n[22] 5.26fF
C9317 VDD a_42240_29423# 0.78fF
C9318 VDD a_30118_7890# 0.33fF
C9319 pmat.col_n[27] ctopp 2.02fF
C9320 a_42258_11500# a_42258_10496# 1.00fF
C9321 a_23182_69182# vcm 0.62fF
C9322 VDD a_2727_58470# 3.89fF
C9323 _1194_.B1 a_11067_30287# 0.33fF
C9324 a_18546_23546# a_29114_23954# 0.35fF
C9325 a_23182_23548# a_24186_23548# 0.97fF
C9326 ANTENNA__1183__B1.DIODE a_14365_22351# 0.51fF
C9327 a_13275_48783# a_40628_39429# 0.40fF
C9328 a_10055_31591# ANTENNA__1196__A2.DIODE 0.45fF
C9329 a_11497_38543# a_14600_37607# 0.96fF
C9330 a_18546_9490# a_33130_9898# 0.35fF
C9331 a_25190_9492# a_26194_9492# 0.97fF
C9332 a_47278_61150# a_48282_61150# 0.97fF
C9333 pmat.rowon_n[14] a_18162_70226# 1.19fF
C9334 a_18546_70228# a_19074_70186# 0.35fF
C9335 a_32218_59142# vcm 0.62fF
C9336 a_32218_12504# a_32218_11500# 1.00fF
C9337 nmat.rowon_n[7] a_10515_13967# 0.46fF
C9338 pmat.rowon_n[6] vcm 0.58fF
C9339 a_18546_55168# a_18162_55166# 2.55fF
C9340 a_38851_28327# a_37820_30485# 0.98fF
C9341 a_22499_49783# a_9411_2215# 0.93fF
C9342 pmat.rowon_n[3] a_2411_43301# 0.59fF
C9343 a_27198_56130# ctopp 3.40fF
C9344 VDD a_36234_56130# 0.54fF
C9345 a_41254_20536# a_42258_20536# 0.97fF
C9346 pmat.row_n[5] pmat.row_n[1] 13.91fF
C9347 _1224_.X clk_ena 4.55fF
C9348 VDD a_1761_9839# 0.59fF
C9349 a_18546_72236# a_30118_72194# 0.35fF
C9350 VDD m3_32120_72146# 0.33fF
C9351 a_9411_2215# a_8583_29199# 1.09fF
C9352 a_17996_41831# a_17625_42902# 0.51fF
C9353 a_18546_62196# a_50198_62154# 0.35fF
C9354 ANTENNA__1395__A1.DIODE a_24867_53135# 1.21fF
C9355 a_18546_66212# a_46182_66170# 0.35fF
C9356 a_40250_9492# a_40250_8488# 1.00fF
C9357 a_30210_66170# ctopp 3.58fF
C9358 a_1586_50247# a_1591_50095# 0.34fF
C9359 VDD a_39246_66170# 0.52fF
C9360 a_22178_21540# a_23182_21540# 0.97fF
C9361 VDD a_34887_36919# 0.63fF
C9362 nmat.sw a_18975_40871# 1.14fF
C9363 a_23182_63158# ctopp 3.58fF
C9364 a_10883_3303# nmat.col_n[13] 0.70fF
C9365 VDD a_32218_63158# 0.52fF
C9366 a_2952_25045# a_3305_27791# 0.81fF
C9367 a_18546_61192# a_31122_61150# 0.35fF
C9368 m2_37008_54946# m2_38012_54946# 0.96fF
C9369 a_23182_71190# a_23182_70186# 1.00fF
C9370 a_37238_58138# a_38242_58138# 0.97fF
C9371 a_11067_64015# a_11067_16359# 2.29fF
C9372 VDD a_10867_43447# 0.59fF
C9373 VDD a_31631_51701# 0.76fF
C9374 a_32218_19532# vcm 0.65fF
C9375 a_5682_56311# a_11902_56775# 0.32fF
C9376 VDD a_21815_34191# 0.31fF
C9377 a_31214_10496# vcm 0.65fF
C9378 a_18546_13506# a_25098_13914# 0.35fF
C9379 a_21174_13508# a_22178_13508# 0.97fF
C9380 VDD a_1644_72917# 0.31fF
C9381 a_5651_66975# a_9463_50877# 0.53fF
C9382 nmat.col[14] ctopn 1.97fF
C9383 a_3339_59879# a_11067_16359# 0.33fF
C9384 a_32218_71190# m2_31988_72014# 1.00fF
C9385 _1192_.A2 vcm 1.25fF
C9386 nmat.rowon_n[14] vcm 0.53fF
C9387 VDD a_26242_49257# 0.47fF
C9388 a_37238_61150# a_37238_60146# 1.00fF
C9389 a_28202_67174# ctopp 3.58fF
C9390 nmat.col_n[3] a_3571_13627# 0.98fF
C9391 VDD a_32035_38825# 0.64fF
C9392 a_45270_19532# a_45270_18528# 1.00fF
C9393 a_3576_17143# clk_dig 0.71fF
C9394 a_18546_70228# a_48190_70186# 0.35fF
C9395 VDD a_37238_67174# 0.52fF
C9396 a_19166_11500# a_20170_11500# 0.97fF
C9397 VDD a_34924_37253# 1.32fF
C9398 VDD a_11261_41245# 1.23fF
C9399 VDD a_26194_14512# 0.52fF
C9400 a_47278_62154# vcm 0.62fF
C9401 VDD a_25190_64162# 0.52fF
C9402 inn_analog nmat.col[28] 2.88fF
C9403 nmat.col_n[18] ANTENNA__1190__A2.DIODE 2.13fF
C9404 a_11067_49871# a_11067_30287# 0.60fF
C9405 VDD a_7079_40277# 0.60fF
C9406 a_18546_17522# a_43170_17930# 0.35fF
C9407 pmat.rowon_n[0] pmat.rowoff_n[1] 1.09fF
C9408 a_18546_57176# a_39154_57134# 0.35fF
C9409 a_13529_34951# cgen.dlycontrol1_in[3] 0.43fF
C9410 VDD vcm.sky130_fd_sc_hd__nand2_1_1.A 0.79fF
C9411 VDD a_13073_54997# 0.39fF
C9412 a_38242_59142# a_38242_58138# 1.00fF
C9413 _1194_.B1 _1192_.A2 2.18fF
C9414 a_6451_67655# a_5081_53135# 1.30fF
C9415 a_1674_57711# a_10239_14183# 0.82fF
C9416 pmat.rowoff_n[8] pmat.rowon_n[7] 1.01fF
C9417 pmat.rowoff_n[12] start_conversion_in 0.37fF
C9418 a_30210_15516# a_31214_15516# 0.97fF
C9419 a_18546_15514# a_43170_15922# 0.35fF
C9420 a_4351_55527# a_4025_54965# 1.08fF
C9421 a_29206_69182# a_30210_69182# 0.97fF
C9422 VDD a_1761_7119# 0.71fF
C9423 VDD a_22357_35877# 1.32fF
C9424 a_46274_70186# vcm 0.62fF
C9425 VDD pmat.col_n[20] 5.49fF
C9426 a_33222_11500# vcm 0.65fF
C9427 VDD a_4075_31591# 14.04fF
C9428 VDD a_12985_62581# 0.65fF
C9429 a_23395_53135# _1192_.B1 1.03fF
C9430 ANTENNA__1187__B1.DIODE a_11067_27239# 6.05fF
C9431 ANTENNA__1197__B.DIODE a_24591_28327# 0.41fF
C9432 a_2263_43719# a_14887_46377# 1.85fF
C9433 a_43262_17524# a_43262_16520# 1.00fF
C9434 a_18162_8488# ctopn 1.30fF
C9435 a_30663_50087# a_30111_47911# 0.88fF
C9436 ctopp ctopn 2.23fF
C9437 a_18546_56172# a_22086_56130# 0.35fF
C9438 pmat.row_n[15] a_11897_21263# 0.31fF
C9439 inn_analog m2_50060_24282# 0.71fF
C9440 VDD a_20170_24552# 0.60fF
C9441 a_8439_69653# a_9135_69679# 0.63fF
C9442 a_10515_61839# nmat.en_bit_n[1] 7.95fF
C9443 a_49286_12504# a_50290_12504# 0.97fF
C9444 VDD a_10641_52815# 0.64fF
C9445 a_35230_19532# ctopn 3.58fF
C9446 VDD a_22541_43131# 1.44fF
C9447 a_1823_74557# a_2124_69947# 0.37fF
C9448 a_18546_14510# a_18162_14512# 2.61fF
C9449 VDD a_28202_65166# 0.52fF
C9450 a_2007_25597# a_20310_28029# 0.72fF
C9451 pmat.row_n[6] a_18162_14512# 25.57fF
C9452 VDD a_10957_28879# 0.32fF
C9453 ANTENNA__1190__B1.DIODE a_38913_31055# 0.62fF
C9454 VDD a_35230_21540# 0.52fF
C9455 a_38242_59142# a_39246_59142# 0.97fF
C9456 a_34226_10496# ctopn 3.58fF
C9457 a_18546_68220# a_30118_68178# 0.35fF
C9458 VDD a_23352_30761# 0.44fF
C9459 a_41254_58138# ctopp 3.58fF
C9460 a_37238_68178# vcm 0.62fF
C9461 VDD a_6179_69831# 0.53fF
C9462 a_11067_30287# a_8749_47381# 0.55fF
C9463 VDD a_50290_58138# 0.54fF
C9464 nmat.sw a_6467_29415# 2.80fF
C9465 a_27198_23548# a_27198_22544# 1.00fF
C9466 VDD pmat.col[24] 4.43fF
C9467 VDD a_6051_74183# 1.61fF
C9468 a_26194_60146# a_27198_60146# 0.97fF
C9469 a_18546_60188# a_35138_60146# 0.35fF
C9470 VDD a_51202_23954# 0.30fF
C9471 m2_51064_19262# m2_51064_20266# 0.99fF
C9472 pmat.row_n[8] nmat.sample 0.35fF
C9473 m2_51064_7214# m3_51196_7346# 2.79fF
C9474 VDD a_7364_63303# 0.37fF
C9475 comp.adc_nor_latch_0.QN comp_latch 1.08fF
C9476 nmat.col[1] a_3571_13627# 0.37fF
C9477 a_45019_38645# a_44757_37289# 0.41fF
C9478 m2_28976_54946# m3_29108_55078# 2.79fF
C9479 VDD m2_19940_72014# 1.16fF
C9480 a_34226_68178# a_34226_67174# 1.00fF
C9481 a_15660_31029# clk_ena 0.37fF
C9482 a_42258_23548# vcm 0.65fF
C9483 a_33222_69182# ctopp 3.58fF
C9484 a_44266_9492# vcm 0.65fF
C9485 VDD a_42258_69182# 0.52fF
C9486 pmat.row_n[11] cgen.dlycontrol2_in[3] 0.53fF
C9487 m2_22952_72014# m2_23956_72014# 0.96fF
C9488 a_37820_30485# a_37827_30793# 0.46fF
C9489 VDD a_15420_44007# 1.15fF
C9490 a_20170_15516# a_20170_14512# 1.00fF
C9491 pmat.col_n[10] m2_28976_54946# 0.37fF
C9492 VDD a_36532_46805# 0.49fF
C9493 VDD a_2715_51969# 0.44fF
C9494 pmat.rowon_n[8] a_1957_43567# 1.11fF
C9495 a_42258_59142# ctopp 3.58fF
C9496 VDD a_20267_27497# 0.38fF
C9497 a_36234_11500# ctopn 3.58fF
C9498 a_13091_28327# nmat.col[15] 1.19fF
C9499 _1154_.X _1192_.A2 2.27fF
C9500 _1154_.A a_13091_28327# 0.34fF
C9501 _1179_.X ANTENNA__1197__B.DIODE 2.56fF
C9502 _1192_.B1 a_46027_44905# 0.50fF
C9503 a_24867_53135# ANTENNA__1196__A2.DIODE 1.32fF
C9504 a_33467_46261# a_43315_48437# 0.36fF
C9505 ANTENNA__1197__B.DIODE a_33423_47695# 0.69fF
C9506 a_32218_16520# a_33222_16520# 0.97fF
C9507 a_18546_16518# a_47186_16926# 0.35fF
C9508 m2_43032_24282# vcm 0.42fF
C9509 a_22178_67174# a_22178_66170# 1.00fF
C9510 a_10595_53361# a_10409_53903# 0.59fF
C9511 pmat.row_n[10] ctopp 1.65fF
C9512 a_10589_22351# nmat.col_n[13] 0.36fF
C9513 VDD a_19166_67174# 0.56fF
C9514 a_2419_53351# a_4081_61127# 0.36fF
C9515 VDD a_28202_61150# 0.52fF
C9516 a_2199_13887# a_1591_8213# 0.34fF
C9517 nmat.col[31] a_31339_31787# 1.19fF
C9518 VDD a_25879_31591# 8.94fF
C9519 a_40250_13508# vcm 0.65fF
C9520 VDD a_39321_42333# 1.18fF
C9521 a_38905_28853# a_41237_28585# 0.39fF
C9522 a_21739_29415# a_31339_31787# 0.50fF
C9523 VDD a_1895_63866# 0.89fF
C9524 a_20616_27791# nmat.col[10] 1.95fF
C9525 a_38242_18528# vcm 0.65fF
C9526 VDD a_22178_20536# 0.52fF
C9527 a_21174_17524# a_22178_17524# 0.97fF
C9528 pmat.row_n[7] pmat.row_n[5] 1.58fF
C9529 a_2407_49289# a_1769_13103# 0.37fF
C9530 a_4351_55527# a_2407_49289# 0.49fF
C9531 _1179_.X a_31675_47695# 0.37fF
C9532 a_24186_20536# a_24186_19532# 1.00fF
C9533 m2_51064_58962# m2_51064_57958# 0.99fF
C9534 a_33423_47695# a_31675_47695# 1.25fF
C9535 a_49286_15516# vcm 0.65fF
C9536 VDD a_34226_17524# 0.52fF
C9537 a_22178_8488# a_23182_8488# 0.97fF
C9538 a_18546_8486# a_27106_8894# 0.35fF
C9539 a_18546_65208# a_24094_65166# 0.35fF
C9540 m2_43032_72014# m3_43164_72146# 2.79fF
C9541 VDD a_14839_20871# 1.05fF
C9542 a_41254_70186# a_41254_69182# 1.00fF
C9543 VDD a_35230_8488# 0.55fF
C9544 a_18546_21538# a_38150_21946# 0.35fF
C9545 VDD a_22085_36374# 1.13fF
C9546 a_30210_14512# a_30210_13508# 1.00fF
C9547 a_45270_23548# ctopn 3.40fF
C9548 a_35230_56130# a_35230_55126# 1.00fF
C9549 a_47278_9492# ctopn 3.57fF
C9550 a_27763_27221# nmat.col_n[31] 0.36fF
C9551 a_18546_67216# a_24094_67174# 0.35fF
C9552 a_34226_57134# a_34226_56130# 1.00fF
C9553 pmat.rowon_n[12] ctopp 1.57fF
C9554 VDD a_10959_23983# 1.52fF
C9555 ANTENNA__1195__A1.DIODE nmat.col[12] 0.38fF
C9556 a_38242_19532# a_39246_19532# 0.97fF
C9557 a_34204_27765# nmat.col_n[19] 0.38fF
C9558 a_45270_60146# vcm 0.62fF
C9559 nmat.rowon_n[7] a_2835_13077# 1.23fF
C9560 VDD a_50290_10496# 0.54fF
C9561 a_10873_38517# a_11225_35836# 0.92fF
C9562 a_28915_50959# a_10883_3303# 1.02fF
C9563 a_11041_40948# a_21981_34191# 1.18fF
C9564 a_19166_57134# m2_18936_55950# 0.99fF
C9565 a_2411_43301# a_4128_46983# 0.39fF
C9566 a_1781_9308# a_5131_13255# 0.37fF
C9567 a_18546_7482# a_24094_7890# 0.35fF
C9568 VDD a_7644_16341# 4.28fF
C9569 pmat.rowon_n[0] a_4523_21276# 0.75fF
C9570 a_18243_28327# a_15667_27239# 1.30fF
C9571 VDD a_47011_31029# 0.64fF
C9572 a_17139_30503# nmat.col[15] 0.39fF
C9573 a_37238_10496# a_38242_10496# 0.97fF
C9574 a_19166_68178# vcm 0.61fF
C9575 VDD a_30210_12504# 0.52fF
C9576 a_11067_16359# a_3571_13627# 0.31fF
C9577 a_2149_45717# a_1586_63927# 1.37fF
C9578 a_2879_57487# a_3866_57399# 1.73fF
C9579 VDD a_13349_72405# 0.63fF
C9580 a_2149_45717# a_1769_47919# 1.81fF
C9581 a_9135_60967# nmat.sw 0.91fF
C9582 a_48282_56130# a_49286_56130# 0.97fF
C9583 a_43262_13508# ctopn 3.58fF
C9584 _1196_.B1 ANTENNA__1187__B1.DIODE 0.90fF
C9585 VDD a_10058_60431# 0.51fF
C9586 pmat.col[15] vcm 5.88fF
C9587 a_38242_57134# vcm 0.62fF
C9588 a_37238_71190# vcm 0.60fF
C9589 a_10515_15055# a_9963_13967# 3.38fF
C9590 a_41254_18528# ctopn 3.58fF
C9591 VDD a_33765_41317# 1.18fF
C9592 a_24186_58138# vcm 0.62fF
C9593 a_13459_28111# a_25695_28111# 0.31fF
C9594 ANTENNA__1196__A2.DIODE a_38851_28327# 0.31fF
C9595 m2_50060_24282# clk_ena 0.56fF
C9596 VDD a_29159_39783# 0.56fF
C9597 a_2163_61761# a_2124_61635# 0.75fF
C9598 m2_17932_55950# m2_18936_55950# 0.96fF
C9599 VDD m3_19068_7346# 0.37fF
C9600 a_30210_22544# a_31214_22544# 0.97fF
C9601 VDD config_1_in[15] 1.32fF
C9602 VDD a_13985_44581# 1.33fF
C9603 VDD a_8767_16055# 0.52fF
C9604 pmat.row_n[4] a_1586_18231# 0.38fF
C9605 nmat.rowoff_n[6] a_7717_14735# 1.08fF
C9606 a_3746_58487# a_4707_32156# 0.32fF
C9607 a_17139_30503# a_11711_50959# 1.16fF
C9608 pmat.row_n[3] pmat.row_n[2] 2.08fF
C9609 VDD nmat.col_n[9] 5.44fF
C9610 a_4583_68021# a_4075_68583# 0.36fF
C9611 VDD a_14287_31599# 0.38fF
C9612 VDD a_23090_7890# 0.34fF
C9613 a_2419_69455# a_4081_61127# 0.36fF
C9614 VDD a_1775_35113# 0.45fF
C9615 a_18546_23546# a_22086_23954# 0.35fF
C9616 ANTENNA__1197__A.DIODE a_36453_29199# 0.34fF
C9617 VDD ndecision_finish 7.79fF
C9618 a_44266_63158# a_45270_63158# 0.97fF
C9619 m2_39016_54946# vcm 0.42fF
C9620 a_18546_9490# a_26102_9898# 0.35fF
C9621 a_49286_22544# vcm 0.65fF
C9622 a_19166_61150# a_19166_60146# 1.00fF
C9623 a_47278_68178# ctopp 3.58fF
C9624 ANTENNA__1183__B1.DIODE nmat.col[26] 0.46fF
C9625 VDD a_7899_67477# 0.66fF
C9626 a_40105_47375# a_7109_29423# 1.86fF
C9627 a_25190_59142# vcm 0.62fF
C9628 a_34226_55126# m2_32992_54946# 0.96fF
C9629 pmat.col_n[22] vcm 2.80fF
C9630 a_24407_31375# nmat.sw 1.46fF
C9631 a_32687_46607# a_28336_29967# 0.88fF
C9632 nmat.col[25] nmat.col[26] 0.45fF
C9633 a_20170_18528# vcm 0.65fF
C9634 a_20170_56130# ctopp 3.28fF
C9635 a_1923_69823# a_3136_72515# 0.30fF
C9636 VDD a_29206_56130# 0.55fF
C9637 a_6283_31591# a_31675_47695# 0.98fF
C9638 a_22178_8488# m2_21948_7214# 1.00fF
C9639 VDD a_18162_70226# 2.73fF
C9640 VDD m2_46044_7214# 0.93fF
C9641 a_6283_31591# a_24374_29941# 0.38fF
C9642 a_10781_42869# a_14497_42658# 1.36fF
C9643 VDD a_12815_74581# 0.54fF
C9644 a_18546_62196# a_43170_62154# 0.35fF
C9645 a_18546_66212# a_39154_66170# 0.35fF
C9646 a_23182_66170# ctopp 3.58fF
C9647 a_22199_30287# nmat.col_n[26] 0.46fF
C9648 _1154_.A a_26891_28327# 1.31fF
C9649 VDD a_7387_33231# 0.45fF
C9650 VDD a_32218_66170# 0.52fF
C9651 a_39246_11500# a_40250_11500# 0.97fF
C9652 ANTENNA__1197__A.DIODE nmat.col_n[31] 1.28fF
C9653 pmat.row_n[13] pmat.row_n[7] 0.77fF
C9654 VDD a_25190_63158# 0.52fF
C9655 pmat.en_bit_n[2] a_22216_30761# 0.32fF
C9656 a_41254_64162# a_41254_63158# 1.00fF
C9657 m2_51064_59966# vcm 0.51fF
C9658 a_44266_10496# a_44266_9492# 1.00fF
C9659 a_18546_61192# a_24094_61150# 0.35fF
C9660 a_41254_58138# a_41254_57134# 1.00fF
C9661 VDD a_33765_39141# 1.18fF
C9662 a_4257_34319# a_4307_35639# 0.40fF
C9663 VDD a_46950_43719# 0.52fF
C9664 m2_17932_16250# m3_18064_16382# 2.76fF
C9665 a_25190_19532# vcm 0.65fF
C9666 a_45270_60146# a_45270_59142# 1.00fF
C9667 a_33222_18528# a_33222_17524# 1.00fF
C9668 cgen.dlycontrol1_in[2] a_3091_33402# 0.52fF
C9669 a_18546_71232# ctopp 1.30fF
C9670 _1154_.A _1184_.A2 0.49fF
C9671 a_28901_48437# a_30189_48437# 0.52fF
C9672 a_24186_10496# vcm 0.65fF
C9673 ANTENNA__1197__B.DIODE nmat.sample_n 2.91fF
C9674 a_33222_63158# a_33222_62154# 1.00fF
C9675 nmat.rowoff_n[1] ctopn 0.60fF
C9676 a_49286_67174# a_50290_67174# 0.97fF
C9677 a_10239_14183# a_4383_7093# 0.44fF
C9678 a_1823_60949# a_3136_59459# 0.59fF
C9679 VDD a_2907_22522# 0.41fF
C9680 VDD a_13801_38779# 1.25fF
C9681 a_21174_67174# ctopp 3.58fF
C9682 VDD a_24591_28327# 13.85fF
C9683 a_18546_70228# a_41162_70186# 0.35fF
C9684 VDD a_30210_67174# 0.52fF
C9685 _1192_.A2 a_40837_46261# 0.47fF
C9686 pmat.rowon_n[8] a_2411_33749# 1.43fF
C9687 VDD a_12309_38659# 4.98fF
C9688 a_14600_37607# a_14712_37429# 0.35fF
C9689 a_39246_22544# a_39246_21540# 1.00fF
C9690 a_46274_66170# a_46274_65166# 1.00fF
C9691 a_19166_71190# vcm 0.60fF
C9692 pmat.rowoff_n[15] a_10883_3303# 1.35fF
C9693 VDD a_29036_41831# 1.30fF
C9694 VDD a_18162_14512# 2.74fF
C9695 a_9581_56079# a_9213_53903# 0.46fF
C9696 a_38242_14512# a_39246_14512# 0.97fF
C9697 a_40250_62154# vcm 0.62fF
C9698 nmat.col[29] nmat.col_n[24] 3.96fF
C9699 pmat.row_n[2] pmat.row_n[1] 5.10fF
C9700 a_18546_17522# a_36142_17930# 0.35fF
C9701 a_37238_64162# a_38242_64162# 0.97fF
C9702 a_43262_68178# a_44266_68178# 0.97fF
C9703 a_18546_57176# a_32126_57134# 0.35fF
C9704 pmat.col[12] m2_30984_54946# 0.40fF
C9705 a_41254_8488# m2_41024_7214# 1.00fF
C9706 a_32218_13508# a_32218_12504# 1.00fF
C9707 pmat.rowoff_n[12] nmat.rowon_n[7] 3.59fF
C9708 pmat.row_n[11] pmat.row_n[7] 3.06fF
C9709 a_6283_31591# a_14691_27399# 0.43fF
C9710 a_18546_15514# a_36142_15922# 0.35fF
C9711 VDD m2_17932_54946# 1.28fF
C9712 VDD a_32371_47349# 0.53fF
C9713 VDD a_6200_70919# 3.84fF
C9714 a_1923_61759# a_2163_67645# 0.32fF
C9715 VDD a_27443_32143# 0.51fF
C9716 VDD a_6559_57167# 0.35fF
C9717 nmat.col_n[23] ctopn 2.02fF
C9718 a_39246_70186# vcm 0.62fF
C9719 a_9411_2215# nmat.col[15] 0.72fF
C9720 a_26194_11500# vcm 0.65fF
C9721 _1154_.A a_9411_2215# 0.62fF
C9722 a_13459_28111# a_12987_26159# 1.52fF
C9723 ANTENNA__1183__B1.DIODE clk_ena 0.91fF
C9724 a_5731_58951# a_5682_56311# 0.31fF
C9725 VDD a_13768_22325# 0.71fF
C9726 pmat.rowon_n[7] a_4707_32156# 2.28fF
C9727 a_28202_19532# ctopn 3.58fF
C9728 VDD cgen.dlycontrol2_in[4] 5.77fF
C9729 nmat.col[11] nmat.col_n[11] 0.75fF
C9730 m2_17932_13238# m3_18064_13370# 2.76fF
C9731 VDD a_21174_65166# 0.52fF
C9732 a_2419_69455# a_2935_38279# 0.41fF
C9733 a_10239_14183# a_14457_15823# 0.61fF
C9734 VDD a_43659_28853# 0.77fF
C9735 a_2407_49289# a_3339_70759# 0.74fF
C9736 VDD a_28202_21540# 0.52fF
C9737 a_39246_65166# a_39246_64162# 1.00fF
C9738 a_27198_10496# ctopn 3.58fF
C9739 a_48282_57134# ctopp 3.57fF
C9740 a_18546_68220# a_23090_68178# 0.35fF
C9741 a_47278_71190# ctopp 3.40fF
C9742 a_10515_13967# a_2683_22089# 0.53fF
C9743 a_34226_58138# ctopp 3.58fF
C9744 a_30210_68178# vcm 0.62fF
C9745 VDD a_43262_58138# 0.52fF
C9746 a_48282_23548# a_49286_23548# 0.97fF
C9747 VDD _1179_.X 19.97fF
C9748 a_28202_16520# a_28202_15516# 1.00fF
C9749 a_21174_62154# a_22178_62154# 0.97fF
C9750 m2_51064_15246# m2_51064_14242# 0.99fF
C9751 a_12987_26159# a_6829_26703# 0.69fF
C9752 VDD a_33423_47695# 12.89fF
C9753 a_8481_10396# comp_latch 0.42fF
C9754 a_18546_60188# a_28110_60146# 0.35fF
C9755 pmat.rowon_n[4] ctopp 1.57fF
C9756 a_13357_37429# a_10873_36341# 0.80fF
C9757 a_10515_61839# a_9963_13967# 1.88fF
C9758 pmat.rowoff_n[7] nmat.rowoff_n[8] 20.45fF
C9759 a_35230_23548# vcm 0.65fF
C9760 a_26194_69182# ctopp 3.58fF
C9761 a_37238_9492# vcm 0.65fF
C9762 VDD a_35230_69182# 0.52fF
C9763 a_13643_29415# nmat.rowon_n[12] 0.32fF
C9764 a_1739_47893# a_1895_20346# 0.34fF
C9765 VDD a_35290_44527# 0.36fF
C9766 pmat.col_n[6] m2_24960_54946# 0.38fF
C9767 a_2124_59067# a_2163_58941# 0.70fF
C9768 a_40250_65166# a_41254_65166# 0.97fF
C9769 a_35230_59142# ctopp 3.58fF
C9770 a_29206_11500# ctopn 3.58fF
C9771 VDD a_14917_23983# 1.66fF
C9772 VDD a_44266_59142# 0.52fF
C9773 pmat.col_n[30] ctopp 2.01fF
C9774 a_47278_21540# a_48282_21540# 0.97fF
C9775 VDD a_27049_35515# 1.40fF
C9776 nmat.en_bit_n[1] a_13091_28327# 0.32fF
C9777 a_11067_27239# a_18243_28327# 2.27fF
C9778 nmat.col[29] ctopn 2.00fF
C9779 a_10985_44220# a_10927_43421# 0.41fF
C9780 a_18546_16518# a_40158_16926# 0.35fF
C9781 a_22153_37179# a_13357_37429# 1.24fF
C9782 nmat.col[31] inn_analog 0.52fF
C9783 a_20170_70186# a_21174_70186# 0.97fF
C9784 a_48282_71190# a_48282_70186# 1.00fF
C9785 VDD a_21174_61150# 0.52fF
C9786 a_14773_38306# a_16981_37462# 0.41fF
C9787 pmat.rowon_n[10] nmat.rowon_n[7] 0.46fF
C9788 cgen.dlycontrol4_in[3] a_1923_31743# 3.50fF
C9789 a_33222_13508# vcm 0.65fF
C9790 ANTENNA__1187__B1.DIODE a_45019_38645# 0.87fF
C9791 VDD a_23741_42567# 1.14fF
C9792 ANTENNA__1190__A1.DIODE _1192_.A2 1.14fF
C9793 pmat.col[23] m2_42028_54946# 0.39fF
C9794 m2_17932_10226# m3_18064_10358# 2.76fF
C9795 m2_49056_7214# m2_50060_7214# 0.96fF
C9796 ANTENNA__1395__B1.DIODE clk_vcm 1.30fF
C9797 a_31214_18528# vcm 0.65fF
C9798 VDD a_4976_16091# 4.55fF
C9799 a_10515_15055# nmat.rowon_n[4] 0.73fF
C9800 nmat.col[15] nmat.col[13] 4.08fF
C9801 a_26891_28327# a_37291_29397# 0.39fF
C9802 a_46274_13508# a_47278_13508# 0.97fF
C9803 a_18546_72236# a_33130_72194# 0.35fF
C9804 VDD m3_47180_72146# 0.42fF
C9805 a_42258_15516# vcm 0.65fF
C9806 VDD a_27198_17524# 0.52fF
C9807 a_22361_41479# a_11389_40443# 0.34fF
C9808 cgen.start_conv_in a_25997_42902# 0.38fF
C9809 a_2263_43719# a_12263_50959# 5.05fF
C9810 ANTENNA__1395__A2.DIODE a_20616_27791# 0.46fF
C9811 ANTENNA__1190__B1.DIODE a_24867_53135# 0.53fF
C9812 a_18546_8486# a_19074_8894# 0.35fF
C9813 a_44266_18528# a_45270_18528# 0.97fF
C9814 VDD a_28202_8488# 0.55fF
C9815 a_18546_21538# a_31122_21946# 0.35fF
C9816 VDD cgen.dlycontrol1_in[4] 6.06fF
C9817 VDD pmat.row_n[15] 18.01fF
C9818 a_31214_62154# a_31214_61150# 1.00fF
C9819 pmat.rowoff_n[12] a_1769_13103# 2.16fF
C9820 m2_51064_7214# vcm 0.34fF
C9821 a_18162_17524# vcm 6.95fF
C9822 a_38242_23548# ctopn 3.40fF
C9823 a_23821_35279# a_11681_35823# 0.40fF
C9824 VDD a_44266_19532# 0.52fF
C9825 a_40250_9492# ctopn 3.57fF
C9826 m2_24960_24282# m3_25092_24414# 2.79fF
C9827 pmat.row_n[0] nmat.sample 0.34fF
C9828 VDD a_9441_20189# 3.80fF
C9829 a_4955_40277# a_6830_44655# 0.70fF
C9830 a_38242_60146# vcm 0.62fF
C9831 VDD a_43262_10496# 0.52fF
C9832 VDD a_15921_38550# 1.73fF
C9833 VDD a_6375_15279# 0.46fF
C9834 a_31214_15516# a_31214_14512# 1.00fF
C9835 VDD a_6830_22895# 1.24fF
C9836 a_6292_65479# a_5403_67655# 0.72fF
C9837 VDD pmat.col[0] 14.07fF
C9838 VDD a_6981_21263# 1.01fF
C9839 a_18546_58180# a_50198_58138# 0.35fF
C9840 VDD a_27340_31055# 0.32fF
C9841 a_33222_69182# a_33222_68178# 1.00fF
C9842 a_5497_62839# a_4843_54826# 0.33fF
C9843 a_18546_10494# a_50198_10902# 0.35fF
C9844 a_41254_21540# a_41254_20536# 1.00fF
C9845 a_40677_48437# a_40949_48437# 0.49fF
C9846 VDD a_23182_12504# 0.52fF
C9847 a_50290_62154# ctopp 3.43fF
C9848 pmat.col_n[28] pmat.col[29] 5.92fF
C9849 nmat.col[2] nmat.col_n[1] 6.73fF
C9850 a_44266_16520# vcm 0.65fF
C9851 pmat.sw ANTENNA__1183__B1.DIODE 0.39fF
C9852 VDD a_6283_31591# 22.48fF
C9853 VDD a_47223_38671# 0.41fF
C9854 a_36234_13508# ctopn 3.58fF
C9855 a_31214_57134# vcm 0.62fF
C9856 VDD a_10651_37683# 0.54fF
C9857 a_30210_71190# vcm 0.60fF
C9858 pmat.row_n[7] pmat.row_n[2] 0.47fF
C9859 a_34226_18528# ctopn 3.58fF
C9860 m2_17932_7214# m3_18064_7346# 2.79fF
C9861 m2_17932_62978# vcm 0.44fF
C9862 a_2935_38279# cgen.dlycontrol4_in[3] 0.41fF
C9863 a_49286_70186# ctopp 3.56fF
C9864 a_45270_15516# ctopn 3.58fF
C9865 VDD a_45270_11500# 0.52fF
C9866 VDD m3_51196_21402# 0.33fF
C9867 nmat.col[3] m2_21948_24282# 0.39fF
C9868 a_4719_30287# a_6283_31591# 0.48fF
C9869 VDD a_12875_16341# 0.65fF
C9870 VDD a_6830_44655# 0.47fF
C9871 cgen.dlycontrol2_in[2] a_10873_38517# 1.07fF
C9872 a_4985_51433# a_1586_50247# 1.51fF
C9873 VDD a_45282_32143# 1.41fF
C9874 a_18546_69224# a_45178_69182# 0.35fF
C9875 a_35230_11500# a_35230_10496# 1.00fF
C9876 VDD a_33765_35877# 1.32fF
C9877 VDD pmat.col_n[23] 5.52fF
C9878 VDD a_5784_52423# 1.79fF
C9879 a_14641_57711# pmat.rowon_n[8] 0.37fF
C9880 a_42258_22544# vcm 0.65fF
C9881 a_40250_61150# a_41254_61150# 0.97fF
C9882 a_40250_68178# ctopp 3.58fF
C9883 nmat.sw a_10873_38517# 2.74fF
C9884 VDD a_49286_68178# 0.52fF
C9885 a_13459_28111# comp_latch 0.32fF
C9886 a_25190_12504# a_25190_11500# 1.00fF
C9887 a_40837_46261# a_18597_31599# 0.53fF
C9888 a_9963_13967# a_4339_27804# 0.42fF
C9889 a_23182_63158# pmat.col[4] 0.31fF
C9890 a_42240_29423# a_41949_30761# 1.26fF
C9891 VDD a_22178_56130# 0.55fF
C9892 a_18546_20534# a_51202_20942# 0.35fF
C9893 a_34226_20536# a_35230_20536# 0.97fF
C9894 a_47278_16520# ctopn 3.58fF
C9895 VDD nmat.col[7] 6.88fF
C9896 pmat.sample_n pmat.row_n[15] 0.83fF
C9897 VDD nmat.col[17] 4.35fF
C9898 a_9528_20407# nmat.rowon_n[2] 1.11fF
C9899 a_8831_24501# a_8305_20871# 1.10fF
C9900 VDD m2_31988_7214# 1.05fF
C9901 ANTENNA__1187__B1.DIODE nmat.sw 5.88fF
C9902 a_18546_62196# a_36142_62154# 0.35fF
C9903 a_47278_67174# a_47278_66170# 1.00fF
C9904 a_18546_66212# a_32126_66170# 0.35fF
C9905 a_33222_9492# a_33222_8488# 1.00fF
C9906 VDD a_4811_22351# 0.33fF
C9907 pmat.rowoff_n[4] a_6467_29415# 0.41fF
C9908 VDD nmat.sample_n 32.44fF
C9909 a_3615_71631# a_12217_66389# 0.55fF
C9910 VDD a_25190_66170# 0.52fF
C9911 a_2791_57703# a_1769_47919# 0.31fF
C9912 pmat.rowoff_n[7] a_2422_29575# 1.04fF
C9913 a_14287_70543# vcm 0.44fF
C9914 a_7415_29397# a_8443_20719# 0.87fF
C9915 a_6829_26703# comp_latch 1.86fF
C9916 a_20170_23548# ctopn 3.28fF
C9917 a_46274_17524# a_47278_17524# 0.97fF
C9918 a_20310_28029# clk_ena 0.46fF
C9919 a_44266_57134# a_45270_57134# 0.97fF
C9920 pmat.rowoff_n[12] pmat.rowoff_n[11] 0.55fF
C9921 a_49286_20536# a_49286_19532# 1.00fF
C9922 a_43262_71190# a_44266_71190# 0.97fF
C9923 pmat.rowoff_n[4] a_13091_52047# 0.89fF
C9924 VDD a_17113_39141# 1.24fF
C9925 a_30210_58138# a_31214_58138# 0.97fF
C9926 pmat.row_n[8] pmat.row_n[3] 2.33fF
C9927 VDD a_11041_39860# 7.36fF
C9928 a_50290_14512# vcm 0.65fF
C9929 a_49286_64162# vcm 0.62fF
C9930 a_47278_8488# a_48282_8488# 0.97fF
C9931 a_18546_55168# ctopp 0.38fF
C9932 VDD a_6743_31061# 0.45fF
C9933 a_5651_66975# a_10883_3303# 0.34fF
C9934 a_6787_47607# a_8907_48437# 0.32fF
C9935 nmat.col[7] nmat.rowoff_n[2] 4.83fF
C9936 m2_17932_61974# m2_17932_60970# 0.99fF
C9937 _1194_.B1 a_16311_28327# 0.61fF
C9938 nmat.en_bit_n[1] _1184_.A2 1.09fF
C9939 a_45270_22544# ctopn 3.57fF
C9940 cgen.dlycontrol4_in[3] a_11497_40719# 4.42fF
C9941 VDD a_50290_18528# 0.54fF
C9942 a_6679_15492# a_6375_15279# 0.48fF
C9943 m2_51064_24282# vcm 0.47fF
C9944 VDD m2_51064_64986# 1.02fF
C9945 VDD a_5639_49007# 0.46fF
C9946 a_30210_61150# a_30210_60146# 1.00fF
C9947 a_38242_19532# a_38242_18528# 1.00fF
C9948 a_18546_70228# a_34134_70186# 0.35fF
C9949 VDD a_23182_67174# 0.52fF
C9950 VDD a_14261_42043# 1.29fF
C9951 _1194_.A2 a_15667_27239# 2.63fF
C9952 a_33222_62154# vcm 0.62fF
C9953 a_18546_17522# a_29114_17930# 0.35fF
C9954 a_18546_64204# a_50198_64162# 0.35fF
C9955 VDD a_83656_2767# 0.64fF
C9956 a_18546_57176# a_25098_57134# 0.35fF
C9957 VDD nmat.col_n[6] 5.51fF
C9958 a_31214_59142# a_31214_58138# 1.00fF
C9959 ANTENNA__1395__B1.DIODE a_9963_28111# 0.56fF
C9960 pmat.col_n[13] pmat.col[14] 6.16fF
C9961 a_18546_15514# a_29114_15922# 0.35fF
C9962 a_23182_15516# a_24186_15516# 0.97fF
C9963 a_10515_13967# a_11948_49783# 0.64fF
C9964 ANTENNA__1195__A1.DIODE a_28915_50959# 0.34fF
C9965 a_48282_60146# ctopp 3.58fF
C9966 m2_48052_72014# m3_48184_72146# 2.79fF
C9967 VDD a_22199_32149# 0.35fF
C9968 a_22178_69182# a_23182_69182# 0.97fF
C9969 VDD pmat.rowon_n[3] 15.44fF
C9970 pmat.row_n[4] a_18162_12504# 25.57fF
C9971 nmat.col_n[11] ctopn 2.02fF
C9972 a_1591_50095# a_1757_50095# 0.66fF
C9973 VDD a_29404_36165# 1.28fF
C9974 a_32218_70186# vcm 0.62fF
C9975 a_18162_11500# vcm 6.95fF
C9976 nmat.en_bit_n[1] a_9411_2215# 0.90fF
C9977 cgen.dlycontrol4_in[1] a_3325_26159# 0.51fF
C9978 pmat.en_bit_n[2] a_28812_29575# 0.69fF
C9979 a_36234_17524# a_36234_16520# 1.00fF
C9980 pmat.row_n[9] a_18546_17522# 0.35fF
C9981 m2_17932_24282# m2_18936_24282# 0.96fF
C9982 a_11927_27399# a_11235_26159# 0.64fF
C9983 a_42258_12504# a_43262_12504# 0.97fF
C9984 a_13432_62581# a_10515_61839# 0.40fF
C9985 cgen.dlycontrol4_in[4] a_1775_35113# 0.40fF
C9986 a_21174_19532# ctopn 3.58fF
C9987 pmat.rowon_n[7] ctopp 1.57fF
C9988 VDD a_39469_43493# 1.34fF
C9989 a_2400_13763# a_2129_12559# 0.67fF
C9990 VDD a_12889_64789# 0.66fF
C9991 a_13459_28111# nmat.col[28] 0.33fF
C9992 VDD m2_17932_19262# 1.01fF
C9993 pmat.col_n[4] _1192_.A2 0.77fF
C9994 a_24374_29941# nmat.col_n[12] 0.76fF
C9995 a_4351_55527# a_5257_69679# 0.39fF
C9996 VDD a_21174_21540# 0.52fF
C9997 a_31214_59142# a_32218_59142# 0.97fF
C9998 a_18546_59184# a_45178_59142# 0.35fF
C9999 ANTENNA__1395__B1.DIODE ANTENNA__1195__A1.DIODE 1.35fF
C10000 a_41254_57134# ctopp 3.57fF
C10001 VDD a_2648_29397# 10.28fF
C10002 a_40250_71190# ctopp 3.40fF
C10003 VDD a_50290_57134# 0.54fF
C10004 a_27198_58138# ctopp 3.58fF
C10005 a_23182_68178# vcm 0.62fF
C10006 VDD comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top 0.93fF
C10007 VDD a_49286_71190# 0.55fF
C10008 ANTENNA__1197__A.DIODE _1183_.A2 16.67fF
C10009 VDD a_36234_58138# 0.52fF
C10010 VDD a_18546_72236# 33.37fF
C10011 a_24186_62154# pmat.col[5] 0.31fF
C10012 a_18546_60188# a_21082_60146# 0.35fF
C10013 _1154_.X a_16311_28327# 0.41fF
C10014 a_15667_27239# a_44444_32233# 0.35fF
C10015 a_7109_29423# a_6981_28879# 0.30fF
C10016 a_2129_10383# config_1_in[2] 0.32fF
C10017 a_13459_28111# a_20475_49783# 0.39fF
C10018 pmat.en_bit_n[2] a_22459_28879# 0.41fF
C10019 a_11067_27239# nmat.col_n[1] 0.46fF
C10020 nmat.col_n[1] nmat.rowoff_n[3] 0.35fF
C10021 VDD a_38935_39913# 0.64fF
C10022 a_27198_68178# a_27198_67174# 1.00fF
C10023 a_28202_23548# vcm 0.65fF
C10024 a_30210_9492# vcm 0.65fF
C10025 a_32687_46607# a_29937_31055# 1.99fF
C10026 VDD a_28202_69182# 0.52fF
C10027 a_18546_22542# a_47186_22950# 0.35fF
C10028 VDD config_1_in[6] 0.97fF
C10029 VDD a_22541_44581# 1.37fF
C10030 nmat.sw a_5179_31591# 0.86fF
C10031 pmat.col_n[2] m2_20944_54946# 0.37fF
C10032 VDD m2_29980_24282# 0.62fF
C10033 a_46274_20536# vcm 0.65fF
C10034 a_12345_39100# a_25755_38695# 0.69fF
C10035 a_28202_59142# ctopp 3.58fF
C10036 a_22178_11500# ctopn 3.58fF
C10037 pmat.row_n[12] pmat.rowoff_n[12] 21.17fF
C10038 VDD a_30412_31751# 0.37fF
C10039 VDD pmat.rowoff_n[2] 2.66fF
C10040 VDD a_37238_59142# 0.52fF
C10041 pmat.col[26] vcm 5.88fF
C10042 cgen.dlycontrol3_in[4] a_10873_36341# 0.43fF
C10043 pmat.sw nmat.col[31] 6.74fF
C10044 _1196_.B1 a_30571_50959# 0.76fF
C10045 a_18546_16518# a_33130_16926# 0.35fF
C10046 a_25190_16520# a_26194_16520# 0.97fF
C10047 ANTENNA__1197__A.DIODE a_34204_27765# 0.38fF
C10048 VDD a_2879_60975# 0.33fF
C10049 a_36234_55126# m2_37008_54946# 0.96fF
C10050 pmat.col_n[25] vcm 2.80fF
C10051 a_4128_64391# a_6559_57167# 0.52fF
C10052 nmat.rowon_n[14] a_2422_29575# 0.92fF
C10053 a_26194_13508# vcm 0.65fF
C10054 m2_42028_7214# m2_43032_7214# 0.96fF
C10055 a_24186_18528# vcm 0.65fF
C10056 a_2411_33749# a_5823_40303# 0.34fF
C10057 ANTENNA_fanout52_A.DIODE vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.45fF
C10058 m2_17932_17254# m2_17932_16250# 0.99fF
C10059 VDD nmat.rowoff_n[5] 2.50fF
C10060 a_30663_50087# a_10883_3303# 0.48fF
C10061 VDD a_9217_23983# 1.47fF
C10062 VDD m3_19068_72146# 0.41fF
C10063 _1196_.B1 ANTENNA__1190__A2.DIODE 1.18fF
C10064 a_35230_15516# vcm 0.65fF
C10065 a_3339_59879# a_5053_59575# 0.79fF
C10066 a_2563_34837# a_2467_35015# 0.36fF
C10067 a_2263_43719# a_12447_16143# 0.57fF
C10068 a_12723_64789# a_12889_64789# 0.69fF
C10069 VDD a_6343_32661# 0.51fF
C10070 a_34226_70186# a_34226_69182# 1.00fF
C10071 VDD a_21174_8488# 0.55fF
C10072 a_4339_27804# a_4516_21531# 1.72fF
C10073 a_12345_36924# a_10873_36341# 0.85fF
C10074 a_4955_40277# a_4705_39759# 0.66fF
C10075 a_18546_21538# a_24094_21946# 0.35fF
C10076 VDD a_12131_71829# 0.30fF
C10077 a_23182_14512# a_23182_13508# 1.00fF
C10078 a_1586_50247# cgen.dlycontrol3_in[1] 0.55fF
C10079 a_31214_23548# ctopn 3.40fF
C10080 a_11067_16359# a_6467_29415# 0.38fF
C10081 VDD a_37238_19532# 0.52fF
C10082 a_4523_21276# a_9441_20189# 0.40fF
C10083 a_33222_9492# ctopn 3.57fF
C10084 VDD m2_49056_72014# 0.98fF
C10085 ANTENNA__1197__A.DIODE ANTENNA__1395__A1.DIODE 1.95fF
C10086 a_27198_57134# a_27198_56130# 1.00fF
C10087 a_13459_28111# a_22307_27791# 0.42fF
C10088 a_31214_19532# a_32218_19532# 0.97fF
C10089 a_31214_60146# vcm 0.62fF
C10090 VDD a_36234_10496# 0.52fF
C10091 a_9411_2215# a_3688_17179# 0.64fF
C10092 ANTENNA__1395__B1.DIODE a_7415_29397# 1.17fF
C10093 pmat.rowon_n[8] pmat.row_n[8] 21.17fF
C10094 a_11067_30287# a_10287_29941# 0.55fF
C10095 a_29937_31055# a_37471_32149# 0.52fF
C10096 a_49286_20536# ctopn 3.57fF
C10097 pmat.row_n[1] a_15899_47939# 2.08fF
C10098 VDD pmat.en_bit_n[2] 11.34fF
C10099 a_18546_58180# a_43170_58138# 0.35fF
C10100 VDD a_3770_57399# 0.36fF
C10101 a_12345_36924# cgen.dlycontrol1_in[3] 2.83fF
C10102 a_30210_10496# a_31214_10496# 0.97fF
C10103 a_18546_10494# a_43170_10902# 0.35fF
C10104 VDD a_1761_11471# 0.31fF
C10105 a_43262_62154# ctopp 3.58fF
C10106 a_19166_13508# a_20170_13508# 0.97fF
C10107 a_37238_16520# vcm 0.65fF
C10108 a_12985_62581# a_12429_62607# 0.50fF
C10109 a_41254_56130# a_42258_56130# 0.97fF
C10110 VDD nmat.rowoff_n[0] 2.05fF
C10111 a_29206_13508# ctopn 3.58fF
C10112 a_24186_57134# vcm 0.62fF
C10113 a_23182_71190# vcm 0.60fF
C10114 a_27198_18528# ctopn 3.58fF
C10115 VDD a_34924_41605# 1.47fF
C10116 a_5081_53135# a_5462_62215# 1.74fF
C10117 a_7840_27247# nmat.col[7] 1.06fF
C10118 a_12079_31061# a_12245_31061# 0.72fF
C10119 VDD a_4705_39759# 1.02fF
C10120 _1194_.A2 a_46386_33231# 1.24fF
C10121 a_42258_70186# ctopp 3.57fF
C10122 a_38242_15516# ctopn 3.58fF
C10123 a_24407_31375# a_41731_49525# 1.15fF
C10124 VDD a_38242_11500# 0.52fF
C10125 a_10641_52815# a_9463_53511# 0.46fF
C10126 a_23182_22544# a_24186_22544# 0.97fF
C10127 a_6283_31591# a_8583_29199# 0.68fF
C10128 VDD a_4745_45519# 0.49fF
C10129 a_46274_62154# a_47278_62154# 0.97fF
C10130 VDD m2_25964_54946# 0.62fF
C10131 a_44266_66170# a_45270_66170# 0.97fF
C10132 VDD dummypin[0] 0.81fF
C10133 a_18546_69224# a_38150_69182# 0.35fF
C10134 VDD a_19166_59142# 0.58fF
C10135 a_11317_36924# cgen.dlycontrol1_in[1] 1.27fF
C10136 VDD a_5363_33551# 12.81fF
C10137 VDD a_13985_35877# 1.33fF
C10138 pmat.col_n[1] pmat.col_n[2] 0.45fF
C10139 a_25839_49783# a_30111_47911# 0.31fF
C10140 a_38851_28327# inn_analog 2.07fF
C10141 VDD a_10391_62911# 0.56fF
C10142 cgen.dlycontrol4_in[5] a_11317_40188# 3.79fF
C10143 a_37238_63158# a_38242_63158# 0.97fF
C10144 VDD m2_17932_67998# 1.01fF
C10145 nmat.col[30] nmat.col_n[24] 10.97fF
C10146 a_25879_31591# nmat.col[15] 0.46fF
C10147 _1154_.A a_25879_31591# 1.06fF
C10148 a_35230_22544# vcm 0.65fF
C10149 VDD a_10513_24135# 0.53fF
C10150 a_33222_68178# ctopp 3.58fF
C10151 a_16311_28327# nmat.col_n[7] 1.03fF
C10152 a_20170_19532# a_20170_18528# 1.00fF
C10153 _1196_.B1 nmat.col_n[1] 1.17fF
C10154 VDD a_42258_68178# 0.52fF
C10155 a_12197_38306# a_13837_37981# 0.33fF
C10156 VDD a_14113_43132# 1.26fF
C10157 a_49286_63158# vcm 0.62fF
C10158 VDD a_4068_25615# 3.72fF
C10159 ANTENNA__1197__A.DIODE ANTENNA__1395__A2.DIODE 0.40fF
C10160 VDD a_28336_29967# 4.82fF
C10161 VDD a_11202_55687# 2.16fF
C10162 a_18546_20534# a_44174_20942# 0.35fF
C10163 a_40250_16520# ctopn 3.58fF
C10164 VDD a_1895_27962# 0.68fF
C10165 VDD m2_17932_7214# 1.38fF
C10166 VDD a_10995_76207# 0.34fF
C10167 a_18546_62196# a_29114_62154# 0.35fF
C10168 VDD a_4128_46983# 2.22fF
C10169 a_18546_66212# a_25098_66170# 0.35fF
C10170 pmat.row_n[8] pmat.row_n[7] 0.44fF
C10171 VDD a_47278_23548# 0.55fF
C10172 a_45270_70186# a_46274_70186# 0.97fF
C10173 VDD a_49286_9492# 0.52fF
C10174 VDD nmat.col[3] 7.71fF
C10175 _1192_.A2 nmat.col[12] 0.63fF
C10176 a_12437_28879# a_16966_29673# 0.75fF
C10177 a_32218_11500# a_33222_11500# 0.97fF
C10178 a_18546_11498# a_47186_11906# 0.35fF
C10179 a_20439_27247# a_12053_27497# 0.59fF
C10180 VDD a_43776_30287# 3.73fF
C10181 a_18546_66212# pmat.rowoff_n[10] 4.09fF
C10182 a_2835_13077# a_12171_18005# 0.35fF
C10183 a_17842_27497# nmat.col_n[3] 0.39fF
C10184 nmat.rowon_n[10] a_18162_13508# 1.33fF
C10185 a_1781_9308# a_2021_11043# 0.69fF
C10186 VDD a_19166_19532# 0.56fF
C10187 nmat.rowon_n[7] pmat.rowoff_n[4] 0.34fF
C10188 a_34226_64162# a_34226_63158# 1.00fF
C10189 nmat.col_n[27] m2_46044_24282# 0.44fF
C10190 a_37238_10496# a_37238_9492# 1.00fF
C10191 a_4128_64391# a_6283_31591# 0.41fF
C10192 a_34226_58138# a_34226_57134# 1.00fF
C10193 VDD a_19283_49783# 2.63fF
C10194 pmat.rowoff_n[4] a_14653_53458# 0.36fF
C10195 a_43262_14512# vcm 0.65fF
C10196 a_42258_64162# vcm 0.62fF
C10197 a_38242_60146# a_38242_59142# 1.00fF
C10198 a_26194_18528# a_26194_17524# 1.00fF
C10199 ANTENNA__1190__A2.DIODE a_2835_13077# 0.56fF
C10200 VDD nmat.col_n[12] 11.92fF
C10201 VDD a_1643_56597# 0.35fF
C10202 a_21279_48999# a_13275_48783# 1.15fF
C10203 VDD a_45270_13508# 0.52fF
C10204 a_38242_22544# ctopn 3.57fF
C10205 VDD a_43262_18528# 0.52fF
C10206 cgen.enable_dlycontrol_in a_21981_34191# 1.75fF
C10207 a_26194_63158# a_26194_62154# 1.00fF
C10208 VDD pmat.col[11] 4.64fF
C10209 a_11067_64015# cgen.enable_dlycontrol_in 0.40fF
C10210 a_42258_67174# a_43262_67174# 0.97fF
C10211 cgen.dlycontrol3_in[1] cgen.start_conv_in 0.69fF
C10212 cgen.dlycontrol3_in[3] a_12197_41570# 1.38fF
C10213 nmat.col_n[26] vcm 3.62fF
C10214 a_5363_70543# a_10409_53903# 0.61fF
C10215 m2_51064_24282# m2_51064_23278# 0.99fF
C10216 a_18546_70228# a_27106_70186# 0.35fF
C10217 nmat.col[21] nmat.col[18] 3.41fF
C10218 a_2715_51969# a_2676_51843# 0.42fF
C10219 a_2411_43301# a_1683_45205# 0.34fF
C10220 a_39246_66170# a_39246_65166# 1.00fF
C10221 a_3305_15823# a_4976_16091# 0.55fF
C10222 a_32218_22544# a_32218_21540# 1.00fF
C10223 VDD a_27519_42359# 0.58fF
C10224 ANTENNA__1197__A.DIODE ANTENNA__1196__A2.DIODE 0.56fF
C10225 VDD a_10791_14191# 0.42fF
C10226 a_31214_14512# a_32218_14512# 0.97fF
C10227 a_18546_14510# a_45178_14918# 0.35fF
C10228 a_26194_62154# vcm 0.62fF
C10229 m2_51064_14242# vcm 0.62fF
C10230 pmat.rowoff_n[4] nmat.rowoff_n[11] 20.25fF
C10231 VDD a_18546_20534# 32.63fF
C10232 a_18546_17522# a_22086_17930# 0.35fF
C10233 a_18546_64204# a_43170_64162# 0.35fF
C10234 a_30210_64162# a_31214_64162# 0.97fF
C10235 a_36234_68178# a_37238_68178# 0.97fF
C10236 VDD a_35559_30209# 0.45fF
C10237 a_14589_40726# a_18975_40871# 0.34fF
C10238 a_10239_77295# a_6795_76989# 0.33fF
C10239 a_20170_15516# ctopn 3.57fF
C10240 a_18243_28327# nmat.sw 5.11fF
C10241 VDD a_20170_11500# 0.52fF
C10242 a_25190_13508# a_25190_12504# 1.00fF
C10243 a_11149_40188# a_11347_40214# 0.31fF
C10244 a_18546_72236# a_36142_72194# 0.35fF
C10245 nmat.col[30] ctopn 2.01fF
C10246 pmat.row_n[11] nmat.rowon_n[14] 4.83fF
C10247 a_18546_15514# a_22086_15922# 0.35fF
C10248 a_45270_65166# vcm 0.62fF
C10249 a_43262_63158# pmat.col[24] 0.31fF
C10250 pmat.row_n[15] a_3305_15823# 0.97fF
C10251 a_41254_60146# ctopp 3.58fF
C10252 a_18546_69224# a_20078_69182# 0.35fF
C10253 VDD a_50290_60146# 0.54fF
C10254 a_13091_52047# a_11067_49871# 1.34fF
C10255 a_8443_20719# a_9395_27791# 0.39fF
C10256 a_2411_43301# a_6007_42479# 0.69fF
C10257 a_3866_57399# a_2419_53351# 0.69fF
C10258 a_25190_70186# vcm 0.62fF
C10259 VDD a_22086_72194# 0.32fF
C10260 a_10055_31591# a_12447_16143# 0.36fF
C10261 m2_29980_24282# m3_30112_24414# 2.79fF
C10262 a_30571_50959# a_45019_38645# 0.89fF
C10263 VDD a_3399_24787# 0.54fF
C10264 a_8305_20871# a_9155_17455# 0.34fF
C10265 a_46274_14512# ctopn 3.58fF
C10266 VDD a_25393_43493# 1.20fF
C10267 VDD a_10575_15253# 0.42fF
C10268 pmat.col_n[12] pmat.col[13] 6.05fF
C10269 a_3339_59879# a_4991_69831# 2.35fF
C10270 a_18546_59184# a_38150_59142# 0.35fF
C10271 a_32218_65166# a_32218_64162# 1.00fF
C10272 pmat.row_n[3] pmat.row_n[0] 0.96fF
C10273 a_34226_57134# ctopp 3.58fF
C10274 a_33222_71190# ctopp 3.40fF
C10275 VDD a_43262_57134# 0.52fF
C10276 a_20170_58138# ctopp 3.57fF
C10277 VDD a_42258_71190# 0.55fF
C10278 VDD a_29206_58138# 0.52fF
C10279 VDD a_5271_71855# 0.41fF
C10280 a_41254_23548# a_42258_23548# 0.97fF
C10281 a_11149_40188# a_11497_40719# 1.40fF
C10282 a_21174_16520# a_21174_15516# 1.00fF
C10283 a_37238_71190# m2_37008_72014# 1.00fF
C10284 VDD a_5383_48783# 0.37fF
C10285 a_43262_9492# a_44266_9492# 0.97fF
C10286 _1192_.B1 ANTENNA__1195__A1.DIODE 0.51fF
C10287 VDD a_6816_60699# 0.62fF
C10288 a_32687_46607# a_35312_31599# 1.52fF
C10289 a_50290_12504# a_50290_11500# 1.00fF
C10290 VDD a_6099_37039# 0.44fF
C10291 ANTENNA__1196__A2.DIODE a_11051_8903# 0.33fF
C10292 m2_22952_7214# m3_23084_7346# 2.79fF
C10293 a_18546_24550# a_43170_24958# 0.35fF
C10294 nmat.col_n[1] a_2835_13077# 0.32fF
C10295 a_9963_28111# a_10441_21263# 0.32fF
C10296 nmat.col_n[31] nmat.col_n[29] 1.11fF
C10297 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col[30] 0.32fF
C10298 pmat.col[1] ctopp 1.92fF
C10299 VDD a_16171_40157# 1.02fF
C10300 VDD a_23700_39655# 1.22fF
C10301 a_21174_23548# vcm 0.65fF
C10302 a_23182_9492# vcm 0.65fF
C10303 VDD a_21174_69182# 0.52fF
C10304 a_1586_50247# a_4259_31375# 0.56fF
C10305 a_45270_61150# vcm 0.62fF
C10306 _1196_.B1 _1194_.A2 2.35fF
C10307 ANTENNA__1190__A1.DIODE a_16311_28327# 2.06fF
C10308 a_18546_22542# a_40158_22950# 0.35fF
C10309 VDD a_1586_8439# 9.33fF
C10310 VDD nmat.col_n[18] 10.81fF
C10311 ANTENNA__1184__B1.DIODE nmat.col[10] 1.80fF
C10312 VDD m2_49056_54946# 0.64fF
C10313 a_39246_20536# vcm 0.65fF
C10314 a_33222_65166# a_34226_65166# 0.97fF
C10315 a_10873_39605# a_14533_39631# 1.71fF
C10316 a_21174_59142# ctopp 3.58fF
C10317 VDD a_2124_31867# 0.63fF
C10318 VDD a_30210_59142# 0.52fF
C10319 a_3746_58487# a_4259_31375# 0.70fF
C10320 a_40250_21540# a_41254_21540# 0.97fF
C10321 VDD pmat.col_n[26] 5.28fF
C10322 a_20170_22544# ctopn 3.56fF
C10323 a_18243_28327# a_22199_30287# 0.58fF
C10324 a_13091_28327# a_28131_50069# 0.34fF
C10325 a_7717_14735# a_8307_23439# 0.39fF
C10326 a_18546_16518# a_26102_16926# 0.35fF
C10327 m2_30984_54946# vcm 0.42fF
C10328 a_11883_62063# a_12217_66389# 0.46fF
C10329 a_41254_71190# a_41254_70186# 1.00fF
C10330 VDD a_2163_67645# 0.52fF
C10331 pmat.col[4] ctopp 1.97fF
C10332 a_18162_13508# vcm 6.95fF
C10333 VDD a_44774_40821# 1.36fF
C10334 ANTENNA__1190__A2.DIODE a_8861_24527# 0.48fF
C10335 a_2411_43301# a_8583_47381# 0.55fF
C10336 m2_35000_7214# m2_36004_7214# 0.96fF
C10337 a_13909_39605# a_11339_39319# 0.69fF
C10338 a_10959_23983# a_11892_21959# 0.72fF
C10339 a_11067_64015# a_2411_33749# 0.65fF
C10340 a_12449_22895# nmat.col[3] 0.39fF
C10341 a_3866_57399# a_2419_69455# 0.46fF
C10342 VDD a_2021_9563# 3.36fF
C10343 a_39246_13508# a_40250_13508# 0.97fF
C10344 a_11892_21959# a_7644_16341# 0.51fF
C10345 a_6283_31591# a_18241_31698# 0.88fF
C10346 a_28202_15516# vcm 0.65fF
C10347 pmat.rowoff_n[12] a_1586_18231# 1.01fF
C10348 VDD a_5266_17143# 1.65fF
C10349 VDD a_13091_50095# 0.76fF
C10350 VDD a_42191_48071# 0.50fF
C10351 a_12815_8213# a_12981_8213# 0.75fF
C10352 VDD a_14005_22589# 0.58fF
C10353 _1183_.A2 nmat.col[19] 0.89fF
C10354 a_10515_15055# nmat.rowon_n[12] 0.41fF
C10355 a_37238_18528# a_38242_18528# 0.97fF
C10356 VDD a_3091_33402# 0.97fF
C10357 a_3615_71631# a_1586_63927# 0.42fF
C10358 a_28202_62154# pmat.col[9] 0.31fF
C10359 a_24186_62154# a_24186_61150# 1.00fF
C10360 a_47278_12504# vcm 0.65fF
C10361 a_19166_14512# a_19166_13508# 1.00fF
C10362 a_20310_28029# a_15753_28879# 0.55fF
C10363 a_24186_23548# ctopn 3.40fF
C10364 VDD a_30210_19532# 0.52fF
C10365 a_26194_9492# ctopn 3.57fF
C10366 m2_40020_54946# m3_40152_55078# 2.79fF
C10367 _1196_.B1 a_44444_32233# 0.86fF
C10368 pmat.row_n[1] pmat.row_n[0] 1.38fF
C10369 VDD m2_35000_72014# 1.36fF
C10370 nmat.rowon_n[7] clk_dig 1.37fF
C10371 a_31675_47695# a_29937_31055# 0.42fF
C10372 a_24186_60146# vcm 0.62fF
C10373 VDD a_29206_10496# 0.52fF
C10374 VDD a_25755_38695# 1.08fF
C10375 nmat.rowon_n[7] a_11067_16359# 1.63fF
C10376 a_10055_31591# a_11435_58791# 0.53fF
C10377 a_42258_20536# ctopn 3.58fF
C10378 VDD a_29627_43983# 0.57fF
C10379 a_48282_15516# a_49286_15516# 0.97fF
C10380 a_24186_15516# a_24186_14512# 1.00fF
C10381 nmat.col[6] vcm 5.76fF
C10382 nmat.sw a_2046_30184# 0.46fF
C10383 a_18546_59184# a_20078_59142# 0.35fF
C10384 a_1858_25615# a_5253_32687# 0.61fF
C10385 pmat.row_n[3] nmat.sample 0.35fF
C10386 a_18546_58180# a_36142_58138# 0.35fF
C10387 a_47278_69182# a_48282_69182# 0.97fF
C10388 a_26194_69182# a_26194_68178# 1.00fF
C10389 VDD a_9577_58229# 0.57fF
C10390 _1154_.A _1179_.X 2.10fF
C10391 a_18546_10494# a_36142_10902# 0.35fF
C10392 _1154_.X a_24407_31375# 3.16fF
C10393 a_34226_21540# a_34226_20536# 1.00fF
C10394 VDD a_26767_34967# 0.57fF
C10395 nmat.col[15] a_33423_47695# 0.83fF
C10396 ANTENNA__1197__B.DIODE a_15667_27239# 0.64fF
C10397 a_36234_62154# ctopp 3.58fF
C10398 VDD a_45270_62154# 0.52fF
C10399 a_30210_16520# vcm 0.65fF
C10400 a_23700_36391# clk_dig 0.32fF
C10401 a_14773_43746# a_12197_43746# 1.59fF
C10402 a_17139_30503# a_28131_50069# 5.13fF
C10403 pmat.row_n[8] a_18546_16518# 0.35fF
C10404 nmat.rowon_n[7] nmat.rowoff_n[13] 0.52fF
C10405 VDD a_2563_34837# 2.13fF
C10406 a_22178_13508# ctopn 3.58fF
C10407 a_5081_53135# a_4985_51433# 4.27fF
C10408 VDD a_23847_40183# 0.65fF
C10409 a_34204_27765# nmat.col[19] 1.21fF
C10410 pmat.en_bit_n[2] a_8583_29199# 0.36fF
C10411 a_1923_69823# a_9135_69679# 0.56fF
C10412 cgen.enable_dlycontrol_in cgen.dlycontrol3_in[0] 1.50fF
C10413 a_35230_70186# ctopp 3.57fF
C10414 VDD a_10497_54697# 0.81fF
C10415 a_3339_59879# a_6787_47607# 1.94fF
C10416 a_18546_67216# vcm 0.40fF
C10417 a_31214_15516# ctopn 3.58fF
C10418 VDD a_44266_70186# 0.52fF
C10419 VDD a_31214_11500# 0.52fF
C10420 a_5363_70543# a_4075_31591# 0.62fF
C10421 pmat.col[16] vcm 5.88fF
C10422 a_45270_23548# a_45270_22544# 1.00fF
C10423 _1194_.B1 a_17842_27497# 0.93fF
C10424 nmat.rowon_n[7] vcm 0.58fF
C10425 VDD a_5713_77295# 0.60fF
C10426 a_44266_60146# a_45270_60146# 0.97fF
C10427 a_50290_12504# ctopn 3.43fF
C10428 a_18546_69224# a_31122_69182# 0.35fF
C10429 a_7779_22583# a_6173_22895# 0.72fF
C10430 nmat.col[16] ctopn 2.03fF
C10431 a_28202_11500# a_28202_10496# 1.00fF
C10432 a_46274_56130# vcm 0.62fF
C10433 a_8491_47911# a_9135_60967# 0.63fF
C10434 a_26891_28327# a_35244_32411# 0.45fF
C10435 a_7415_29397# a_10441_21263# 0.71fF
C10436 a_18563_27791# a_28715_28879# 0.35fF
C10437 config_1_in[15] config_1_in[14] 0.51fF
C10438 a_18546_63200# a_50198_63158# 0.35fF
C10439 a_28202_22544# vcm 0.65fF
C10440 a_33222_61150# a_34226_61150# 0.97fF
C10441 a_26194_68178# ctopp 3.58fF
C10442 ANTENNA__1184__B1.DIODE _1183_.A2 2.13fF
C10443 VDD config_2_in[12] 1.77fF
C10444 a_49286_66170# vcm 0.62fF
C10445 VDD a_35230_68178# 0.52fF
C10446 a_20170_55126# m2_18936_54946# 0.96fF
C10447 VDD nmat.rowoff_n[10] 2.00fF
C10448 nmat.rowon_n[10] nmat.rowoff_n[9] 0.31fF
C10449 a_42258_63158# vcm 0.62fF
C10450 pmat.col_n[31] m2_50060_54946# 0.62fF
C10451 a_14287_31599# a_14453_31599# 0.39fF
C10452 pmat.row_n[6] nmat.rowon_n[9] 21.59fF
C10453 pmat.rowon_n[7] a_4259_31375# 1.24fF
C10454 a_11023_76359# a_10995_76207# 0.34fF
C10455 a_5081_53135# a_3746_58487# 0.42fF
C10456 a_13091_28327# a_42292_47893# 0.41fF
C10457 a_2046_30184# a_1858_25615# 0.66fF
C10458 a_10873_36341# cgen.dlycontrol1_in[3] 0.54fF
C10459 a_27198_20536# a_28202_20536# 0.97fF
C10460 a_18546_20534# a_37146_20942# 0.35fF
C10461 a_33222_16520# ctopn 3.58fF
C10462 VDD result_out[4] 0.74fF
C10463 a_11921_35286# clk_dig 3.75fF
C10464 a_13503_43421# a_15921_38550# 0.37fF
C10465 VDD a_4123_76181# 1.38fF
C10466 a_18546_62196# a_22086_62154# 0.35fF
C10467 a_40250_67174# a_40250_66170# 1.00fF
C10468 a_26194_9492# a_26194_8488# 1.00fF
C10469 VDD a_40250_23548# 0.55fF
C10470 VDD a_1644_65845# 0.31fF
C10471 VDD a_42258_9492# 0.52fF
C10472 a_43533_30761# a_43776_30287# 3.83fF
C10473 a_18546_11498# a_40158_11906# 0.35fF
C10474 VDD a_21999_37737# 0.61fF
C10475 a_11067_64015# nmat.rowoff_n[6] 0.58fF
C10476 nmat.col_n[28] nmat.col[18] 1.80fF
C10477 inp_analog _1192_.A2 0.92fF
C10478 a_38242_56130# m2_38012_54946# 0.99fF
C10479 a_26891_28327# a_28131_50069# 0.30fF
C10480 a_18563_27791# a_25575_31055# 0.82fF
C10481 VDD a_2879_19093# 0.52fF
C10482 a_39246_17524# a_40250_17524# 0.97fF
C10483 pmat.row_n[1] nmat.sample 0.34fF
C10484 a_37238_57134# a_38242_57134# 0.97fF
C10485 a_18546_19530# a_20078_19938# 0.35fF
C10486 a_18162_19532# nmat.rowon_n[4] 1.33fF
C10487 a_10239_14183# comp_latch 0.37fF
C10488 a_42258_20536# a_42258_19532# 1.00fF
C10489 a_47278_67174# vcm 0.62fF
C10490 a_5081_53135# a_1674_57711# 0.53fF
C10491 a_36234_71190# a_37238_71190# 0.97fF
C10492 VDD a_23971_50228# 0.35fF
C10493 a_23182_58138# a_24186_58138# 0.97fF
C10494 VDD a_32256_44869# 0.99fF
C10495 a_17139_30503# a_44763_34293# 0.39fF
C10496 a_36234_14512# vcm 0.65fF
C10497 a_35230_64162# vcm 0.62fF
C10498 VDD m2_39016_24282# 0.62fF
C10499 VDD a_25681_46831# 0.41fF
C10500 a_44266_62154# pmat.col[25] 0.31fF
C10501 a_40250_8488# a_41254_8488# 0.97fF
C10502 VDD nmat.col_n[25] 5.54fF
C10503 ANTENNA_fanout52_A.DIODE a_37820_30485# 0.92fF
C10504 pmat.col_n[0] a_19579_52789# 0.52fF
C10505 VDD a_16381_35286# 1.17fF
C10506 VDD a_38242_13508# 0.52fF
C10507 a_18546_62196# ctopp 1.59fF
C10508 a_48282_14512# a_48282_13508# 1.00fF
C10509 a_9963_13967# nmat.rowon_n[13] 0.46fF
C10510 a_3615_71631# pmat.rowoff_n[4] 1.37fF
C10511 ANTENNA__1197__A.DIODE a_19405_28853# 1.15fF
C10512 a_31214_22544# ctopn 3.57fF
C10513 a_31978_43439# a_11149_40188# 0.37fF
C10514 ANTENNA__1195__A1.DIODE a_30663_50087# 0.65fF
C10515 VDD a_36234_18528# 0.52fF
C10516 m2_20944_24282# vcm 0.42fF
C10517 a_23182_61150# a_23182_60146# 1.00fF
C10518 a_31214_19532# a_31214_18528# 1.00fF
C10519 VDD pmat.row_n[4] 24.55fF
C10520 a_7415_29397# a_5991_23983# 0.43fF
C10521 a_40837_46261# nmat.col_n[26] 0.51fF
C10522 pmat.col_n[28] vcm 2.81fF
C10523 _1179_.X pmat.col[31] 14.36fF
C10524 a_4128_64391# a_5363_33551# 0.61fF
C10525 VDD a_13167_42359# 0.62fF
C10526 VDD a_47278_15516# 0.52fF
C10527 a_18546_14510# a_38150_14918# 0.35fF
C10528 a_10873_38517# clk_dig 1.30fF
C10529 VDD a_2847_20479# 0.37fF
C10530 a_18546_64204# a_36142_64162# 0.35fF
C10531 a_21981_34191# a_25671_40719# 0.35fF
C10532 a_24186_59142# a_24186_58138# 1.00fF
C10533 a_27198_8488# m2_26968_7214# 1.00fF
C10534 nmat.rowon_n[2] ctopn 1.40fF
C10535 a_4075_50087# a_6175_60039# 0.32fF
C10536 a_38242_65166# vcm 0.62fF
C10537 ANTENNA__1395__A1.DIODE ANTENNA__1184__B1.DIODE 6.21fF
C10538 a_45270_21540# vcm 0.65fF
C10539 VDD a_18546_22542# 32.63fF
C10540 a_34226_60146# ctopp 3.58fF
C10541 a_10515_61839# nmat.rowon_n[12] 0.42fF
C10542 VDD a_43262_60146# 0.52fF
C10543 a_12513_36924# a_11057_35836# 3.91fF
C10544 VDD a_5779_71285# 1.68fF
C10545 a_29206_17524# a_29206_16520# 1.00fF
C10546 ANTENNA__1197__A.DIODE ANTENNA__1190__B1.DIODE 1.05fF
C10547 a_18546_19530# a_49194_19938# 0.35fF
C10548 a_39246_14512# ctopn 3.58fF
C10549 a_12263_50959# a_13643_29415# 1.11fF
C10550 ANTENNA__1190__A1.DIODE a_47147_44655# 0.43fF
C10551 a_35230_12504# a_36234_12504# 0.97fF
C10552 _1187_.A2 nmat.col[29] 0.32fF
C10553 a_48282_22544# a_49286_22544# 0.97fF
C10554 VDD a_13837_43421# 1.32fF
C10555 VDD a_49286_16520# 0.52fF
C10556 a_14497_42658# a_11921_41814# 3.33fF
C10557 VDD a_32319_50345# 0.89fF
C10558 a_26891_28327# nmat.col_n[31] 1.20fF
C10559 a_24186_59142# a_25190_59142# 0.97fF
C10560 a_18546_59184# a_31122_59142# 0.35fF
C10561 nmat.col[15] nmat.col[7] 1.06fF
C10562 a_11435_58791# a_6559_33767# 1.51fF
C10563 a_27198_57134# ctopp 3.57fF
C10564 a_26194_71190# ctopp 3.40fF
C10565 VDD a_36234_57134# 0.52fF
C10566 VDD a_35230_71190# 0.55fF
C10567 VDD a_22178_58138# 0.52fF
C10568 VDD a_10751_72917# 0.41fF
C10569 pmat.row_n[12] nmat.col_n[3] 0.61fF
C10570 a_11113_39747# cgen.dlycontrol4_in[2] 1.07fF
C10571 nmat.col_n[15] ctopn 2.04fF
C10572 VDD a_32947_38825# 0.59fF
C10573 nmat.col[5] nmat.col_n[5] 0.75fF
C10574 a_13357_37429# a_12585_37179# 0.83fF
C10575 a_12263_50959# a_16083_50069# 1.05fF
C10576 VDD a_36161_37462# 1.45fF
C10577 a_1781_9308# a_4333_30511# 0.59fF
C10578 VDD a_1591_40853# 0.44fF
C10579 a_18546_55168# a_47186_55126# 0.35fF
C10580 a_18546_24550# a_36142_24958# 0.39fF
C10581 nmat.col_n[30] ANTENNA__1190__A2.DIODE 2.93fF
C10582 VDD a_2283_39189# 0.36fF
C10583 a_20170_68178# a_20170_67174# 1.00fF
C10584 a_20616_27791# clk_ena 0.37fF
C10585 pmat.row_n[3] a_10883_3303# 0.31fF
C10586 a_44444_32233# a_45019_38645# 0.36fF
C10587 a_46274_8488# m2_46044_7214# 1.00fF
C10588 a_38242_61150# vcm 0.62fF
C10589 a_37238_23548# m2_37008_24282# 0.99fF
C10590 a_18546_22542# a_33130_22950# 0.35fF
C10591 a_48282_21540# ctopn 3.58fF
C10592 nmat.rowoff_n[9] vcm 0.30fF
C10593 VDD a_29937_31055# 8.47fF
C10594 a_32218_20536# vcm 0.65fF
C10595 pmat.row_n[8] pmat.rowoff_n[7] 1.15fF
C10596 VDD a_47278_22544# 0.52fF
C10597 a_4081_61127# pmat.rowon_n[0] 0.32fF
C10598 a_5363_70543# a_7899_67477# 0.50fF
C10599 VDD a_7939_7125# 0.52fF
C10600 VDD a_23182_59142# 0.52fF
C10601 a_18546_17522# ctopn 1.59fF
C10602 VDD a_20170_13508# 0.52fF
C10603 VDD a_15655_50613# 0.46fF
C10604 _1192_.B1 a_39939_29967# 0.38fF
C10605 ANTENNA__1197__B.DIODE a_11067_27239# 1.58fF
C10606 ANTENNA__1184__B1.DIODE ANTENNA__1395__A2.DIODE 1.20fF
C10607 a_44266_17524# vcm 0.65fF
C10608 cgen.dlycontrol4_in[5] cgen.dlycontrol4_in[0] 0.39fF
C10609 a_19166_8488# ctopn 3.24fF
C10610 a_5307_67655# a_5595_65301# 0.90fF
C10611 nmat.col_n[2] nmat.col[3] 6.61fF
C10612 a_8439_69653# a_9301_69679# 0.60fF
C10613 a_45270_8488# vcm 0.64fF
C10614 nmat.col[20] m2_39016_24282# 0.39fF
C10615 VDD a_11737_53359# 0.44fF
C10616 cgen.dlycontrol2_in[2] cgen.dlycontrol2_in[1] 1.88fF
C10617 VDD a_11389_40443# 2.51fF
C10618 nmat.col[28] nmat.col_n[24] 5.16fF
C10619 m2_27972_7214# m2_28976_7214# 0.96fF
C10620 ANTENNA__1190__A1.DIODE nmat.col_n[26] 0.60fF
C10621 nmat.sw cgen.dlycontrol1_in[2] 0.82fF
C10622 a_1923_69823# a_7847_73493# 0.35fF
C10623 VDD a_18162_56170# 2.76fF
C10624 VDD a_8439_69653# 1.00fF
C10625 a_4383_7093# a_8703_6202# 0.48fF
C10626 a_6830_22895# a_11892_21959# 0.62fF
C10627 VDD a_3305_27791# 3.82fF
C10628 a_21174_15516# vcm 0.65fF
C10629 a_12228_40693# a_20438_35431# 1.31fF
C10630 a_11041_39860# a_23700_42919# 0.37fF
C10631 VDD a_15667_27239# 14.24fF
C10632 VDD a_10383_75637# 0.42fF
C10633 a_13091_28327# a_34705_51959# 0.36fF
C10634 VDD a_4579_47919# 0.66fF
C10635 a_7109_29423# a_46013_42997# 0.50fF
C10636 pmat.rowoff_n[12] a_2411_43301# 0.37fF
C10637 a_18546_18526# a_50198_18934# 0.35fF
C10638 a_27198_70186# a_27198_69182# 1.00fF
C10639 VDD nmat.rowon_n[15] 3.20fF
C10640 VDD a_1895_36666# 0.53fF
C10641 a_40250_12504# vcm 0.65fF
C10642 a_45270_64162# ctopp 3.58fF
C10643 pmat.row_n[7] nmat.sample 0.35fF
C10644 VDD a_7321_63151# 0.48fF
C10645 a_23821_35279# cgen.dlycontrol1_in[4] 1.01fF
C10646 VDD a_23182_19532# 0.52fF
C10647 a_18162_9492# ctopn 1.49fF
C10648 VDD m2_20944_72014# 0.98fF
C10649 a_20170_57134# a_20170_56130# 1.00fF
C10650 pmat.rowon_n[0] a_1923_31743# 0.77fF
C10651 _1192_.A2 ANTENNA__1395__B1.DIODE 0.33fF
C10652 a_24186_19532# a_25190_19532# 0.97fF
C10653 VDD a_22178_10496# 0.52fF
C10654 a_13091_28327# nmat.col[10] 1.71fF
C10655 a_50290_13508# a_50290_12504# 1.00fF
C10656 a_35230_20536# ctopn 3.58fF
C10657 VDD a_16837_44219# 1.16fF
C10658 VDD nmat.col[2] 4.36fF
C10659 a_18546_58180# a_29114_58138# 0.35fF
C10660 a_23182_10496# a_24186_10496# 0.97fF
C10661 a_18546_10494# a_29114_10902# 0.35fF
C10662 VDD a_18546_57176# 32.63fF
C10663 ANTENNA_fanout52_A.DIODE ANTENNA__1395__A2.DIODE 0.85fF
C10664 ANTENNA__1184__B1.DIODE ANTENNA__1196__A2.DIODE 1.72fF
C10665 a_5411_48695# a_5383_48783# 0.35fF
C10666 a_47278_17524# ctopn 3.58fF
C10667 a_9963_13967# a_4075_31591# 0.39fF
C10668 a_29206_62154# ctopp 3.58fF
C10669 VDD a_38242_62154# 0.52fF
C10670 pmat.rowon_n[11] a_13643_29415# 7.07fF
C10671 a_23182_16520# vcm 0.65fF
C10672 m2_44036_24282# vcm 0.42fF
C10673 a_48282_8488# ctopn 3.40fF
C10674 VDD a_40415_49551# 0.52fF
C10675 a_10515_61839# ANTENNA__1196__A2.DIODE 1.26fF
C10676 a_11067_64015# ANTENNA__1395__B1.DIODE 0.39fF
C10677 a_8111_11209# comp_latch 0.94fF
C10678 a_34226_56130# a_35230_56130# 0.97fF
C10679 a_18546_56172# a_51202_56130# 0.35fF
C10680 a_11202_55687# a_10955_55687# 0.32fF
C10681 a_10055_31591# a_19541_28879# 1.64fF
C10682 nmat.rowon_n[5] vcm 0.86fF
C10683 VDD a_2099_8725# 0.69fF
C10684 cgen.dlycontrol3_in[2] a_20221_40835# 2.31fF
C10685 _1154_.X ANTENNA__1187__B1.DIODE 0.45fF
C10686 nmat.col[10] m2_28976_24282# 0.41fF
C10687 a_48282_65166# ctopp 3.58fF
C10688 VDD a_37923_42359# 0.59fF
C10689 VDD nmat.rowon_n[9] 3.33fF
C10690 ANTENNA__1190__A1.DIODE a_24407_31375# 0.31fF
C10691 a_18546_55168# a_30118_55126# 0.35fF
C10692 a_30278_30511# clk_ena 1.51fF
C10693 a_28202_70186# ctopp 3.57fF
C10694 a_1858_25615# cgen.dlycontrol1_in[2] 1.37fF
C10695 a_1586_18231# a_1757_18005# 0.50fF
C10696 a_18546_71232# a_19074_71190# 0.35fF
C10697 a_24186_15516# ctopn 3.58fF
C10698 VDD a_37238_70186# 0.52fF
C10699 VDD a_24186_11500# 0.52fF
C10700 a_18546_72236# a_39154_72194# 0.35fF
C10701 VDD m3_51196_59094# 0.34fF
C10702 a_6283_31591# a_14453_31599# 0.58fF
C10703 VDD a_21341_28585# 1.13fF
C10704 nmat.en_bit_n[1] a_14917_23983# 0.53fF
C10705 a_46274_16520# a_46274_15516# 1.00fF
C10706 a_39246_62154# a_40250_62154# 0.97fF
C10707 m2_51064_13238# m2_51064_12234# 0.99fF
C10708 a_37238_66170# a_38242_66170# 0.97fF
C10709 pmat.row_n[14] ctopn 1.64fF
C10710 a_19166_62154# m2_17932_61974# 0.96fF
C10711 a_43262_12504# ctopn 3.58fF
C10712 a_18546_69224# a_24094_69182# 0.35fF
C10713 nmat.col[28] ctopn 2.01fF
C10714 a_39246_56130# vcm 0.62fF
C10715 VDD a_23663_36649# 0.62fF
C10716 a_6451_67655# a_5535_57993# 0.37fF
C10717 VDD a_25098_72194# 0.32fF
C10718 pmat.col[3] vcm 5.88fF
C10719 a_2315_44124# a_2389_45859# 0.48fF
C10720 a_30210_63158# a_31214_63158# 0.97fF
C10721 a_18546_63200# a_43170_63158# 0.35fF
C10722 pmat.sw a_20616_27791# 2.15fF
C10723 a_2952_25045# a_5320_27023# 0.66fF
C10724 a_21174_22544# vcm 0.65fF
C10725 VDD a_12075_24847# 0.42fF
C10726 a_34204_27765# nmat.col_n[29] 0.73fF
C10727 a_42258_66170# vcm 0.62fF
C10728 VDD a_28202_68178# 0.52fF
C10729 VDD a_26515_43447# 0.59fF
C10730 VDD a_3063_14741# 0.51fF
C10731 a_35230_63158# vcm 0.62fF
C10732 m2_51064_15246# m3_51196_15378# 2.76fF
C10733 pmat.col_n[27] m2_46044_54946# 0.43fF
C10734 a_18241_31698# nmat.col_n[12] 1.80fF
C10735 VDD a_14943_26703# 1.18fF
C10736 VDD a_49194_55126# 0.44fF
C10737 a_18546_20534# a_30118_20942# 0.35fF
C10738 a_33423_47695# a_43315_48437# 0.96fF
C10739 a_11067_30287# a_15899_47939# 1.03fF
C10740 a_26194_16520# ctopn 3.58fF
C10741 m2_50060_24282# ctopn 0.69fF
C10742 VDD a_21063_48723# 0.40fF
C10743 pmat.rowon_n[5] pmat.rowoff_n[6] 0.89fF
C10744 VDD a_33222_23548# 0.55fF
C10745 a_48282_61150# ctopp 3.58fF
C10746 _1196_.B1 ANTENNA__1197__B.DIODE 1.44fF
C10747 a_38242_70186# a_39246_70186# 0.97fF
C10748 VDD a_35230_9492# 0.52fF
C10749 nmat.col[30] m2_49056_24282# 0.39fF
C10750 a_2411_33749# a_5087_32687# 0.34fF
C10751 VDD a_10878_58487# 1.70fF
C10752 a_25190_11500# a_26194_11500# 0.97fF
C10753 a_18546_11498# a_33130_11906# 0.35fF
C10754 VDD a_39781_41245# 1.40fF
C10755 pmat.sw a_13643_29415# 3.16fF
C10756 a_13459_28111# a_38851_28327# 0.65fF
C10757 m2_27972_7214# m3_28104_7346# 2.79fF
C10758 a_42240_29423# a_41227_29423# 0.34fF
C10759 a_8399_6037# a_8565_6037# 0.72fF
C10760 a_27198_64162# a_27198_63158# 1.00fF
C10761 a_1899_35051# cgen.dlycontrol4_in[5] 0.51fF
C10762 nmat.sample a_9307_31068# 1.24fF
C10763 m2_18936_55950# m3_19068_56082# 2.76fF
C10764 a_2124_67771# a_2163_67645# 0.46fF
C10765 a_30210_10496# a_30210_9492# 1.00fF
C10766 pmat.col[7] m2_25964_54946# 0.40fF
C10767 nmat.col_n[14] nmat.col_n[19] 0.35fF
C10768 a_40250_67174# vcm 0.62fF
C10769 a_18546_71232# a_48190_71190# 0.35fF
C10770 ANTENNA__1395__A1.DIODE nmat.col_n[29] 3.80fF
C10771 a_22567_47381# a_22733_47381# 0.69fF
C10772 _1192_.A2 a_30111_47911# 1.01fF
C10773 a_27198_58138# a_27198_57134# 1.00fF
C10774 a_3325_20175# a_4613_19087# 1.85fF
C10775 VDD config_1_in[13] 1.07fF
C10776 VDD a_12255_44535# 0.59fF
C10777 a_29206_14512# vcm 0.65fF
C10778 pmat.row_n[11] a_3351_27249# 1.76fF
C10779 VDD a_9411_15831# 0.34fF
C10780 a_1586_33927# a_2411_33749# 1.04fF
C10781 _1194_.B1 a_25575_31055# 1.66fF
C10782 a_28202_64162# vcm 0.62fF
C10783 a_31214_60146# a_31214_59142# 1.00fF
C10784 a_18546_11498# ctopn 1.59fF
C10785 a_14287_70543# pmat.row_n[11] 0.44fF
C10786 a_1674_57711# a_1823_66941# 2.07fF
C10787 a_11067_16359# a_2683_22089# 1.55fF
C10788 pmat.row_n[12] vcm 1.21fF
C10789 VDD pmat.col_n[29] 6.64fF
C10790 a_49286_62154# a_49286_61150# 1.00fF
C10791 VDD a_31214_13508# 0.52fF
C10792 a_20439_27247# nmat.col_n[10] 1.54fF
C10793 a_30571_50959# a_47207_35951# 0.31fF
C10794 a_24186_22544# ctopn 3.57fF
C10795 a_13091_28327# _1183_.A2 0.55fF
C10796 VDD a_29206_18528# 0.52fF
C10797 VDD config_2_in[5] 0.83fF
C10798 pmat.sw nmat.en_bit_n[0] 0.36fF
C10799 m2_40020_54946# vcm 0.42fF
C10800 a_35230_67174# a_36234_67174# 0.97fF
C10801 a_11497_38543# a_13597_37571# 0.32fF
C10802 ANTENNA__1183__B1.DIODE nmat.col_n[24] 0.70fF
C10803 a_31701_37462# a_30431_37683# 0.40fF
C10804 a_7068_11703# a_2021_9563# 0.31fF
C10805 a_25190_22544# a_25190_21540# 1.00fF
C10806 a_4075_68583# a_4317_62215# 0.34fF
C10807 a_32218_66170# a_32218_65166# 1.00fF
C10808 VDD a_40250_15516# 0.52fF
C10809 nmat.col[25] nmat.col_n[24] 6.58fF
C10810 a_18546_14510# a_31122_14918# 0.35fF
C10811 a_24186_14512# a_25190_14512# 0.97fF
C10812 a_49286_15516# a_49286_14512# 1.00fF
C10813 pmat.col[5] vcm 5.88fF
C10814 m2_51064_12234# m3_51196_12366# 2.76fF
C10815 ANTENNA__1190__A1.DIODE a_17842_27497# 1.22fF
C10816 a_23182_64162# a_24186_64162# 0.97fF
C10817 a_18546_64204# a_29114_64162# 0.35fF
C10818 a_18546_57176# pmat.rowoff_n[1] 4.09fF
C10819 a_29206_68178# a_30210_68178# 0.97fF
C10820 VDD a_3622_29967# 0.51fF
C10821 a_3305_15823# a_5266_17143# 0.83fF
C10822 VDD a_19166_70186# 0.56fF
C10823 VDD a_5223_11079# 0.44fF
C10824 a_4075_31591# a_1923_31743# 0.59fF
C10825 VDD m2_47048_7214# 1.33fF
C10826 VDD a_10423_16055# 0.57fF
C10827 VDD a_12981_74581# 0.35fF
C10828 a_31214_65166# vcm 0.62fF
C10829 a_38242_21540# vcm 0.65fF
C10830 a_27198_60146# ctopp 3.58fF
C10831 m2_19940_72014# m3_20072_72146# 2.79fF
C10832 VDD a_46386_33231# 1.45fF
C10833 VDD a_4254_7351# 0.32fF
C10834 VDD a_36234_60146# 0.52fF
C10835 a_11921_37462# a_11057_35836# 0.34fF
C10836 a_3351_27249# a_6579_21583# 0.38fF
C10837 VDD a_19891_36919# 0.60fF
C10838 ANTENNA__1197__A.DIODE inn_analog 1.49fF
C10839 a_1923_61759# a_8031_64789# 0.47fF
C10840 a_16478_29423# clk_ena 1.40fF
C10841 m2_17932_58962# vcm 0.44fF
C10842 m2_45040_54946# m3_45172_55078# 2.79fF
C10843 nmat.col[24] nmat.col_n[31] 1.23fF
C10844 a_6664_26159# clk_ena 0.78fF
C10845 a_18546_19530# a_42166_19938# 0.35fF
C10846 m2_28976_54946# m2_29980_54946# 0.96fF
C10847 a_32218_14512# ctopn 3.58fF
C10848 a_13091_28327# a_34204_27765# 0.42fF
C10849 a_18546_12502# a_46182_12910# 0.35fF
C10850 VDD result_out[15] 0.59fF
C10851 VDD cgen.dlycontrol4_in[1] 12.96fF
C10852 VDD a_42258_16520# 0.52fF
C10853 a_18546_59184# a_24094_59142# 0.35fF
C10854 a_25190_65166# a_25190_64162# 1.00fF
C10855 pmat.col[19] m2_38012_54946# 0.39fF
C10856 VDD a_32126_55126# 0.43fF
C10857 a_20170_57134# ctopp 3.56fF
C10858 nmat.en_bit_n[1] nmat.col[7] 0.37fF
C10859 VDD a_9525_58255# 0.39fF
C10860 a_17139_30503# a_37820_30485# 1.52fF
C10861 VDD a_29206_57134# 0.52fF
C10862 a_2879_57487# a_5267_65479# 0.74fF
C10863 a_4976_16091# a_3688_17179# 1.20fF
C10864 VDD a_2847_33749# 0.33fF
C10865 a_45270_69182# vcm 0.62fF
C10866 a_13158_71285# a_13102_71311# 0.78fF
C10867 VDD a_28202_71190# 0.55fF
C10868 a_1717_13647# a_2021_11043# 1.06fF
C10869 a_34226_23548# a_35230_23548# 0.97fF
C10870 a_18546_23546# a_51202_23954# 0.35fF
C10871 ANTENNA__1395__B1.DIODE a_45187_38129# 1.24fF
C10872 pmat.row_n[7] a_10883_3303# 1.43fF
C10873 a_1769_47919# a_1769_14735# 0.53fF
C10874 a_17139_30503# _1183_.A2 3.59fF
C10875 VDD a_44870_48437# 0.60fF
C10876 a_1781_9308# cgen.start_conv_in 0.56fF
C10877 a_36234_9492# a_37238_9492# 0.97fF
C10878 a_10883_3303# a_7415_29397# 1.34fF
C10879 VDD a_11067_27239# 16.04fF
C10880 a_11067_64015# a_15899_47939# 1.24fF
C10881 VDD nmat.rowoff_n[3] 4.17fF
C10882 a_43262_12504# a_43262_11500# 1.00fF
C10883 VDD a_19689_38053# 1.12fF
C10884 VDD a_19166_14512# 0.56fF
C10885 a_21174_56130# m2_20944_54946# 0.99fF
C10886 m2_51064_9222# m3_51196_9354# 2.76fF
C10887 VDD a_18546_64204# 32.64fF
C10888 a_18546_55168# a_40158_55126# 0.35fF
C10889 a_18546_24550# a_29114_24958# 0.35fF
C10890 a_20475_49783# a_21279_48999# 0.44fF
C10891 a_3339_59879# a_10864_68565# 0.44fF
C10892 VDD a_35312_31599# 2.43fF
C10893 a_9305_58229# a_9577_58229# 0.48fF
C10894 ANTENNA__1196__A2.DIODE a_10223_26703# 0.39fF
C10895 a_49286_56130# ctopp 3.39fF
C10896 a_1923_69823# a_3267_74817# 0.34fF
C10897 a_31214_61150# vcm 0.62fF
C10898 ANTENNA__1395__B1.DIODE a_18597_31599# 0.45fF
C10899 a_5257_69679# a_4265_71543# 0.55fF
C10900 nmat.col[0] ctopn 1.55fF
C10901 a_18546_22542# a_26102_22950# 0.35fF
C10902 a_41254_21540# ctopn 3.58fF
C10903 VDD a_1683_45205# 0.48fF
C10904 a_12658_42895# a_11389_40443# 0.46fF
C10905 VDD a_4241_28335# 0.61fF
C10906 VDD m2_18936_54946# 0.66fF
C10907 a_25190_20536# vcm 0.65fF
C10908 a_26194_65166# a_27198_65166# 0.97fF
C10909 VDD a_40250_22544# 0.52fF
C10910 a_2215_47375# a_19541_28879# 0.56fF
C10911 nmat.col[25] ctopn 1.97fF
C10912 a_33222_21540# a_34226_21540# 0.97fF
C10913 VDD a_1591_13103# 0.30fF
C10914 a_45270_63158# ctopp 3.58fF
C10915 VDD a_4025_54965# 3.04fF
C10916 pmat.rowoff_n[8] a_21215_48071# 1.27fF
C10917 a_37238_17524# vcm 0.65fF
C10918 pmat.row_n[4] a_5411_48695# 0.89fF
C10919 m2_50060_24282# m3_50768_24414# 0.80fF
C10920 a_1823_58237# a_1586_50247# 0.43fF
C10921 VDD a_3387_22869# 0.52fF
C10922 m2_25964_24282# m2_26968_24282# 0.96fF
C10923 a_34226_71190# a_34226_70186# 1.00fF
C10924 a_38242_8488# vcm 0.64fF
C10925 a_48282_58138# a_49286_58138# 0.97fF
C10926 a_11711_50959# a_19283_49783# 0.55fF
C10927 VDD a_6007_42479# 0.43fF
C10928 a_4259_73807# a_3838_70455# 0.66fF
C10929 m2_20944_7214# m2_21948_7214# 0.96fF
C10930 VDD a_20695_30485# 0.36fF
C10931 VDD a_5730_54965# 0.87fF
C10932 m2_17932_59966# m2_17932_58962# 0.99fF
C10933 pmat.row_n[4] cgen.dlycontrol4_in[4] 0.37fF
C10934 a_18546_13506# a_47186_13914# 0.35fF
C10935 a_32218_13508# a_33222_13508# 0.97fF
C10936 _1183_.A2 a_11927_27399# 1.37fF
C10937 a_6375_15279# a_6541_15279# 0.50fF
C10938 VDD m2_51064_60970# 1.02fF
C10939 VDD a_43261_48783# 0.40fF
C10940 a_20170_21540# vcm 0.65fF
C10941 a_10955_55687# a_10497_54697# 0.87fF
C10942 a_48282_61150# a_48282_60146# 1.00fF
C10943 a_50290_67174# ctopp 3.43fF
C10944 a_26891_28327# a_37820_30485# 1.55fF
C10945 a_30210_18528# a_31214_18528# 0.97fF
C10946 a_18546_18526# a_43170_18934# 0.35fF
C10947 VDD a_10515_13967# 18.21fF
C10948 a_12345_36924# a_12585_37179# 1.37fF
C10949 a_11921_37462# a_11113_36483# 2.36fF
C10950 VDD a_33341_37692# 1.15fF
C10951 a_13432_62581# a_4075_31591# 0.59fF
C10952 a_33222_12504# vcm 0.65fF
C10953 a_38242_64162# ctopp 3.58fF
C10954 VDD a_48282_14512# 0.52fF
C10955 VDD a_47278_64162# 0.52fF
C10956 a_26891_28327# _1183_.A2 0.47fF
C10957 pmat.sample_n cgen.dlycontrol4_in[1] 0.30fF
C10958 VDD a_7131_19407# 0.39fF
C10959 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top ANTENNA__1183__B1.DIODE 0.51fF
C10960 a_49286_59142# a_49286_58138# 1.00fF
C10961 nmat.rowon_n[1] a_14195_7351# 0.31fF
C10962 ANTENNA__1395__A1.DIODE a_17139_30503# 1.27fF
C10963 a_1674_68047# a_1923_69823# 2.21fF
C10964 a_28202_20536# ctopn 3.58fF
C10965 a_41254_15516# a_42258_15516# 0.97fF
C10966 VDD pmat.col[18] 4.80fF
C10967 pmat.row_n[3] pmat.row_n[1] 14.43fF
C10968 VDD a_11091_26311# 0.93fF
C10969 a_50290_62154# m2_51064_61974# 0.96fF
C10970 a_18546_58180# a_22086_58138# 0.35fF
C10971 a_40250_69182# a_41254_69182# 0.97fF
C10972 a_6835_51183# a_3339_70759# 0.42fF
C10973 cgen.enable_dlycontrol_in a_6467_29415# 3.94fF
C10974 a_18546_10494# a_22086_10902# 0.35fF
C10975 VDD a_8749_57141# 1.23fF
C10976 a_27198_21540# a_27198_20536# 1.00fF
C10977 _1194_.B1 a_18243_28327# 0.92fF
C10978 ANTENNA__1395__A2.DIODE a_13091_28327# 1.32fF
C10979 _1192_.B1 _1192_.A2 1.57fF
C10980 a_33957_48437# a_33685_48437# 0.42fF
C10981 a_33467_46261# a_14887_46377# 0.36fF
C10982 a_40250_17524# ctopn 3.58fF
C10983 a_22178_62154# ctopp 3.58fF
C10984 VDD a_31214_62154# 0.52fF
C10985 a_30155_36893# ndecision_finish 0.58fF
C10986 _1184_.A2 _1183_.A2 3.72fF
C10987 pmat.sw a_6664_26159# 0.55fF
C10988 a_41731_49525# a_44811_36469# 0.44fF
C10989 a_41254_8488# ctopn 3.40fF
C10990 a_18546_56172# a_44174_56130# 0.35fF
C10991 VDD a_43170_24958# 0.44fF
C10992 nmat.col[30] nmat.col[29] 0.40fF
C10993 ANTENNA__1197__A.DIODE clk_ena 1.89fF
C10994 a_16311_28327# nmat.col_n[4] 0.51fF
C10995 pmat.col_n[31] vcm 2.78fF
C10996 a_41254_65166# ctopp 3.58fF
C10997 VDD a_24937_41479# 1.13fF
C10998 VDD a_50290_65166# 0.54fF
C10999 a_18546_55168# a_23090_55126# 0.35fF
C11000 a_49286_59142# a_50290_59142# 0.97fF
C11001 VDD a_30699_29397# 0.70fF
C11002 a_7092_74005# a_7099_74313# 0.91fF
C11003 a_34226_24552# vcm 0.62fF
C11004 a_21174_70186# ctopp 3.57fF
C11005 a_26891_28327# a_34204_27765# 0.37fF
C11006 cgen.dlycontrol2_in[2] a_12345_39100# 5.29fF
C11007 VDD a_30210_70186# 0.52fF
C11008 VDD a_11501_10927# 0.41fF
C11009 nmat.col_n[3] nmat.col_n[1] 0.34fF
C11010 VDD a_7186_25615# 0.57fF
C11011 a_38242_23548# a_38242_22544# 1.00fF
C11012 VDD a_2407_49289# 10.55fF
C11013 ANTENNA__1190__B1.DIODE ANTENNA__1184__B1.DIODE 13.42fF
C11014 ANTENNA__1190__A1.DIODE ANTENNA__1187__B1.DIODE 0.55fF
C11015 VDD a_8583_47381# 0.44fF
C11016 a_18546_8486# a_20078_8894# 0.35fF
C11017 a_37238_60146# a_38242_60146# 0.97fF
C11018 a_36234_12504# ctopn 3.58fF
C11019 a_21174_11500# a_21174_10496# 1.00fF
C11020 a_32218_56130# vcm 0.62fF
C11021 a_31675_47695# a_45019_38645# 3.43fF
C11022 VDD a_11225_35836# 1.00fF
C11023 VDD a_19074_72194# 0.33fF
C11024 a_3345_62839# a_5682_56311# 0.43fF
C11025 VDD _1196_.B1 24.73fF
C11026 a_15101_29423# ANTENNA__1183__B1.DIODE 1.48fF
C11027 a_19166_17524# vcm 0.65fF
C11028 cgen.dlycontrol4_in[5] cgen.dlycontrol4_in[3] 0.40fF
C11029 a_18546_63200# a_36142_63158# 0.35fF
C11030 _1183_.A2 a_9411_2215# 0.82fF
C11031 a_45270_68178# a_45270_67174# 1.00fF
C11032 a_26194_61150# a_27198_61150# 0.97fF
C11033 a_35230_66170# vcm 0.62fF
C11034 a_20170_8488# vcm 0.64fF
C11035 VDD a_21174_68178# 0.52fF
C11036 m2_45040_72014# m2_46044_72014# 0.96fF
C11037 VDD a_17902_43439# 1.18fF
C11038 a_28202_63158# vcm 0.62fF
C11039 pmat.col_n[23] m2_42028_54946# 0.37fF
C11040 a_19166_16520# m2_17932_16250# 0.96fF
C11041 VDD a_14466_28879# 0.33fF
C11042 a_4259_73807# a_2879_57487# 1.20fF
C11043 a_43776_30287# a_37291_29397# 0.40fF
C11044 a_10878_58487# a_10595_53361# 0.37fF
C11045 VDD a_42166_55126# 0.42fF
C11046 pmat.row_n[11] a_13091_52047# 0.93fF
C11047 a_1923_61759# a_1586_63927# 2.51fF
C11048 VDD a_9785_28879# 3.19fF
C11049 ANTENNA__1395__A2.DIODE a_13145_26935# 0.47fF
C11050 a_11057_35836# a_14589_35286# 0.51fF
C11051 a_18546_20534# a_23090_20942# 0.35fF
C11052 a_18162_16520# ctopn 1.49fF
C11053 ANTENNA__1395__A1.DIODE a_26891_28327# 0.33fF
C11054 a_7521_47081# a_6787_47607# 0.32fF
C11055 pmat.row_n[5] a_18162_13508# 25.57fF
C11056 a_2046_30184# clk_dig 0.87fF
C11057 a_10781_42869# a_31095_42367# 0.34fF
C11058 a_43262_16520# a_44266_16520# 0.97fF
C11059 m2_51064_22274# vcm 0.50fF
C11060 a_33222_67174# a_33222_66170# 1.00fF
C11061 VDD a_26194_23548# 0.55fF
C11062 a_41254_61150# ctopp 3.58fF
C11063 a_12309_38659# a_30155_36893# 1.06fF
C11064 VDD a_28202_9492# 0.52fF
C11065 VDD a_50290_61150# 0.54fF
C11066 a_18546_11498# a_26102_11906# 0.35fF
C11067 VDD a_3659_39733# 1.10fF
C11068 VDD a_44266_20536# 0.52fF
C11069 a_32218_17524# a_33222_17524# 0.97fF
C11070 VDD a_15549_39867# 1.48fF
C11071 a_30210_57134# a_31214_57134# 0.97fF
C11072 a_35230_20536# a_35230_19532# 1.00fF
C11073 a_29206_71190# a_30210_71190# 0.97fF
C11074 a_18546_71232# a_41162_71190# 0.35fF
C11075 a_33222_67174# vcm 0.62fF
C11076 a_13459_28111# a_20616_27791# 1.01fF
C11077 ANTENNA_fanout52_A.DIODE ANTENNA__1190__B1.DIODE 0.99fF
C11078 a_42258_62154# pmat.col[23] 0.31fF
C11079 ANTENNA__1184__B1.DIODE a_7109_29423# 0.45fF
C11080 ANTENNA__1395__A1.DIODE _1184_.A2 2.93fF
C11081 _1194_.B1 a_18547_51565# 0.51fF
C11082 pmat.rowoff_n[12] pmat.row_n[6] 0.78fF
C11083 a_18546_65208# pmat.rowoff_n[9] 4.09fF
C11084 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top a_52398_39208# 0.59fF
C11085 a_22178_14512# vcm 0.65fF
C11086 a_21174_64162# vcm 0.62fF
C11087 cgen.dlycontrol2_in[2] a_32072_38567# 0.59fF
C11088 a_33222_8488# a_34226_8488# 0.97fF
C11089 a_18546_8486# a_49194_8894# 0.35fF
C11090 pmat.row_n[1] a_18546_9490# 0.35fF
C11091 a_18546_65208# a_46182_65166# 0.35fF
C11092 nmat.col[1] nmat.col_n[1] 0.66fF
C11093 a_11317_36924# a_11921_35286# 0.38fF
C11094 a_12934_35823# cgen.dlycontrol1_in[1] 0.63fF
C11095 VDD a_24186_13508# 0.52fF
C11096 a_2648_29397# a_3688_17179# 0.32fF
C11097 a_41254_14512# a_41254_13508# 1.00fF
C11098 VDD a_10286_60405# 1.31fF
C11099 VDD a_22178_18528# 0.52fF
C11100 a_3339_59879# a_5651_66975# 0.31fF
C11101 a_9963_13967# a_9441_20189# 0.53fF
C11102 a_18546_67216# a_46182_67174# 0.35fF
C11103 _1192_.A2 a_43720_32143# 0.42fF
C11104 a_45270_57134# a_45270_56130# 1.00fF
C11105 a_24186_19532# a_24186_18528# 1.00fF
C11106 a_49286_19532# a_50290_19532# 0.97fF
C11107 a_18546_59184# vcm 0.40fF
C11108 a_40837_46261# a_42791_32375# 0.38fF
C11109 VDD a_33489_43131# 1.17fF
C11110 a_2007_25597# a_4339_27804# 0.86fF
C11111 VDD a_33222_15516# 0.52fF
C11112 a_18546_14510# a_24094_14918# 0.35fF
C11113 a_18546_7482# a_46182_7890# 0.35fF
C11114 a_18546_64204# a_22086_64162# 0.35fF
C11115 cgen.dlycontrol3_in[4] nmat.rowon_n[14] 0.37fF
C11116 ANTENNA__1196__A2.DIODE a_17139_30503# 0.34fF
C11117 pmat.col_n[15] a_34226_55126# 0.31fF
C11118 pmat.row_n[14] ctopp 1.85fF
C11119 a_48282_10496# a_49286_10496# 0.97fF
C11120 ANTENNA__1395__A2.DIODE a_11927_27399# 0.55fF
C11121 VDD a_10391_69653# 0.39fF
C11122 a_18546_72236# a_18162_72234# 2.62fF
C11123 pmat.sample pmat.row_n[15] 0.42fF
C11124 nmat.col[31] ctopn 2.20fF
C11125 VDD m2_32992_7214# 0.91fF
C11126 ANTENNA__1197__B.DIODE nmat.sw 0.66fF
C11127 VDD a_4399_51157# 3.03fF
C11128 _1183_.A2 nmat.col[13] 0.75fF
C11129 a_25879_31591# nmat.col_n[31] 0.87fF
C11130 a_48282_62154# pmat.col[29] 0.31fF
C11131 a_24186_65166# vcm 0.62fF
C11132 nmat.col_n[2] nmat.col[2] 0.71fF
C11133 VDD a_20879_47893# 0.47fF
C11134 a_31214_21540# vcm 0.65fF
C11135 pmat.sw ANTENNA__1197__A.DIODE 1.50fF
C11136 a_20170_60146# ctopp 3.57fF
C11137 VDD a_29206_60146# 0.52fF
C11138 _1194_.B1 a_30571_50959# 0.34fF
C11139 a_25879_31591# a_44763_34293# 0.31fF
C11140 a_13641_23439# a_19405_28853# 0.82fF
C11141 a_21739_29415# a_10147_29415# 0.32fF
C11142 a_46274_58138# vcm 0.62fF
C11143 ANTENNA__1190__A2.DIODE vcm 2.34fF
C11144 VDD a_18546_63200# 32.63fF
C11145 a_22178_17524# a_22178_16520# 1.00fF
C11146 nmat.rowon_n[7] pmat.row_n[5] 0.32fF
C11147 pmat.sample pmat.col[0] 0.52fF
C11148 cgen.dlycontrol3_in[3] a_24833_40719# 1.33fF
C11149 a_20895_30199# clk_ena 0.65fF
C11150 a_18546_19530# a_35138_19938# 0.35fF
C11151 m2_21948_54946# m2_22952_54946# 0.96fF
C11152 a_8079_46519# a_8051_46607# 0.38fF
C11153 a_25190_14512# ctopn 3.58fF
C11154 a_13459_28111# nmat.en_bit_n[0] 0.64fF
C11155 a_28202_12504# a_29206_12504# 0.97fF
C11156 a_18546_12502# a_39154_12910# 0.35fF
C11157 a_10873_38517# a_11317_36924# 1.49fF
C11158 pmat.rowoff_n[4] _1194_.A2 0.88fF
C11159 a_41254_22544# a_42258_22544# 0.97fF
C11160 VDD a_10873_39605# 8.09fF
C11161 VDD a_35230_16520# 0.52fF
C11162 nmat.sw a_24374_29941# 0.45fF
C11163 a_18546_19530# vcm 0.40fF
C11164 VDD a_25098_55126# 0.42fF
C11165 VDD a_6909_31061# 0.62fF
C11166 VDD a_45178_7890# 0.33fF
C11167 pmat.col_n[1] a_19579_52789# 0.37fF
C11168 VDD a_22178_57134# 0.52fF
C11169 ANTENNA__1395__A2.DIODE _1184_.A2 6.21fF
C11170 a_3339_70759# a_5682_56311# 1.54fF
C11171 a_38242_69182# vcm 0.62fF
C11172 VDD a_21174_71190# 0.55fF
C11173 a_18546_23546# a_44174_23954# 0.35fF
C11174 _1194_.A2 nmat.col_n[3] 1.06fF
C11175 m2_17932_16250# m2_17932_15246# 0.99fF
C11176 m2_17932_23278# vcm 0.44fF
C11177 a_23182_71190# m2_22952_72014# 1.00fF
C11178 VDD m2_17932_63982# 1.11fF
C11179 a_18546_9490# a_48190_9898# 0.35fF
C11180 VDD a_2835_13077# 12.75fF
C11181 a_18546_13506# ctopn 1.59fF
C11182 a_47278_59142# vcm 0.62fF
C11183 VDD a_16505_40157# 1.25fF
C11184 a_21981_34191# a_12345_36924# 1.33fF
C11185 VDD a_15383_42089# 0.64fF
C11186 VDD a_4075_13653# 0.46fF
C11187 VDD a_6568_59887# 0.91fF
C11188 a_18546_24550# a_22086_24958# 0.35fF
C11189 a_6743_31061# a_7047_31226# 0.39fF
C11190 a_31339_31787# a_13641_23439# 0.49fF
C11191 pmat.row_n[5] nmat.rowoff_n[11] 0.62fF
C11192 a_42258_56130# ctopp 3.40fF
C11193 a_20221_40835# a_20605_40719# 0.30fF
C11194 a_24186_61150# vcm 0.62fF
C11195 a_18546_72236# a_42166_72194# 0.35fF
C11196 a_34226_21540# ctopn 3.58fF
C11197 a_19166_70186# m2_17932_70006# 0.96fF
C11198 a_16311_28327# a_28915_50959# 0.52fF
C11199 ANTENNA__1196__A2.DIODE a_26891_28327# 0.57fF
C11200 _1192_.A2 a_30663_50087# 0.45fF
C11201 VDD a_33222_22544# 0.52fF
C11202 a_45270_66170# ctopp 3.58fF
C11203 a_10515_15055# a_12263_50959# 0.33fF
C11204 pmat.col_n[2] ctopp 2.02fF
C11205 VDD a_32035_36649# 0.67fF
C11206 VDD a_28110_72194# 0.32fF
C11207 a_5639_49007# a_5805_49007# 0.69fF
C11208 nmat.rowon_n[7] a_1957_43567# 0.48fF
C11209 a_19166_11500# vcm 0.65fF
C11210 a_38242_63158# ctopp 3.58fF
C11211 ANTENNA__1395__A2.DIODE a_9411_2215# 1.96fF
C11212 a_2199_13887# a_8695_12801# 0.33fF
C11213 VDD a_47278_63158# 0.52fF
C11214 a_30210_17524# vcm 0.65fF
C11215 a_2263_43719# a_21279_48999# 0.30fF
C11216 a_5687_38279# a_5659_38127# 0.38fF
C11217 m2_41024_24282# m3_41156_24414# 2.79fF
C11218 pmat.row_n[2] a_13091_52047# 0.35fF
C11219 _1154_.X a_30571_50959# 0.31fF
C11220 a_18546_61192# a_46182_61150# 0.35fF
C11221 ANTENNA__1197__B.DIODE a_22199_30287# 0.39fF
C11222 a_31214_8488# vcm 0.64fF
C11223 a_7840_27247# a_11091_26311# 0.83fF
C11224 VDD dummypin[13] 1.11fF
C11225 a_9135_60967# a_2411_33749# 0.69fF
C11226 VDD a_35715_43447# 0.62fF
C11227 ANTENNA__1195__A1.DIODE nmat.col[21] 0.98fF
C11228 _1194_.A2 a_41731_49525# 0.43fF
C11229 a_47278_19532# vcm 0.65fF
C11230 ANTENNA__1395__B1.DIODE a_16311_28327# 3.32fF
C11231 ANTENNA__1196__A2.DIODE _1184_.A2 1.60fF
C11232 a_44266_18528# a_44266_17524# 1.00fF
C11233 m2_51064_71010# vcm 0.50fF
C11234 nmat.col_n[1] vcm 2.79fF
C11235 a_46274_10496# vcm 0.65fF
C11236 a_18546_13506# a_40158_13914# 0.35fF
C11237 a_20170_23548# a_20170_22544# 1.00fF
C11238 a_44266_63158# a_44266_62154# 1.00fF
C11239 a_42258_71190# m2_42028_72014# 1.00fF
C11240 _1154_.X ANTENNA__1190__A2.DIODE 0.62fF
C11241 pmat.row_n[15] a_18546_23546# 0.35fF
C11242 a_43262_67174# ctopp 3.58fF
C11243 a_18546_18526# a_36142_18934# 0.35fF
C11244 a_20170_70186# a_20170_69182# 1.00fF
C11245 VDD a_12217_66389# 2.43fF
C11246 VDD a_1591_58799# 0.84fF
C11247 VDD a_16981_37462# 1.13fF
C11248 a_50290_22544# a_50290_21540# 1.00fF
C11249 a_25695_28111# nmat.col_n[11] 1.10fF
C11250 a_26194_12504# vcm 0.65fF
C11251 a_31214_64162# ctopp 3.58fF
C11252 a_24407_31375# a_22628_30485# 0.52fF
C11253 VDD a_41254_14512# 0.52fF
C11254 a_49286_14512# a_50290_14512# 0.97fF
C11255 m2_51064_10226# vcm 0.51fF
C11256 m2_32992_7214# m3_33124_7346# 2.79fF
C11257 VDD a_40250_64162# 0.52fF
C11258 a_18546_24550# a_51202_24958# 0.35fF
C11259 VDD a_33084_40743# 1.15fF
C11260 a_48282_64162# a_49286_64162# 0.97fF
C11261 VDD a_45019_38645# 5.30fF
C11262 a_18243_28327# a_40837_46261# 0.33fF
C11263 a_43262_13508# a_43262_12504# 1.00fF
C11264 a_18546_12502# a_21082_12910# 0.35fF
C11265 a_11067_30287# a_5535_29980# 0.57fF
C11266 ANTENNA__1195__A1.DIODE a_45829_35407# 0.79fF
C11267 a_21174_20536# ctopn 3.58fF
C11268 VDD a_20811_44535# 0.60fF
C11269 VDD a_8937_15823# 0.67fF
C11270 _1224_.X nmat.col[29] 0.78fF
C11271 VDD m2_30984_24282# 0.62fF
C11272 VDD a_13091_7655# 10.70fF
C11273 a_22199_32149# a_22365_32149# 0.42fF
C11274 VDD a_31210_31751# 0.77fF
C11275 ANTENNA__1196__A2.DIODE a_9411_2215# 5.04fF
C11276 VDD a_51202_72194# 0.39fF
C11277 a_21215_48071# a_21279_48999# 3.49fF
C11278 a_33222_17524# ctopn 3.58fF
C11279 a_48282_11500# vcm 0.65fF
C11280 pmat.row_n[13] nmat.rowon_n[7] 1.48fF
C11281 VDD a_24186_62154# 0.52fF
C11282 _1194_.A2 nmat.rowoff_n[14] 2.39fF
C11283 a_34226_8488# ctopn 3.40fF
C11284 a_27198_56130# a_28202_56130# 0.97fF
C11285 a_18546_56172# a_37146_56130# 0.35fF
C11286 VDD a_36142_24958# 0.39fF
C11287 m2_49056_24282# m2_50060_24282# 0.93fF
C11288 a_1586_63927# a_1591_63701# 0.43fF
C11289 a_50290_19532# ctopn 3.43fF
C11290 a_34226_65166# ctopp 3.58fF
C11291 a_7717_14735# a_36459_29673# 0.49fF
C11292 VDD a_6369_39465# 0.95fF
C11293 VDD a_43262_65166# 0.52fF
C11294 a_13091_52047# a_28901_48437# 0.78fF
C11295 a_9963_28111# a_7415_29397# 0.33fF
C11296 VDD a_50290_21540# 0.56fF
C11297 a_4128_64391# a_4025_54965# 2.11fF
C11298 a_50290_65166# a_50290_64162# 1.00fF
C11299 a_49286_10496# ctopn 3.57fF
C11300 VDD a_5967_5461# 0.37fF
C11301 a_18546_68220# a_45178_68178# 0.35fF
C11302 _1179_.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.47fF
C11303 a_5779_71285# a_5497_62839# 0.43fF
C11304 VDD a_23182_70186# 0.52fF
C11305 nmat.col[15] a_29937_31055# 0.98fF
C11306 a_19541_28879# a_13643_29415# 0.58fF
C11307 VDD a_8861_24527# 2.55fF
C11308 pmat.rowoff_n[4] a_18162_12504# 1.33fF
C11309 a_3746_58487# cgen.dlycontrol3_in[2] 0.33fF
C11310 a_32218_62154# a_33222_62154# 0.97fF
C11311 a_39246_16520# a_39246_15516# 1.00fF
C11312 a_30210_66170# a_31214_66170# 0.97fF
C11313 a_1586_63927# a_3175_59585# 0.82fF
C11314 a_18546_60188# a_50198_60146# 0.35fF
C11315 m2_24960_72014# m3_25092_72146# 2.79fF
C11316 a_29206_12504# ctopn 3.58fF
C11317 a_25190_56130# vcm 0.62fF
C11318 VDD a_30489_36893# 1.30fF
C11319 VDD a_13605_71017# 0.55fF
C11320 a_6175_60039# a_4843_54826# 0.89fF
C11321 a_14287_70543# pmat.row_n[8] 1.16fF
C11322 pmat.row_n[5] nmat.rowoff_n[9] 0.43fF
C11323 a_18546_63200# a_29114_63158# 0.35fF
C11324 a_23182_63158# a_24186_63158# 0.97fF
C11325 m2_50060_54946# m3_50192_55078# 0.85fF
C11326 VDD m2_50060_72014# 1.03fF
C11327 a_11927_27399# a_12053_27497# 0.36fF
C11328 pmat.rowon_n[11] a_18162_67214# 1.19fF
C11329 pmat.row_n[11] a_18546_67216# 0.35fF
C11330 a_48282_69182# ctopp 3.58fF
C11331 a_1899_35051# a_2389_45859# 1.94fF
C11332 m2_51064_55950# m2_51064_54946# 0.99fF
C11333 a_28202_66170# vcm 0.62fF
C11334 VDD pmat.rowoff_n[12] 16.09fF
C11335 a_10239_14183# a_6559_33767# 5.18fF
C11336 m2_38012_72014# m2_39016_72014# 0.96fF
C11337 pmat.rowon_n[8] pmat.row_n[7] 0.84fF
C11338 a_14839_66103# pmat.rowon_n[7] 2.24fF
C11339 a_10515_15055# pmat.rowon_n[5] 0.38fF
C11340 a_4128_64391# a_10515_13967# 0.39fF
C11341 a_10781_42364# a_21981_34191# 0.88fF
C11342 a_21174_63158# vcm 0.62fF
C11343 pmat.col_n[19] m2_38012_54946# 0.37fF
C11344 _1224_.X _1187_.A2 1.35fF
C11345 a_2199_13887# a_6487_5629# 0.35fF
C11346 _1196_.B1 a_8583_29199# 0.35fF
C11347 a_15667_27239# nmat.col[15] 6.47fF
C11348 VDD a_12255_34473# 0.61fF
C11349 VDD a_9103_73791# 0.39fF
C11350 VDD dummypin[3] 1.02fF
C11351 a_2263_43719# a_22567_47381# 0.71fF
C11352 a_11113_39747# a_30819_40191# 1.33fF
C11353 a_2215_47375# a_10239_14183# 0.40fF
C11354 a_6283_31591# a_35244_32411# 0.44fF
C11355 a_19166_71190# m2_17932_71010# 0.96fF
C11356 VDD a_18162_23548# 2.77fF
C11357 a_34226_61150# ctopp 3.58fF
C11358 m2_51064_23278# m2_51064_22274# 0.99fF
C11359 a_31214_70186# a_32218_70186# 0.97fF
C11360 a_13091_18535# nmat.rowon_n[14] 1.12fF
C11361 VDD a_21174_9492# 0.52fF
C11362 VDD a_43262_61150# 0.52fF
C11363 nmat.rowon_n[7] nmat.rowon_n[1] 0.34fF
C11364 VDD a_27795_38007# 0.57fF
C11365 a_10055_31591# a_4707_32156# 2.23fF
C11366 VDD a_37739_42089# 0.64fF
C11367 a_4128_64391# a_8749_57141# 0.45fF
C11368 a_10883_3303# a_11067_30287# 0.55fF
C11369 VDD a_37238_20536# 0.52fF
C11370 VDD cgen.dlycontrol2_in[2] 6.91fF
C11371 a_20170_64162# a_20170_63158# 1.00fF
C11372 a_1923_31743# a_6743_31061# 0.34fF
C11373 a_23182_10496# a_23182_9492# 1.00fF
C11374 a_18546_71232# a_34134_71190# 0.35fF
C11375 a_26194_67174# vcm 0.62fF
C11376 a_2935_38279# a_6830_44655# 0.93fF
C11377 a_20170_58138# a_20170_57134# 1.00fF
C11378 a_4383_7093# comp_latch 0.84fF
C11379 ANTENNA__1190__A1.DIODE a_18243_28327# 0.98fF
C11380 a_6451_67655# a_13102_71311# 0.63fF
C11381 VDD a_5921_44629# 0.51fF
C11382 pmat.col_n[30] pmat.col[30] 1.07fF
C11383 VDD a_49286_17524# 0.52fF
C11384 a_11021_43011# a_10781_42364# 0.81fF
C11385 a_10873_39605# a_11113_40835# 0.51fF
C11386 VDD m2_26968_54946# 0.62fF
C11387 a_18546_8486# a_42166_8894# 0.35fF
C11388 a_24186_60146# a_24186_59142# 1.00fF
C11389 a_18546_65208# a_39154_65166# 0.35fF
C11390 VDD nmat.sw 33.51fF
C11391 VDD a_50290_8488# 0.58fF
C11392 a_12069_36341# a_15049_36374# 0.45fF
C11393 a_11067_64015# a_5535_29980# 0.30fF
C11394 _1194_.A2 vcm 1.20fF
C11395 a_42258_62154# a_42258_61150# 1.00fF
C11396 VDD a_8031_13353# 0.47fF
C11397 a_5731_58951# a_5785_48463# 0.55fF
C11398 VDD pmat.col[29] 4.61fF
C11399 VDD a_13427_18303# 0.54fF
C11400 a_11142_64783# a_10921_64786# 0.48fF
C11401 a_28202_67174# a_29206_67174# 0.97fF
C11402 a_18546_67216# a_39154_67174# 0.35fF
C11403 a_18546_56172# a_18162_56170# 2.62fF
C11404 a_25190_66170# a_25190_65166# 1.00fF
C11405 VDD a_15049_42902# 1.31fF
C11406 VDD a_26194_15516# 0.52fF
C11407 a_1823_74557# a_1674_57711# 0.30fF
C11408 a_42258_15516# a_42258_14512# 1.00fF
C11409 ANTENNA__1395__A1.DIODE nmat.col_n[22] 0.42fF
C11410 a_4719_30287# nmat.sw 0.78fF
C11411 VDD a_6579_29199# 0.34fF
C11412 a_18546_7482# a_39154_7890# 0.35fF
C11413 _1194_.A2 _1194_.B1 18.30fF
C11414 a_30571_50959# a_40837_46261# 0.44fF
C11415 a_13641_23439# a_7026_24527# 0.56fF
C11416 pmat.rowon_n[3] a_1923_31743# 0.97fF
C11417 a_44266_69182# a_44266_68178# 1.00fF
C11418 a_22178_68178# a_23182_68178# 0.97fF
C11419 VDD a_45405_30511# 0.34fF
C11420 a_18546_24550# vcm 0.37fF
C11421 a_11057_35836# cgen.dlycontrol1_in[0] 0.43fF
C11422 VDD a_13091_54447# 0.81fF
C11423 a_19166_8488# m2_17932_8218# 0.96fF
C11424 VDD a_45270_12504# 0.52fF
C11425 pmat.col[30] ctopp 1.99fF
C11426 a_5651_66975# a_10049_60663# 2.31fF
C11427 a_4583_68021# pmat.rowoff_n[7] 1.31fF
C11428 VDD m2_18936_7214# 1.27fF
C11429 a_6927_30503# a_6467_29415# 1.10fF
C11430 VDD pmat.col[12] 4.42fF
C11431 nmat.rowon_n[7] a_2659_35015# 2.19fF
C11432 VDD a_4071_47919# 0.39fF
C11433 a_24186_21540# vcm 0.65fF
C11434 VDD pmat.rowon_n[10] 4.02fF
C11435 VDD a_22178_60146# 0.52fF
C11436 a_1591_36501# a_1895_36666# 0.48fF
C11437 a_2021_9563# a_3663_9269# 0.72fF
C11438 VDD a_11149_36924# 4.03fF
C11439 a_2835_13077# a_12337_18005# 0.38fF
C11440 a_39246_58138# vcm 0.62fF
C11441 a_43262_56130# m2_43032_54946# 0.99fF
C11442 cgen.enable_dlycontrol_in a_10873_38517# 0.58fF
C11443 a_50290_15516# m2_51064_15246# 0.96fF
C11444 _1187_.A2 comp_latch 15.49fF
C11445 a_1923_31743# a_2648_29397# 1.08fF
C11446 a_11067_16359# pmat.rowoff_n[9] 0.31fF
C11447 a_18546_19530# a_28110_19938# 0.35fF
C11448 VDD a_18546_10494# 32.63fF
C11449 a_18546_12502# a_32126_12910# 0.35fF
C11450 ANTENNA__1184__B1.DIODE nmat.col_n[10] 4.25fF
C11451 VDD a_12585_39355# 2.52fF
C11452 a_4351_55527# a_5211_57172# 0.43fF
C11453 VDD a_28202_16520# 0.52fF
C11454 a_50290_70186# m2_51064_70006# 0.96fF
C11455 VDD a_31053_47081# 0.40fF
C11456 VDD pmat.col[27] 4.56fF
C11457 a_12237_38772# a_12345_39100# 0.38fF
C11458 VDD a_38150_7890# 0.33fF
C11459 pmat.rowon_n[15] ctopp 1.26fF
C11460 a_46274_11500# a_46274_10496# 1.00fF
C11461 VDD a_2124_56891# 0.39fF
C11462 VDD a_1858_25615# 7.25fF
C11463 a_31214_69182# vcm 0.62fF
C11464 a_25802_48169# a_24602_48169# 0.47fF
C11465 pmat.col_n[4] pmat.col[5] 6.15fF
C11466 a_27198_23548# a_28202_23548# 0.97fF
C11467 a_18546_23546# a_37146_23954# 0.35fF
C11468 _1192_.A2 a_10883_3303# 0.34fF
C11469 a_29206_9492# a_30210_9492# 0.97fF
C11470 a_18546_9490# a_41162_9898# 0.35fF
C11471 nmat.col[23] vcm 5.76fF
C11472 a_3688_17179# a_5266_17143# 0.75fF
C11473 VDD a_13973_66933# 0.84fF
C11474 a_40250_59142# vcm 0.62fF
C11475 VDD a_11339_39319# 4.34fF
C11476 a_36234_12504# a_36234_11500# 1.00fF
C11477 VDD a_22199_30287# 21.22fF
C11478 VDD a_12116_40871# 5.47fF
C11479 a_13091_52047# ANTENNA__1395__B1.DIODE 0.32fF
C11480 ANTENNA__1197__A.DIODE a_13459_28111# 0.64fF
C11481 a_12449_22895# a_8861_24527# 0.34fF
C11482 nmat.col[10] nmat.col_n[9] 6.62fF
C11483 m2_17932_13238# vcm 0.44fF
C11484 pmat.en_bit_n[0] a_20616_27791# 0.36fF
C11485 nmat.col_n[28] nmat.col[21] 5.17fF
C11486 a_2149_45717# a_2347_46070# 0.30fF
C11487 ANTENNA__1195__A1.DIODE nmat.col_n[28] 0.50fF
C11488 VDD a_12999_3855# 0.45fF
C11489 a_35230_56130# ctopp 3.51fF
C11490 VDD a_44266_56130# 0.55fF
C11491 a_45270_20536# a_46274_20536# 0.97fF
C11492 cgen.dlycontrol3_in[2] cgen.dlycontrol3_in[1] 6.67fF
C11493 a_32218_8488# m2_31988_7214# 1.00fF
C11494 a_27198_21540# ctopn 3.58fF
C11495 pmat.rowon_n[3] a_2935_38279# 0.82fF
C11496 _1154_.X _1194_.A2 1.64fF
C11497 a_6292_65479# a_5779_71285# 0.32fF
C11498 a_44266_9492# a_44266_8488# 1.00fF
C11499 VDD a_26194_22544# 0.52fF
C11500 a_38242_66170# ctopp 3.58fF
C11501 VDD a_47278_66170# 0.52fF
C11502 a_26194_21540# a_27198_21540# 0.97fF
C11503 VDD a_16837_36603# 1.18fF
C11504 VDD a_14947_26159# 0.73fF
C11505 nmat.rowon_n[7] pmat.row_n[2] 0.39fF
C11506 a_10515_15055# a_12447_16143# 7.63fF
C11507 a_31214_63158# ctopp 3.58fF
C11508 pmat.rowon_n[3] nmat.rowon_n[4] 2.21fF
C11509 VDD a_40250_63158# 0.52fF
C11510 a_23182_17524# vcm 0.65fF
C11511 a_21174_63158# pmat.col[2] 0.31fF
C11512 a_19166_67174# a_20170_67174# 0.97fF
C11513 a_18546_61192# a_39154_61150# 0.35fF
C11514 VDD a_4337_22351# 1.39fF
C11515 m2_45040_54946# m2_46044_54946# 0.96fF
C11516 a_2791_57703# a_4075_68583# 0.53fF
C11517 a_27198_71190# a_27198_70186# 1.00fF
C11518 a_24186_8488# vcm 0.64fF
C11519 a_19541_28879# a_16478_29423# 1.27fF
C11520 pmat.col_n[8] pmat.col[8] 1.06fF
C11521 a_15667_27239# a_37291_29397# 0.43fF
C11522 pmat.rowon_n[11] a_10515_61839# 3.03fF
C11523 a_41254_58138# a_42258_58138# 0.97fF
C11524 a_1781_9308# a_23933_32143# 0.86fF
C11525 a_25879_31591# _1183_.A2 1.40fF
C11526 ANTENNA_fanout52_A.DIODE clk_ena 0.65fF
C11527 VDD a_8031_64789# 0.49fF
C11528 a_32957_30287# a_31339_31787# 0.58fF
C11529 a_40250_19532# vcm 0.65fF
C11530 a_18546_7482# a_21082_7890# 0.35fF
C11531 a_2263_43719# a_1586_50247# 1.27fF
C11532 a_3615_71631# a_1957_43567# 1.45fF
C11533 a_11113_36483# cgen.dlycontrol1_in[0] 0.49fF
C11534 VDD a_36946_34191# 0.50fF
C11535 ANTENNA__1190__A1.DIODE a_30571_50959# 1.12fF
C11536 a_39246_10496# vcm 0.65fF
C11537 a_25190_13508# a_26194_13508# 0.97fF
C11538 a_18546_13506# a_33130_13914# 0.35fF
C11539 VDD a_5257_69679# 0.70fF
C11540 a_12069_38517# a_10873_38517# 3.12fF
C11541 a_11041_39860# a_11497_40719# 5.02fF
C11542 a_41254_61150# a_41254_60146# 1.00fF
C11543 a_36234_67174# ctopp 3.58fF
C11544 VDD pmat.rowon_n[2] 3.96fF
C11545 a_49286_19532# a_49286_18528# 1.00fF
C11546 a_23182_18528# a_24186_18528# 0.97fF
C11547 a_18546_18526# a_29114_18934# 0.35fF
C11548 VDD a_45270_67174# 0.52fF
C11549 nmat.col_n[3] m2_21948_24282# 0.38fF
C11550 a_14712_37429# a_12585_37179# 0.52fF
C11551 a_18162_12504# vcm 6.95fF
C11552 a_24186_64162# ctopp 3.58fF
C11553 VDD a_26317_40726# 1.08fF
C11554 VDD a_34226_14512# 0.52fF
C11555 VDD a_33222_64162# 0.52fF
C11556 a_34226_55126# a_35230_55126# 0.97fF
C11557 pmat.col[13] clk_ena 0.37fF
C11558 a_18546_17522# a_51202_17930# 0.35fF
C11559 a_4075_50087# a_2389_45859# 0.87fF
C11560 a_18546_57176# a_47186_57134# 0.35fF
C11561 nmat.col[21] nmat.col_n[20] 6.60fF
C11562 a_42258_59142# a_42258_58138# 1.00fF
C11563 a_32687_46607# a_33986_47375# 0.80fF
C11564 pmat.rowon_n[8] a_18546_16518# 4.09fF
C11565 a_42258_23548# m2_42028_24282# 0.99fF
C11566 a_23395_53135# a_16311_28327# 0.65fF
C11567 VDD a_2051_44111# 0.51fF
C11568 VDD a_1757_15829# 0.65fF
C11569 pmat.col_n[27] pmat.col[28] 5.90fF
C11570 VDD nmat.col_n[30] 9.79fF
C11571 a_34226_15516# a_35230_15516# 0.97fF
C11572 a_18546_15514# a_51202_15922# 0.35fF
C11573 VDD m2_50060_54946# 0.51fF
C11574 a_7939_31591# a_2007_25597# 2.98fF
C11575 m2_17932_69002# m3_18064_69134# 2.76fF
C11576 a_33222_69182# a_34226_69182# 0.97fF
C11577 a_26194_17524# ctopn 3.58fF
C11578 a_41254_11500# vcm 0.65fF
C11579 _1154_.A a_11067_27239# 0.46fF
C11580 VDD m2_51064_15246# 1.05fF
C11581 nmat.rowoff_n[0] a_18546_23546# 4.09fF
C11582 a_47278_17524# a_47278_16520# 1.00fF
C11583 m2_31988_54946# vcm 0.42fF
C11584 a_27198_8488# ctopn 3.40fF
C11585 a_20170_9492# a_21174_9492# 0.97fF
C11586 a_18546_56172# a_30118_56130# 0.35fF
C11587 VDD a_29114_24958# 0.44fF
C11588 m2_42028_24282# m2_43032_24282# 0.96fF
C11589 a_12447_16143# cgen.dlycontrol4_in[3] 0.46fF
C11590 a_19166_13508# vcm 0.65fF
C11591 a_43262_19532# ctopn 3.58fF
C11592 a_27198_65166# ctopp 3.58fF
C11593 nmat.col_n[19] nmat.col_n[24] 11.33fF
C11594 nmat.col_n[29] nmat.col[26] 1.74fF
C11595 VDD a_36234_65166# 0.52fF
C11596 a_13091_52047# a_30111_47911# 2.80fF
C11597 a_12228_39605# a_14773_38306# 0.71fF
C11598 VDD a_43262_21540# 0.52fF
C11599 a_42258_59142# a_43262_59142# 0.97fF
C11600 a_5462_62215# a_2215_47375# 0.37fF
C11601 a_12116_39783# a_12235_39913# 0.37fF
C11602 a_42258_10496# ctopn 3.58fF
C11603 a_18546_68220# a_38150_68178# 0.35fF
C11604 a_4705_39759# a_4831_40303# 0.34fF
C11605 a_49286_58138# ctopp 3.57fF
C11606 a_45270_68178# vcm 0.62fF
C11607 a_13275_48783# a_22733_47381# 0.46fF
C11608 a_20170_8488# m2_19940_7214# 1.00fF
C11609 VDD a_7283_11484# 0.57fF
C11610 a_13459_28111# a_45119_32661# 0.41fF
C11611 a_31214_23548# a_31214_22544# 1.00fF
C11612 a_11067_30287# a_7717_14735# 1.80fF
C11613 a_9411_2215# a_31339_31787# 0.88fF
C11614 ANTENNA__1190__B1.DIODE a_9411_2215# 0.36fF
C11615 a_50290_71190# m2_51064_71010# 0.96fF
C11616 a_18546_60188# a_43170_60146# 0.35fF
C11617 a_30210_60146# a_31214_60146# 0.97fF
C11618 a_22178_12504# ctopn 3.58fF
C11619 nmat.sw a_11113_40835# 3.54fF
C11620 ANTENNA__1395__A1.DIODE a_25879_31591# 0.33fF
C11621 VDD a_13443_36919# 0.60fF
C11622 a_18546_63200# a_22086_63158# 0.35fF
C11623 VDD m2_36004_72014# 1.12fF
C11624 a_38242_68178# a_38242_67174# 1.00fF
C11625 pmat.rowoff_n[12] a_4523_21276# 1.47fF
C11626 _1184_.A2 a_7109_29423# 0.36fF
C11627 a_50290_23548# vcm 0.65fF
C11628 a_41254_69182# ctopp 3.58fF
C11629 ANTENNA__1395__B1.DIODE a_24407_31375# 1.11fF
C11630 a_21174_66170# vcm 0.62fF
C11631 VDD a_50290_69182# 0.56fF
C11632 a_38905_28853# nmat.col[29] 0.62fF
C11633 ANTENNA__1197__B.DIODE nmat.col_n[3] 0.60fF
C11634 m2_30984_72014# m2_31988_72014# 0.96fF
C11635 a_14641_57711# nmat.rowon_n[7] 0.45fF
C11636 VDD a_28705_39141# 1.36fF
C11637 a_50290_59142# ctopp 3.43fF
C11638 m2_17932_65990# m3_18064_66122# 2.76fF
C11639 a_44266_11500# ctopn 3.58fF
C11640 VDD a_11877_58261# 0.65fF
C11641 VDD a_25687_34743# 0.63fF
C11642 ANTENNA__1395__A2.DIODE pmat.col[24] 0.35fF
C11643 VDD a_12792_12937# 0.30fF
C11644 pmat.col_n[19] pmat.col[19] 0.75fF
C11645 a_18823_50247# a_19283_49783# 1.29fF
C11646 a_36234_16520# a_37238_16520# 0.97fF
C11647 pmat.col[4] m2_22952_54946# 0.39fF
C11648 a_18162_7484# ctopn 0.30fF
C11649 VDD a_21883_48981# 0.32fF
C11650 a_26194_67174# a_26194_66170# 1.00fF
C11651 a_27198_61150# ctopp 3.58fF
C11652 a_20170_55126# vcm 0.58fF
C11653 pmat.row_n[13] pmat.row_n[12] 9.31fF
C11654 VDD a_36234_61150# 0.52fF
C11655 VDD a_28116_39655# 1.17fF
C11656 ANTENNA__1183__B1.DIODE nmat.col[29] 0.60fF
C11657 pmat.sw ANTENNA_fanout52_A.DIODE 5.63fF
C11658 a_1586_33927# a_4831_34561# 0.83fF
C11659 a_48282_13508# vcm 0.65fF
C11660 VDD a_20572_40517# 1.39fF
C11661 a_1591_26159# a_1757_26159# 0.49fF
C11662 a_46274_18528# vcm 0.65fF
C11663 VDD a_30210_20536# 0.52fF
C11664 a_25190_17524# a_26194_17524# 0.97fF
C11665 a_13718_68591# a_13973_66933# 0.30fF
C11666 a_23182_57134# a_24186_57134# 0.97fF
C11667 a_19166_10496# a_19166_9492# 1.00fF
C11668 a_28202_20536# a_28202_19532# 1.00fF
C11669 a_22178_71190# a_23182_71190# 0.97fF
C11670 a_18546_71232# a_27106_71190# 0.35fF
C11671 a_3339_70759# a_5211_57172# 0.81fF
C11672 a_18546_72236# a_45178_72194# 0.35fF
C11673 VDD a_42258_17524# 0.52fF
C11674 pmat.col_n[16] pmat.col[17] 6.06fF
C11675 a_18546_58180# pmat.rowoff_n[2] 4.09fF
C11676 pmat.rowon_n[2] pmat.rowoff_n[1] 0.41fF
C11677 _1192_.B1 pmat.col[26] 0.48fF
C11678 a_18546_8486# a_35138_8894# 0.35fF
C11679 a_26194_8488# a_27198_8488# 0.97fF
C11680 VDD a_1923_69823# 8.01fF
C11681 a_18546_65208# a_32126_65166# 0.35fF
C11682 a_45270_70186# a_45270_69182# 1.00fF
C11683 VDD a_43262_8488# 0.55fF
C11684 VDD a_2944_59048# 0.47fF
C11685 pmat.col_n[5] ctopp 2.02fF
C11686 a_4068_25615# a_4516_21531# 1.51fF
C11687 nmat.col_n[19] ctopn 2.46fF
C11688 a_18546_21538# a_46182_21946# 0.35fF
C11689 VDD a_31122_72194# 0.33fF
C11690 a_10515_13967# a_11711_50959# 1.12fF
C11691 a_24591_28327# a_37820_30485# 0.36fF
C11692 a_34226_14512# a_34226_13508# 1.00fF
C11693 a_28336_29967# a_41227_29423# 0.39fF
C11694 VDD a_1757_18005# 0.62fF
C11695 m2_46044_24282# m3_46176_24414# 2.79fF
C11696 a_18546_67216# a_32126_67174# 0.35fF
C11697 a_38242_57134# a_38242_56130# 1.00fF
C11698 a_24591_28327# _1183_.A2 1.22fF
C11699 VDD config_2_in[9] 1.42fF
C11700 a_42258_19532# a_43262_19532# 0.97fF
C11701 m2_51064_72014# m2_51064_71010# 0.99fF
C11702 a_18546_55168# a_51202_55126# 0.35fF
C11703 a_7109_29423# a_7939_31591# 2.83fF
C11704 VDD a_18162_15516# 2.74fF
C11705 VDD a_18546_65208# 32.63fF
C11706 a_18546_7482# a_32126_7890# 0.35fF
C11707 pmat.rowoff_n[12] a_1895_23610# 0.36fF
C11708 pmat.rowon_n[9] pmat.rowoff_n[10] 0.59fF
C11709 m2_17932_62978# m3_18064_63110# 2.76fF
C11710 a_18546_68220# a_20078_68178# 0.35fF
C11711 a_18546_69224# pmat.rowoff_n[13] 4.09fF
C11712 pmat.row_n[12] pmat.row_n[11] 0.40fF
C11713 a_41254_10496# a_42258_10496# 0.97fF
C11714 VDD a_3967_56311# 0.42fF
C11715 a_4128_46983# a_2935_38279# 0.55fF
C11716 a_41731_49525# a_31675_47695# 2.43fF
C11717 VDD result_out[2] 0.51fF
C11718 VDD a_38242_12504# 0.52fF
C11719 a_34226_63158# pmat.col[15] 0.31fF
C11720 ANTENNA__1395__A1.DIODE ndecision_finish 5.46fF
C11721 VDD a_28573_48463# 0.48fF
C11722 VDD a_1586_63927# 8.42fF
C11723 VDD a_1769_47919# 4.56fF
C11724 a_43776_30287# a_35244_32411# 0.79fF
C11725 a_46274_57134# vcm 0.62fF
C11726 VDD a_21219_36885# 2.05fF
C11727 a_11067_64015# a_7717_14735# 1.29fF
C11728 a_45270_71190# vcm 0.60fF
C11729 pmat.en_bit_n[0] a_16478_29423# 0.70fF
C11730 a_49286_18528# ctopn 3.57fF
C11731 a_11149_40188# clk_ena 0.96fF
C11732 a_32218_58138# vcm 0.62fF
C11733 m2_38012_7214# m3_38144_7346# 2.79fF
C11734 _1187_.A2 ANTENNA__1183__B1.DIODE 0.70fF
C11735 a_7521_47081# a_5651_66975# 0.44fF
C11736 a_1591_31599# a_1586_50247# 1.10fF
C11737 VDD a_24775_50095# 0.51fF
C11738 a_18546_12502# a_25098_12910# 0.35fF
C11739 a_21174_12504# a_22178_12504# 0.97fF
C11740 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[19] 0.41fF
C11741 VDD m3_51196_7346# 0.46fF
C11742 a_34226_22544# a_35230_22544# 0.97fF
C11743 VDD a_21174_16520# 0.52fF
C11744 a_11927_27399# a_7026_24527# 0.48fF
C11745 _1194_.B1 a_46339_31029# 0.50fF
C11746 a_24591_28327# a_34204_27765# 0.42fF
C11747 m2_51064_11230# m2_51064_10226# 0.99fF
C11748 VDD m2_40020_24282# 0.62fF
C11749 VDD a_26321_46831# 0.62fF
C11750 a_33222_62154# pmat.col[14] 0.31fF
C11751 pmat.row_n[12] a_18546_68220# 0.35fF
C11752 a_14641_57167# pmat.rowoff_n[8] 0.99fF
C11753 VDD a_47039_31599# 0.87fF
C11754 VDD a_31122_7890# 0.34fF
C11755 a_40837_46261# a_44444_32233# 0.82fF
C11756 VDD a_19086_34343# 0.52fF
C11757 a_24186_69182# vcm 0.62fF
C11758 a_37820_30485# a_33423_47695# 2.68fF
C11759 pmat.rowoff_n[12] cgen.dlycontrol4_in[4] 1.09fF
C11760 a_18162_62194# ctopp 1.49fF
C11761 a_18546_23546# a_30118_23954# 0.35fF
C11762 a_28336_29967# a_35520_30083# 0.62fF
C11763 _1179_.X _1183_.A2 0.51fF
C11764 a_48282_63158# a_49286_63158# 0.97fF
C11765 m2_21948_24282# vcm 0.42fF
C11766 a_18546_9490# a_34134_9898# 0.35fF
C11767 a_33222_59142# vcm 0.62fF
C11768 VDD a_18546_61192# 32.63fF
C11769 a_14773_38306# a_14600_37607# 1.05fF
C11770 a_4128_64391# nmat.sw 0.37fF
C11771 VDD a_17113_42405# 1.13fF
C11772 a_2407_49289# a_5497_62839# 0.34fF
C11773 _1224_.X nmat.col[30] 0.31fF
C11774 a_17139_30503# nmat.col[26] 0.65fF
C11775 a_1858_25615# a_8583_29199# 0.35fF
C11776 m2_17932_59966# m3_18064_60098# 2.76fF
C11777 a_28202_56130# ctopp 3.40fF
C11778 VDD a_22871_29967# 0.38fF
C11779 a_4259_73807# a_1899_35051# 0.97fF
C11780 a_1899_35051# a_19541_28879# 0.68fF
C11781 VDD a_37238_56130# 0.55fF
C11782 a_1674_68047# a_5047_76983# 0.66fF
C11783 VDD m3_36136_72146# 0.33fF
C11784 a_4259_73807# a_2419_53351# 0.32fF
C11785 VDD a_4601_74005# 0.67fF
C11786 a_18546_62196# a_51202_62154# 0.35fF
C11787 ANTENNA__1395__A1.DIODE a_24591_28327# 0.88fF
C11788 a_13091_52047# _1192_.B1 0.45fF
C11789 a_19584_52423# a_15667_27239# 0.52fF
C11790 a_18546_66212# a_47186_66170# 0.35fF
C11791 a_31214_66170# ctopp 3.58fF
C11792 cgen.dlycontrol3_in[4] cgen.dlycontrol3_in[3] 1.14fF
C11793 m2_29980_72014# m3_30112_72146# 2.79fF
C11794 VDD a_40250_66170# 0.52fF
C11795 a_43262_11500# a_44266_11500# 0.97fF
C11796 a_1586_18231# a_8305_20871# 0.78fF
C11797 VDD a_47207_35951# 0.66fF
C11798 pmat.rowon_n[14] vcm 0.58fF
C11799 a_24186_63158# ctopp 3.58fF
C11800 a_4351_55527# a_4075_68583# 0.41fF
C11801 VDD a_34942_51701# 1.63fF
C11802 VDD a_33222_63158# 0.52fF
C11803 a_45270_64162# a_45270_63158# 1.00fF
C11804 _1194_.A2 ANTENNA__1190__A1.DIODE 0.87fF
C11805 a_48282_10496# a_48282_9492# 1.00fF
C11806 a_18546_61192# a_32126_61150# 0.35fF
C11807 a_13091_28327# nmat.col_n[10] 0.41fF
C11808 nmat.col[10] nmat.col[7] 0.73fF
C11809 pmat.rowon_n[7] a_12328_48168# 0.50fF
C11810 m2_38012_54946# m2_39016_54946# 0.96fF
C11811 a_32687_46607# a_40837_46261# 0.88fF
C11812 a_45270_58138# a_45270_57134# 1.00fF
C11813 a_10515_61839# a_11435_58791# 3.21fF
C11814 a_33423_47695# a_34204_27765# 0.75fF
C11815 VDD a_12237_38772# 1.89fF
C11816 a_13091_28327# clk_ena 0.30fF
C11817 a_10791_14191# a_10957_14191# 0.69fF
C11818 VDD a_5399_65479# 0.41fF
C11819 nmat.sample_n nmat.col[10] 3.43fF
C11820 a_6787_47607# a_3339_70759# 0.31fF
C11821 a_33222_19532# vcm 0.65fF
C11822 a_49286_60146# a_49286_59142# 1.00fF
C11823 a_37238_18528# a_37238_17524# 1.00fF
C11824 VDD a_18563_27791# 7.82fF
C11825 pmat.row_n[15] pmat.rowon_n[1] 0.88fF
C11826 a_18546_20534# a_18162_20536# 2.61fF
C11827 a_32218_10496# vcm 0.65fF
C11828 VDD a_20170_12504# 0.52fF
C11829 a_18546_13506# a_26102_13914# 0.35fF
C11830 VDD a_11232_73211# 0.66fF
C11831 a_35559_30209# a_35520_30083# 0.46fF
C11832 nmat.col_n[16] ctopn 2.04fF
C11833 a_37238_63158# a_37238_62154# 1.00fF
C11834 a_29206_67174# ctopp 3.58fF
C11835 a_18546_18526# a_22086_18934# 0.35fF
C11836 a_18546_70228# a_49194_70186# 0.35fF
C11837 VDD a_38242_67174# 0.52fF
C11838 nmat.col_n[10] m2_28976_24282# 0.38fF
C11839 a_13597_37571# a_12585_37179# 0.71fF
C11840 cgen.dlycontrol2_in[0] a_11317_36924# 1.23fF
C11841 a_50290_66170# a_50290_65166# 1.00fF
C11842 a_43262_22544# a_43262_21540# 1.00fF
C11843 VDD a_1757_40853# 0.35fF
C11844 pmat.row_n[1] nmat.rowon_n[14] 20.44fF
C11845 VDD a_27198_14512# 0.52fF
C11846 a_4128_64391# a_1858_25615# 0.64fF
C11847 a_26194_56130# m2_25964_54946# 0.99fF
C11848 a_42258_14512# a_43262_14512# 0.97fF
C11849 a_48282_62154# vcm 0.62fF
C11850 VDD a_26194_64162# 0.52fF
C11851 a_7717_14735# a_24747_29967# 0.74fF
C11852 a_20475_49783# a_13275_48783# 0.51fF
C11853 a_18546_17522# a_44174_17930# 0.35fF
C11854 a_41254_64162# a_42258_64162# 0.97fF
C11855 m2_17932_56954# m3_18064_57086# 2.76fF
C11856 a_47278_68178# a_48282_68178# 0.97fF
C11857 a_18546_57176# a_40158_57134# 0.35fF
C11858 pmat.col[24] m2_43032_54946# 0.39fF
C11859 a_13459_28111# nmat.col[19] 0.91fF
C11860 _1179_.X ANTENNA__1395__A1.DIODE 3.58fF
C11861 a_36234_13508# a_36234_12504# 1.00fF
C11862 a_29937_31055# a_46130_34319# 0.74fF
C11863 a_35244_32411# nmat.col_n[18] 0.95fF
C11864 nmat.sw a_3305_15823# 2.44fF
C11865 a_18546_14510# vcm 0.41fF
C11866 a_18546_15514# a_44174_15922# 0.35fF
C11867 pmat.row_n[6] vcm 1.15fF
C11868 pmat.row_n[7] pmat.rowoff_n[7] 21.32fF
C11869 pmat.rowon_n[7] a_10055_31591# 3.23fF
C11870 pmat.row_n[8] nmat.rowon_n[7] 20.11fF
C11871 a_1674_57711# a_5535_57993# 0.42fF
C11872 VDD a_25393_35877# 1.39fF
C11873 pmat.sample pmat.row_n[4] 0.41fF
C11874 a_47278_70186# vcm 0.62fF
C11875 a_11067_64015# pmat.row_n[1] 1.75fF
C11876 a_34226_11500# vcm 0.65fF
C11877 _1192_.B1 nmat.col_n[26] 3.31fF
C11878 ANTENNA__1190__A1.DIODE a_44444_32233# 2.03fF
C11879 VDD a_17163_50857# 0.30fF
C11880 VDD pmat.rowoff_n[4] 12.55fF
C11881 ANTENNA__1197__B.DIODE _1194_.B1 7.94fF
C11882 a_2263_43719# a_38391_48469# 0.32fF
C11883 VDD a_18546_18526# 32.63fF
C11884 pmat.en_bit_n[0] ANTENNA__1197__A.DIODE 3.16fF
C11885 a_20170_56130# a_21174_56130# 0.97fF
C11886 a_18546_56172# a_23090_56130# 0.35fF
C11887 a_14641_57711# pmat.rowoff_n[11] 0.53fF
C11888 pmat.row_n[12] pmat.row_n[2] 0.43fF
C11889 VDD a_22086_24958# 0.44fF
C11890 nmat.col[31] nmat.col[29] 0.82fF
C11891 pmat.row_n[6] _1194_.B1 0.38fF
C11892 a_19233_38215# a_19689_38053# 0.49fF
C11893 pmat.rowoff_n[15] a_14653_53458# 0.35fF
C11894 cgen.dlycontrol4_in[4] a_1858_25615# 1.62fF
C11895 a_36234_19532# ctopn 3.58fF
C11896 a_20170_65166# ctopp 3.57fF
C11897 a_4259_73807# a_2419_69455# 3.34fF
C11898 a_17139_30503# clk_ena 0.82fF
C11899 VDD a_29206_65166# 0.52fF
C11900 VDD nmat.col_n[3] 9.28fF
C11901 VDD a_36234_21540# 0.52fF
C11902 a_43262_65166# a_43262_64162# 1.00fF
C11903 a_35230_10496# ctopn 3.58fF
C11904 a_18546_68220# a_31122_68178# 0.35fF
C11905 VDD a_26899_30761# 0.44fF
C11906 a_42258_58138# ctopp 3.58fF
C11907 a_38242_68178# vcm 0.62fF
C11908 a_36234_24552# m2_37008_24282# 0.96fF
C11909 _1194_.B1 a_31675_47695# 1.79fF
C11910 cgen.dlycontrol4_in[2] a_10949_43124# 2.48fF
C11911 VDD a_9581_73487# 1.90fF
C11912 a_32218_16520# a_32218_15516# 1.00fF
C11913 a_25190_62154# a_26194_62154# 0.97fF
C11914 a_23182_66170# a_24186_66170# 0.97fF
C11915 a_18546_60188# a_36142_60146# 0.35fF
C11916 VDD a_1757_8213# 0.60fF
C11917 a_19166_58138# m2_17932_57958# 0.96fF
C11918 m2_17932_18258# m2_17932_19262# 0.99fF
C11919 a_4865_12533# a_5173_9839# 0.71fF
C11920 VDD a_3784_62607# 0.32fF
C11921 a_3325_20175# a_7693_22365# 0.59fF
C11922 a_19166_9492# ctopn 3.42fF
C11923 VDD m2_21948_72014# 0.99fF
C11924 a_4075_28335# a_4241_28335# 0.69fF
C11925 _1192_.A2 ANTENNA__1195__A1.DIODE 3.24fF
C11926 a_43262_23548# vcm 0.65fF
C11927 a_34226_69182# ctopp 3.58fF
C11928 a_45270_9492# vcm 0.65fF
C11929 VDD a_43262_69182# 0.52fF
C11930 a_2215_47375# a_1586_50247# 0.47fF
C11931 a_50290_23548# m2_51064_23278# 0.96fF
C11932 m2_23956_72014# m2_24960_72014# 0.96fF
C11933 VDD a_17959_44265# 0.62fF
C11934 ANTENNA__1190__A1.DIODE a_32687_46607# 0.77fF
C11935 VDD a_4403_51701# 0.31fF
C11936 a_44266_65166# a_45270_65166# 0.97fF
C11937 a_43262_59142# ctopp 3.58fF
C11938 a_37238_11500# ctopn 3.58fF
C11939 VDD a_18162_57174# 2.73fF
C11940 _1179_.X ANTENNA__1395__A2.DIODE 2.72fF
C11941 ANTENNA__1187__B1.DIODE ANTENNA__1395__B1.DIODE 5.90fF
C11942 a_11067_27239# a_43315_48437# 0.40fF
C11943 a_13432_62581# a_13091_50095# 0.44fF
C11944 a_10441_21263# a_17702_29967# 0.36fF
C11945 a_18546_16518# a_48190_16926# 0.35fF
C11946 m2_45040_24282# vcm 0.42fF
C11947 VDD a_41731_49525# 11.01fF
C11948 a_11067_64015# ANTENNA__1195__A1.DIODE 0.34fF
C11949 pmat.col[9] ctopp 1.97fF
C11950 VDD a_51202_24958# 0.50fF
C11951 a_20170_61150# ctopp 3.57fF
C11952 a_24186_70186# a_25190_70186# 0.97fF
C11953 _1183_.A2 nmat.sample_n 0.30fF
C11954 VDD a_4865_8181# 1.07fF
C11955 m2_17932_17254# m3_18064_17386# 2.76fF
C11956 VDD a_29206_61150# 0.52fF
C11957 a_6099_37039# a_6265_37039# 0.69fF
C11958 _1154_.X ANTENNA__1197__B.DIODE 0.51fF
C11959 a_41254_13508# vcm 0.65fF
C11960 VDD a_39079_40947# 1.93fF
C11961 VDD nmat.rowon_n[10] 3.00fF
C11962 VDD a_2847_63999# 0.39fF
C11963 a_20616_27791# a_15101_29423# 0.37fF
C11964 a_39246_18528# vcm 0.65fF
C11965 VDD a_23182_20536# 0.52fF
C11966 a_6292_65479# a_2407_49289# 1.02fF
C11967 VDD a_39496_30199# 0.57fF
C11968 a_5651_66975# a_9135_60967# 1.71fF
C11969 m2_17932_57958# m2_17932_56954# 0.99fF
C11970 VDD a_1643_52789# 0.35fF
C11971 a_6283_31591# nmat.rowon_n[12] 0.33fF
C11972 a_12969_40175# a_13503_39069# 0.63fF
C11973 a_25190_23548# m2_24960_24282# 0.99fF
C11974 VDD nmat.col[1] 10.10fF
C11975 a_1674_57711# a_2215_47375# 0.88fF
C11976 a_26891_28327# clk_ena 0.42fF
C11977 a_50290_15516# vcm 0.65fF
C11978 VDD a_35230_17524# 0.52fF
C11979 VDD m2_51064_56954# 0.99fF
C11980 a_18546_8486# a_28110_8894# 0.35fF
C11981 a_18546_65208# a_25098_65166# 0.35fF
C11982 a_48282_18528# a_49286_18528# 0.97fF
C11983 VDD a_36234_8488# 0.55fF
C11984 a_14773_37218# a_15049_36374# 0.59fF
C11985 a_17675_37001# a_17996_36391# 0.59fF
C11986 a_18546_21538# a_39154_21946# 0.35fF
C11987 VDD a_26497_36603# 1.39fF
C11988 a_35230_62154# a_35230_61150# 1.00fF
C11989 a_2935_38279# config_2_in[12] 0.43fF
C11990 a_46274_23548# ctopn 3.40fF
C11991 a_1586_8439# a_1591_15829# 0.57fF
C11992 nmat.col[30] nmat.col[28] 1.88fF
C11993 a_48282_9492# ctopn 3.57fF
C11994 nmat.col_n[18] nmat.col_n[31] 3.92fF
C11995 a_18546_67216# a_25098_67174# 0.35fF
C11996 a_21174_67174# a_22178_67174# 0.97fF
C11997 a_46274_60146# vcm 0.62fF
C11998 _1184_.A2 clk_ena 0.45fF
C11999 a_35230_15516# a_35230_14512# 1.00fF
C12000 nmat.rowon_n[13] a_18162_10496# 1.33fF
C12001 a_2124_31867# a_2163_31741# 0.55fF
C12002 a_1781_9308# a_5579_12394# 0.58fF
C12003 a_18546_7482# a_25098_7890# 0.35fF
C12004 VDD nmat.rowoff_n[14] 4.58fF
C12005 _1179_.X ANTENNA__1196__A2.DIODE 4.87fF
C12006 ANTENNA_fanout52_A.DIODE a_13459_28111# 0.41fF
C12007 a_37238_69182# a_37238_68178# 1.00fF
C12008 a_45270_21540# a_45270_20536# 1.00fF
C12009 VDD a_31214_12504# 0.52fF
C12010 a_5687_71829# a_9279_71829# 0.54fF
C12011 a_18546_23546# a_18546_22542# 0.36fF
C12012 a_11337_25071# a_13768_22325# 1.09fF
C12013 a_11067_16359# a_4955_40277# 0.46fF
C12014 cgen.dlycontrol3_in[0] cgen.dlycontrol2_in[3] 0.52fF
C12015 VDD a_22459_48463# 0.56fF
C12016 a_44266_13508# ctopn 3.58fF
C12017 nmat.col[0] m2_18936_24282# 0.39fF
C12018 a_39246_57134# vcm 0.62fF
C12019 a_11067_64015# a_9944_32259# 0.61fF
C12020 a_38242_71190# vcm 0.60fF
C12021 a_1586_33927# cgen.dlycontrol1_in[3] 1.14fF
C12022 a_42258_18528# ctopn 3.58fF
C12023 VDD a_34887_41271# 0.64fF
C12024 a_25190_58138# vcm 0.62fF
C12025 a_1899_35051# a_3069_69367# 0.37fF
C12026 pmat.en_bit_n[0] a_20895_30199# 0.63fF
C12027 a_28704_29568# a_23021_29199# 0.37fF
C12028 a_27763_27221# nmat.col_n[24] 0.60fF
C12029 VDD a_22743_41001# 0.64fF
C12030 nmat.col_n[15] nmat.col[16] 6.77fF
C12031 ANTENNA__1395__A1.DIODE nmat.col[17] 0.31fF
C12032 a_9411_2215# nmat.col_n[10] 1.15fF
C12033 VDD a_11455_50237# 0.43fF
C12034 ANTENNA__1395__A2.DIODE pmat.col[0] 0.99fF
C12035 VDD m3_23084_7346# 0.36fF
C12036 VDD config_1_in[11] 0.89fF
C12037 VDD a_13779_43123# 1.44fF
C12038 a_1957_43567# a_1769_14735# 0.83fF
C12039 a_12789_68021# a_11837_68591# 0.61fF
C12040 VDD a_15543_31573# 0.34fF
C12041 VDD a_24094_7890# 0.33fF
C12042 a_39246_11500# a_39246_10496# 1.00fF
C12043 a_21371_50087# a_19283_49783# 3.14fF
C12044 VDD a_6127_35076# 0.51fF
C12045 a_33957_48437# a_30111_47911# 0.72fF
C12046 _1192_.B1 a_17842_27497# 4.40fF
C12047 a_18546_23546# a_23090_23954# 0.35fF
C12048 VDD clk_dig 9.18fF
C12049 a_19166_63158# a_19166_62154# 1.00fF
C12050 m2_41024_54946# vcm 0.42fF
C12051 a_22178_9492# a_23182_9492# 0.97fF
C12052 a_18546_9490# a_27106_9898# 0.35fF
C12053 a_50290_22544# vcm 0.65fF
C12054 a_44266_61150# a_45270_61150# 0.97fF
C12055 a_48282_68178# ctopp 3.58fF
C12056 VDD a_10975_67503# 0.42fF
C12057 a_26194_59142# vcm 0.62fF
C12058 VDD a_11067_16359# 14.72fF
C12059 ANTENNA__1195__A1.DIODE a_24747_29967# 2.02fF
C12060 a_29206_12504# a_29206_11500# 1.00fF
C12061 pmat.rowoff_n[12] a_11711_50959# 0.87fF
C12062 pmat.row_n[11] a_18546_19530# 0.35fF
C12063 a_21174_56130# ctopp 3.39fF
C12064 a_7658_71543# a_11271_73085# 0.82fF
C12065 a_8477_57141# a_8749_57141# 0.41fF
C12066 VDD a_30210_56130# 0.55fF
C12067 a_38242_20536# a_39246_20536# 0.97fF
C12068 a_2952_25045# a_3325_20175# 0.32fF
C12069 VDD a_5320_27023# 0.62fF
C12070 VDD m2_48052_7214# 1.04fF
C12071 pmat.col[28] ctopp 1.97fF
C12072 VDD nmat.rowoff_n[13] 2.84fF
C12073 a_6787_47607# a_11019_71543# 1.38fF
C12074 a_18546_62196# a_44174_62154# 0.35fF
C12075 a_18546_66212# a_40158_66170# 0.35fF
C12076 a_4243_54991# a_4587_53505# 0.71fF
C12077 a_37238_9492# a_37238_8488# 1.00fF
C12078 a_24186_66170# ctopp 3.58fF
C12079 VDD a_33222_66170# 0.52fF
C12080 a_18546_21538# a_21082_21946# 0.35fF
C12081 a_12851_28853# a_12437_28585# 0.32fF
C12082 VDD a_26194_63158# 0.52fF
C12083 a_6664_26159# a_10147_29415# 2.39fF
C12084 a_48282_57134# a_49286_57134# 0.97fF
C12085 a_18546_61192# a_25098_61150# 0.35fF
C12086 a_16311_28327# a_45861_29967# 0.57fF
C12087 a_47278_71190# a_48282_71190# 0.97fF
C12088 a_20170_71190# a_20170_70186# 1.00fF
C12089 a_14379_6567# a_12079_9615# 15.88fF
C12090 inp_analog a_18243_28327# 0.46fF
C12091 a_36234_55126# pmat.col[17] 0.38fF
C12092 a_2879_57487# a_1674_57711# 0.47fF
C12093 a_1957_43567# a_12559_51325# 0.34fF
C12094 pmat.row_n[5] _1194_.A2 0.32fF
C12095 VDD a_37497_38550# 1.25fF
C12096 VDD vcm 293.69fF
C12097 a_34226_58138# a_35230_58138# 0.97fF
C12098 pmat.rowon_n[3] nmat.rowon_n[12] 21.24fF
C12099 a_26194_19532# vcm 0.65fF
C12100 a_25190_10496# vcm 0.65fF
C12101 a_11337_25071# a_9441_20189# 0.75fF
C12102 a_30603_29575# a_30699_29397# 0.32fF
C12103 a_28202_71190# m2_27972_72014# 1.00fF
C12104 VDD a_45370_48169# 0.65fF
C12105 a_12693_38543# a_13503_36893# 0.60fF
C12106 a_1769_13103# config_2_in[3] 0.52fF
C12107 a_34226_61150# a_34226_60146# 1.00fF
C12108 a_22178_67174# ctopp 3.58fF
C12109 VDD a_14923_38825# 0.64fF
C12110 VDD _1194_.B1 39.97fF
C12111 a_9741_28585# a_9075_28023# 0.64fF
C12112 a_42258_19532# a_42258_18528# 1.00fF
C12113 a_18546_70228# a_42166_70186# 0.35fF
C12114 VDD a_31214_67174# 0.52fF
C12115 VDD a_14833_8945# 0.39fF
C12116 VDD a_39387_40183# 0.61fF
C12117 VDD a_18143_38007# 0.62fF
C12118 VDD a_30913_42043# 1.36fF
C12119 a_41254_62154# vcm 0.62fF
C12120 a_14839_20871# a_14365_22351# 0.69fF
C12121 nmat.col[24] nmat.col[26] 3.79fF
C12122 a_18546_17522# a_37146_17930# 0.35fF
C12123 a_33423_47695# a_44966_43255# 0.48fF
C12124 a_18546_57176# a_33130_57134# 0.35fF
C12125 a_35230_59142# a_35230_58138# 1.00fF
C12126 nmat.rowoff_n[2] vcm 0.31fF
C12127 ANTENNA__1196__A2.DIODE a_45282_32143# 1.18fF
C12128 ANTENNA__1197__B.DIODE a_40837_46261# 0.65fF
C12129 a_18546_72236# a_48190_72194# 0.35fF
C12130 a_27198_15516# a_28202_15516# 0.97fF
C12131 a_18546_15514# a_37146_15922# 0.35fF
C12132 VDD a_33986_47375# 1.22fF
C12133 a_25879_31591# a_7109_29423# 0.73fF
C12134 a_26194_69182# a_27198_69182# 0.97fF
C12135 a_2683_22089# a_3325_20175# 0.55fF
C12136 pmat.col_n[8] ctopp 2.02fF
C12137 nmat.col[27] ctopn 1.97fF
C12138 a_40250_70186# vcm 0.62fF
C12139 VDD a_34134_72194# 0.32fF
C12140 a_27198_11500# vcm 0.65fF
C12141 ANTENNA__1183__B1.DIODE nmat.col[30] 10.82fF
C12142 VDD pmat.col[10] 4.80fF
C12143 VDD a_6583_62607# 0.50fF
C12144 a_34226_24552# a_34226_23548# 1.00fF
C12145 a_2263_43719# a_13275_48783# 0.88fF
C12146 a_40250_17524# a_40250_16520# 1.00fF
C12147 a_4516_21531# a_3305_27791# 0.41fF
C12148 m2_51064_24282# m3_51196_24414# 2.79fF
C12149 _1154_.A a_22199_30287# 0.40fF
C12150 a_31675_47695# a_40837_46261# 0.85fF
C12151 a_10223_26703# a_6829_26703# 1.52fF
C12152 a_46274_12504# a_47278_12504# 0.97fF
C12153 a_42240_29423# inn_analog 0.36fF
C12154 a_29206_19532# ctopn 3.58fF
C12155 pmat.sw a_9411_2215# 0.65fF
C12156 VDD a_22178_65166# 0.52fF
C12157 a_13459_28111# nmat.col_n[29] 1.13fF
C12158 pmat.col_n[21] pmat.col[22] 6.08fF
C12159 VDD a_29206_21540# 0.52fF
C12160 a_35230_59142# a_36234_59142# 0.97fF
C12161 a_28202_10496# ctopn 3.58fF
C12162 a_49286_57134# ctopp 3.56fF
C12163 a_18546_68220# a_24094_68178# 0.35fF
C12164 VDD a_22186_30485# 0.46fF
C12165 a_48282_71190# ctopp 3.40fF
C12166 a_35230_58138# ctopp 3.58fF
C12167 a_31214_68178# vcm 0.62fF
C12168 ANTENNA__1196__A2.DIODE nmat.sample_n 1.42fF
C12169 VDD a_44266_58138# 0.52fF
C12170 pmat.rowoff_n[15] a_3615_71631# 0.31fF
C12171 a_5651_66975# a_10569_64489# 0.31fF
C12172 a_24186_23548# a_24186_22544# 1.00fF
C12173 a_15667_27239# a_35244_32411# 1.61fF
C12174 a_13641_23439# a_9528_20407# 0.63fF
C12175 m2_17932_14242# m2_17932_13238# 0.99fF
C12176 a_47278_71190# m2_47048_72014# 1.00fF
C12177 VDD m2_17932_59966# 1.00fF
C12178 a_23182_60146# a_24186_60146# 0.97fF
C12179 a_18546_60188# a_29114_60146# 0.35fF
C12180 VDD a_5595_65301# 1.08fF
C12181 VDD a_18162_60186# 2.73fF
C12182 pmat.row_n[6] pmat.rowoff_n[5] 0.35fF
C12183 a_8583_29199# nmat.col_n[3] 0.30fF
C12184 pmat.sample_n vcm 1.15fF
C12185 m2_43032_7214# m3_43164_7346# 2.79fF
C12186 a_10223_26703# a_8013_25615# 0.86fF
C12187 VDD _1154_.X 33.49fF
C12188 nmat.col_n[29] m2_48052_24282# 0.43fF
C12189 m2_20944_54946# m3_21076_55078# 2.79fF
C12190 a_1957_43567# a_2411_43301# 0.31fF
C12191 a_31214_68178# a_31214_67174# 1.00fF
C12192 a_5651_66975# a_8841_60405# 0.73fF
C12193 a_36234_23548# vcm 0.65fF
C12194 a_27198_69182# ctopp 3.58fF
C12195 a_38242_9492# vcm 0.65fF
C12196 VDD a_36234_69182# 0.52fF
C12197 VDD a_3415_9839# 0.39fF
C12198 VDD a_11067_49871# 4.07fF
C12199 a_24591_28327# a_19405_28853# 2.84fF
C12200 VDD a_42024_46805# 0.98fF
C12201 a_36234_59142# ctopp 3.58fF
C12202 a_30210_11500# ctopn 3.58fF
C12203 a_19166_69182# a_19166_68178# 1.00fF
C12204 VDD a_45270_59142# 0.52fF
C12205 VDD a_28171_35561# 0.63fF
C12206 a_11435_58791# nmat.rowon_n[6] 0.41fF
C12207 a_29206_16520# a_30210_16520# 0.97fF
C12208 a_18546_16518# a_41162_16926# 0.35fF
C12209 a_37820_30485# a_43776_30287# 1.78fF
C12210 a_41731_49525# a_43533_30761# 0.38fF
C12211 pmat.row_n[7] a_3571_13627# 1.46fF
C12212 nmat.col[20] vcm 5.76fF
C12213 VDD a_22178_61150# 0.52fF
C12214 ANTENNA__1196__A2.DIODE a_83656_2767# 0.32fF
C12215 a_19233_38215# a_16981_37462# 0.31fF
C12216 a_34226_13508# vcm 0.65fF
C12217 VDD a_11041_40948# 2.15fF
C12218 ANTENNA__1187__B1.DIODE _1192_.B1 0.86fF
C12219 VDD vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top 109.34fF
C12220 m2_50060_7214# m2_51064_7214# 0.96fF
C12221 nmat.col_n[13] ANTENNA__1190__A2.DIODE 8.61fF
C12222 pmat.en_bit_n[2] ANTENNA__1395__A1.DIODE 0.41fF
C12223 a_12228_39605# cgen.dlycontrol2_in[0] 0.61fF
C12224 a_32218_18528# vcm 0.65fF
C12225 a_4128_64391# pmat.rowoff_n[4] 1.44fF
C12226 m2_51064_66994# vcm 0.51fF
C12227 VDD a_13459_4943# 0.42fF
C12228 nmat.col[15] nmat.col_n[30] 0.92fF
C12229 a_21174_20536# a_21174_19532# 1.00fF
C12230 a_3339_59879# a_6975_76823# 0.64fF
C12231 a_6283_31591# a_11784_47099# 0.60fF
C12232 a_13275_48783# a_40105_47375# 0.46fF
C12233 a_1781_9308# a_2411_16101# 0.61fF
C12234 VDD m3_51196_72146# 0.49fF
C12235 a_43262_15516# vcm 0.65fF
C12236 VDD a_28202_17524# 0.52fF
C12237 a_1586_33927# cgen.dlycontrol2_in[3] 1.56fF
C12238 a_11497_40719# a_11389_40443# 0.49fF
C12239 ANTENNA__1190__A1.DIODE ANTENNA__1197__B.DIODE 0.39fF
C12240 a_23395_53135# ANTENNA__1187__B1.DIODE 0.78fF
C12241 _1187_.A2 a_24867_53135# 0.49fF
C12242 ANTENNA__1190__B1.DIODE a_24591_28327# 0.49fF
C12243 VDD a_8749_47381# 0.61fF
C12244 a_1586_63927# a_2163_58941# 0.40fF
C12245 a_10515_13967# a_9963_13967# 4.17fF
C12246 m2_35000_72014# m3_35132_72146# 2.79fF
C12247 pmat.row_n[11] cgen.dlycontrol1_in[2] 0.44fF
C12248 a_38242_70186# a_38242_69182# 1.00fF
C12249 VDD a_29206_8488# 0.55fF
C12250 a_18546_21538# a_32126_21946# 0.35fF
C12251 a_27198_14512# a_27198_13508# 1.00fF
C12252 a_4351_55527# a_5651_66975# 0.88fF
C12253 VDD pmat.col[2] 5.06fF
C12254 a_38851_28327# nmat.col[29] 0.52fF
C12255 _1192_.B1 a_26479_32117# 0.31fF
C12256 a_39246_23548# ctopn 3.40fF
C12257 VDD a_45270_19532# 0.52fF
C12258 nmat.col[3] a_12463_22351# 0.49fF
C12259 a_41254_9492# ctopn 3.57fF
C12260 a_31214_57134# a_31214_56130# 1.00fF
C12261 a_35230_19532# a_36234_19532# 0.97fF
C12262 a_39246_60146# vcm 0.62fF
C12263 VDD a_44266_10496# 0.52fF
C12264 VDD a_18953_43493# 1.25fF
C12265 VDD a_7631_15253# 0.63fF
C12266 a_29937_31055# a_44763_34293# 0.36fF
C12267 a_13091_28327# a_13459_28111# 2.51fF
C12268 a_43776_30287# a_34204_27765# 0.31fF
C12269 a_18546_58180# a_51202_58138# 0.35fF
C12270 a_6975_76823# a_6292_69831# 0.40fF
C12271 VDD a_29493_31375# 0.30fF
C12272 a_14287_70543# pmat.row_n[3] 2.27fF
C12273 a_3866_57399# a_3770_57399# 0.59fF
C12274 a_18546_10494# a_51202_10902# 0.35fF
C12275 a_34226_10496# a_35230_10496# 0.97fF
C12276 VDD dummypin[6] 1.00fF
C12277 a_19166_16520# ctopn 3.43fF
C12278 VDD a_24186_12504# 0.52fF
C12279 VDD a_8491_47911# 10.75fF
C12280 a_45270_16520# vcm 0.65fF
C12281 m2_17932_21270# vcm 0.44fF
C12282 a_45270_56130# a_46274_56130# 0.97fF
C12283 VDD a_6835_51183# 1.05fF
C12284 a_37238_13508# ctopn 3.58fF
C12285 a_32218_57134# vcm 0.62fF
C12286 VDD a_10591_37737# 0.57fF
C12287 a_31214_71190# vcm 0.60fF
C12288 pmat.sample_n a_11067_49871# 0.78fF
C12289 a_35230_18528# ctopn 3.58fF
C12290 VDD a_12197_41570# 3.14fF
C12291 VDD a_14589_40726# 2.46fF
C12292 a_15667_27239# nmat.col_n[31] 0.31fF
C12293 a_50290_70186# ctopp 3.42fF
C12294 a_12069_38517# cgen.dlycontrol2_in[1] 1.40fF
C12295 a_2879_19093# a_3045_19093# 0.72fF
C12296 a_20170_9492# vcm 0.65fF
C12297 a_46274_15516# ctopn 3.58fF
C12298 VDD a_18546_69224# 32.63fF
C12299 VDD a_46274_11500# 0.52fF
C12300 _1179_.X ANTENNA__1190__B1.DIODE 0.74fF
C12301 a_27198_22544# a_28202_22544# 0.97fF
C12302 pmat.en_bit_n[2] ANTENNA__1395__A2.DIODE 2.65fF
C12303 VDD a_11823_46973# 0.45fF
C12304 a_48282_66170# a_49286_66170# 0.97fF
C12305 a_12345_39100# a_12543_39126# 0.30fF
C12306 pmat.row_n[11] a_2411_43301# 0.93fF
C12307 pmat.rowoff_n[6] ctopp 0.60fF
C12308 pmat.row_n[13] pmat.rowoff_n[13] 0.30fF
C12309 a_18546_69224# a_46182_69182# 0.35fF
C12310 VDD a_12107_62037# 0.67fF
C12311 a_20170_16520# a_21174_16520# 0.97fF
C12312 a_41254_63158# a_42258_63158# 0.97fF
C12313 m2_17932_22274# m3_18064_22406# 2.76fF
C12314 a_1957_43567# a_12907_54997# 0.70fF
C12315 a_18546_9490# a_19074_9898# 0.35fF
C12316 a_43262_22544# vcm 0.65fF
C12317 a_41254_68178# ctopp 3.58fF
C12318 nmat.col[28] comp_latch 0.65fF
C12319 a_10055_31591# a_13275_48783# 0.46fF
C12320 VDD a_50290_68178# 0.54fF
C12321 a_2659_35015# cgen.dlycontrol1_in[2] 0.44fF
C12322 nmat.rowon_n[12] nmat.col_n[12] 2.08fF
C12323 a_40250_62154# pmat.col[21] 0.31fF
C12324 a_24867_53135# pmat.col[1] 0.66fF
C12325 nmat.col[17] nmat.col_n[17] 0.65fF
C12326 VDD nmat.col_n[7] 8.04fF
C12327 ANTENNA__1190__B1.DIODE a_14917_23983# 0.89fF
C12328 a_13459_28111# a_17139_30503# 1.14fF
C12329 pmat.row_n[3] a_18162_11500# 25.57fF
C12330 VDD a_23182_56130# 0.55fF
C12331 VDD a_11391_69831# 0.38fF
C12332 a_48282_16520# ctopn 3.58fF
C12333 VDD a_2327_11477# 0.52fF
C12334 VDD m2_33996_7214# 0.93fF
C12335 a_6283_31591# a_2007_25597# 1.35fF
C12336 a_18546_62196# a_37146_62154# 0.35fF
C12337 a_4259_31375# a_8385_51727# 0.80fF
C12338 VDD a_22895_47893# 0.31fF
C12339 a_18546_66212# a_33130_66170# 0.35fF
C12340 a_18546_12502# ctopn 1.59fF
C12341 m2_51064_21270# m2_51064_20266# 0.99fF
C12342 a_49286_70186# a_50290_70186# 0.97fF
C12343 VDD a_44371_34319# 0.59fF
C12344 VDD a_26194_66170# 0.52fF
C12345 VDD a_9827_8181# 0.53fF
C12346 nmat.col[31] nmat.col[30] 0.63fF
C12347 a_36234_11500# a_37238_11500# 0.97fF
C12348 VDD a_13503_36893# 1.59fF
C12349 a_48282_56130# m2_48052_54946# 0.99fF
C12350 pmat.row_n[6] nmat.rowoff_n[8] 0.32fF
C12351 nmat.col_n[21] a_47011_31029# 0.48fF
C12352 a_10515_15055# a_10239_14183# 0.91fF
C12353 a_38242_64162# a_38242_63158# 1.00fF
C12354 a_11142_64783# a_11797_60431# 0.88fF
C12355 a_37820_30485# a_44774_40821# 0.70fF
C12356 a_41254_10496# a_41254_9492# 1.00fF
C12357 _1192_.A2 pmat.col[17] 0.41fF
C12358 ANTENNA__1395__B1.DIODE a_18547_51565# 0.74fF
C12359 a_33423_47695# a_7109_29423# 0.31fF
C12360 a_38391_47381# a_38557_47381# 0.42fF
C12361 pmat.en_bit_n[0] ANTENNA_fanout52_A.DIODE 2.72fF
C12362 a_38242_58138# a_38242_57134# 1.00fF
C12363 pmat.rowon_n[8] a_1586_33927# 0.32fF
C12364 VDD a_20848_39429# 1.24fF
C12365 a_10515_13967# a_18823_50247# 1.13fF
C12366 _1194_.B1 a_41321_30511# 0.36fF
C12367 pmat.col[20] ctopp 1.97fF
C12368 a_50290_64162# vcm 0.62fF
C12369 VDD m2_51064_23278# 1.05fF
C12370 VDD a_40837_46261# 10.39fF
C12371 a_45277_32687# a_47039_31599# 0.31fF
C12372 a_42258_60146# a_42258_59142# 1.00fF
C12373 a_30210_18528# a_30210_17524# 1.00fF
C12374 a_28915_50959# a_11948_49783# 0.44fF
C12375 VDD a_18235_34743# 0.63fF
C12376 a_13275_48783# a_13688_47893# 0.36fF
C12377 VDD a_8378_12691# 0.30fF
C12378 a_5173_9839# a_6763_13103# 0.33fF
C12379 a_2407_49289# a_4081_61127# 0.69fF
C12380 a_2411_16101# a_2603_22357# 0.34fF
C12381 a_46274_22544# ctopn 3.57fF
C12382 a_30210_63158# a_30210_62154# 1.00fF
C12383 m2_18936_23278# vcm 0.44fF
C12384 m2_17932_19262# m3_18064_19394# 2.76fF
C12385 VDD a_6895_48981# 0.38fF
C12386 a_46274_67174# a_47278_67174# 0.97fF
C12387 a_9581_56079# a_1586_50247# 0.89fF
C12388 VDD a_11041_38772# 1.60fF
C12389 a_18546_70228# a_35138_70186# 0.35fF
C12390 VDD a_24186_67174# 0.52fF
C12391 VDD a_15107_40183# 0.61fF
C12392 a_37827_30793# nmat.col[29] 0.34fF
C12393 a_2411_43301# a_2659_35015# 0.51fF
C12394 a_36234_22544# a_36234_21540# 1.00fF
C12395 a_43262_66170# a_43262_65166# 1.00fF
C12396 VDD a_4241_13653# 0.30fF
C12397 a_13145_26935# a_8013_25615# 0.47fF
C12398 a_35230_14512# a_36234_14512# 0.97fF
C12399 a_34226_62154# vcm 0.62fF
C12400 VDD a_8378_63827# 0.31fF
C12401 a_18546_55168# a_34134_55126# 0.39fF
C12402 a_30527_31573# a_9785_28879# 0.43fF
C12403 a_7047_31226# a_6909_31061# 0.46fF
C12404 a_18546_17522# a_30118_17930# 0.35fF
C12405 a_34226_64162# a_35230_64162# 0.97fF
C12406 a_18546_64204# a_51202_64162# 0.35fF
C12407 _1224_.X ANTENNA__1183__B1.DIODE 1.50fF
C12408 a_40250_68178# a_41254_68178# 0.97fF
C12409 a_18546_57176# a_26102_57134# 0.35fF
C12410 VDD nmat.col_n[0] 5.46fF
C12411 VDD a_3496_51701# 0.69fF
C12412 a_37238_8488# m2_37008_7214# 1.00fF
C12413 a_29206_13508# a_29206_12504# 1.00fF
C12414 pmat.rowon_n[3] a_2983_48071# 0.58fF
C12415 a_18546_22542# a_18162_22544# 2.61fF
C12416 a_18546_15514# a_30118_15922# 0.35fF
C12417 a_4383_7093# a_10995_17782# 0.30fF
C12418 a_49286_60146# ctopp 3.57fF
C12419 pmat.rowoff_n[7] nmat.rowon_n[14] 2.36fF
C12420 VDD pmat.rowoff_n[5] 2.18fF
C12421 VDD a_33309_36039# 1.26fF
C12422 a_33222_70186# vcm 0.62fF
C12423 pmat.en_bit_n[0] a_25681_28879# 0.83fF
C12424 pmat.row_n[9] nmat.rowon_n[6] 20.96fF
C12425 ANTENNA__1187__B1.DIODE a_30663_50087# 0.57fF
C12426 nmat.en_bit_n[1] a_22199_30287# 1.07fF
C12427 pmat.rowon_n[7] a_13643_29415# 0.65fF
C12428 a_40105_47375# a_1781_9308# 0.77fF
C12429 pmat.col_n[3] vcm 2.80fF
C12430 a_22178_19532# ctopn 3.58fF
C12431 VDD a_44739_43567# 0.37fF
C12432 a_11041_40948# a_11113_40835# 0.32fF
C12433 ANTENNA__1395__B1.DIODE ANTENNA__1190__A2.DIODE 2.13fF
C12434 VDD a_21365_27247# 1.60fF
C12435 VDD a_22178_21540# 0.52fF
C12436 a_18546_59184# a_46182_59142# 0.35fF
C12437 a_36234_65166# a_36234_64162# 1.00fF
C12438 ANTENNA__1195__A1.DIODE a_16311_28327# 1.36fF
C12439 m2_17932_70006# vcm 0.44fF
C12440 a_21174_10496# ctopn 3.58fF
C12441 a_42258_57134# ctopp 3.57fF
C12442 VDD a_9595_30511# 0.40fF
C12443 a_41254_71190# ctopp 3.40fF
C12444 cgen.dlycontrol4_in[1] a_3325_23439# 0.42fF
C12445 a_28202_58138# ctopp 3.58fF
C12446 a_24186_68178# vcm 0.62fF
C12447 VDD a_50290_71190# 0.58fF
C12448 a_11067_16359# cgen.dlycontrol4_in[4] 0.37fF
C12449 VDD a_37238_58138# 0.52fF
C12450 a_45270_23548# a_46274_23548# 0.97fF
C12451 a_13503_43421# a_12237_38772# 0.71fF
C12452 cgen.dlycontrol4_in[1] a_11497_40719# 3.67fF
C12453 VDD a_5047_76983# 0.85fF
C12454 a_25190_16520# a_25190_15516# 1.00fF
C12455 a_18546_62196# a_18162_62194# 2.62fF
C12456 VDD a_33685_48437# 0.61fF
C12457 a_47278_9492# a_48282_9492# 0.97fF
C12458 a_18546_60188# a_22086_60146# 0.35fF
C12459 VDD a_5682_56311# 3.23fF
C12460 a_2315_44124# a_4313_44111# 0.37fF
C12461 _1194_.A2 nmat.col_n[13] 0.94fF
C12462 m2_17932_9222# vcm 0.44fF
C12463 pmat.en_bit_n[0] a_13641_23439# 1.40fF
C12464 VDD a_53622_39932# 0.37fF
C12465 a_1899_35051# a_4257_34319# 0.54fF
C12466 a_1923_53055# a_2163_53057# 0.32fF
C12467 a_29206_23548# vcm 0.65fF
C12468 nmat.col[19] nmat.col_n[24] 0.61fF
C12469 a_20170_69182# ctopp 3.57fF
C12470 a_31214_9492# vcm 0.65fF
C12471 VDD a_29206_69182# 0.52fF
C12472 a_6283_31591# a_7109_29423# 1.75fF
C12473 VDD a_12539_10389# 0.52fF
C12474 a_47278_23548# m2_47048_24282# 0.99fF
C12475 a_19166_12504# a_20170_12504# 0.97fF
C12476 a_18546_22542# a_48190_22950# 0.35fF
C12477 pmat.row_n[15] cgen.dlycontrol4_in[5] 0.83fF
C12478 VDD a_25209_44581# 1.14fF
C12479 a_5403_67655# a_6451_67655# 0.33fF
C12480 VDD m2_31988_24282# 0.62fF
C12481 a_22199_32149# a_2007_25597# 0.35fF
C12482 ANTENNA__1190__B1.DIODE nmat.sample_n 2.45fF
C12483 a_47278_20536# vcm 0.65fF
C12484 a_37238_65166# a_38242_65166# 0.97fF
C12485 a_29206_59142# ctopp 3.58fF
C12486 pmat.rowon_n[0] a_5558_9527# 0.58fF
C12487 a_23182_11500# ctopn 3.58fF
C12488 VDD a_33331_31599# 0.40fF
C12489 VDD ANTENNA__1190__A1.DIODE 21.57fF
C12490 VDD a_38242_59142# 0.52fF
C12491 a_44266_21540# a_45270_21540# 0.97fF
C12492 VDD a_13259_35561# 0.60fF
C12493 a_25879_31591# clk_ena 0.95fF
C12494 a_18546_16518# a_34134_16926# 0.35fF
C12495 a_2952_25045# a_5991_23983# 0.35fF
C12496 a_11067_64015# a_11067_30287# 0.97fF
C12497 a_45270_71190# a_45270_70186# 1.00fF
C12498 pmat.row_n[1] a_14195_7351# 0.42fF
C12499 a_20438_35431# a_11297_36091# 0.65fF
C12500 a_27198_13508# vcm 0.65fF
C12501 a_1591_40853# a_1895_41018# 0.61fF
C12502 m2_43032_7214# m2_44036_7214# 0.96fF
C12503 a_2007_25597# a_2648_29397# 1.12fF
C12504 a_25190_18528# vcm 0.65fF
C12505 VDD a_6448_5755# 0.40fF
C12506 VDD a_14465_29575# 0.54fF
C12507 a_6283_31591# cgen.dlycontrol4_in[5] 0.46fF
C12508 nmat.col_n[2] vcm 2.80fF
C12509 a_43262_13508# a_44266_13508# 0.97fF
C12510 VDD m3_23084_72146# 0.39fF
C12511 a_36234_15516# vcm 0.65fF
C12512 _1224_.X pmat.col[30] 0.57fF
C12513 VDD a_21174_17524# 0.52fF
C12514 a_2263_43719# a_1823_58237# 0.79fF
C12515 VDD a_8507_20175# 0.52fF
C12516 a_30571_50959# a_30111_47911# 0.32fF
C12517 a_41254_18528# a_42258_18528# 0.97fF
C12518 VDD a_22178_8488# 0.55fF
C12519 a_18546_21538# a_25098_21946# 0.35fF
C12520 VDD a_29183_36919# 0.61fF
C12521 a_28202_62154# a_28202_61150# 1.00fF
C12522 VDD a_3707_53903# 0.47fF
C12523 a_32218_23548# ctopn 3.40fF
C12524 VDD a_38242_19532# 0.52fF
C12525 a_10515_61839# a_10239_14183# 1.72fF
C12526 pmat.row_n[6] pmat.row_n[5] 0.70fF
C12527 a_34226_9492# ctopn 3.57fF
C12528 VDD m2_51064_72014# 1.84fF
C12529 a_10471_12791# comp_latch 0.41fF
C12530 VDD a_3923_68021# 3.68fF
C12531 a_32218_60146# vcm 0.62fF
C12532 VDD a_37238_10496# 0.52fF
C12533 a_12513_39100# cgen.dlycontrol1_in[4] 0.77fF
C12534 a_33423_47695# nmat.col_n[21] 0.53fF
C12535 a_50290_20536# ctopn 3.43fF
C12536 VDD a_2021_26677# 2.09fF
C12537 a_28202_15516# a_28202_14512# 1.00fF
C12538 a_7939_7125# a_8105_7125# 0.75fF
C12539 a_18546_58180# a_44174_58138# 0.35fF
C12540 a_30210_69182# a_30210_68178# 1.00fF
C12541 a_1717_13647# comp_latch 0.39fF
C12542 a_18546_10494# a_44174_10902# 0.35fF
C12543 a_38242_21540# a_38242_20536# 1.00fF
C12544 VDD a_14923_34473# 0.64fF
C12545 a_44266_62154# ctopp 3.58fF
C12546 VDD m2_51064_11230# 1.17fF
C12547 a_38242_16520# vcm 0.65fF
C12548 a_10781_42869# cgen.start_conv_in 2.90fF
C12549 nmat.col[19] ctopn 2.00fF
C12550 a_12693_38543# a_16890_36911# 0.39fF
C12551 pmat.row_n[12] pmat.row_n[0] 7.95fF
C12552 a_30210_13508# ctopn 3.58fF
C12553 _1192_.B1 a_18243_28327# 0.69fF
C12554 a_1781_9308# a_3183_19258# 0.63fF
C12555 a_25190_57134# vcm 0.62fF
C12556 VDD a_29220_37253# 1.40fF
C12557 a_24186_71190# vcm 0.60fF
C12558 a_28202_18528# ctopn 3.58fF
C12559 VDD a_40352_41831# 1.65fF
C12560 a_9411_2215# a_9528_20407# 0.35fF
C12561 a_11435_58791# nmat.rowon_n[13] 0.32fF
C12562 VDD a_2839_38101# 1.30fF
C12563 a_43262_70186# ctopp 3.57fF
C12564 a_39246_15516# ctopn 3.58fF
C12565 a_46523_39733# a_45019_38645# 0.47fF
C12566 VDD a_39246_11500# 0.52fF
C12567 m3_34128_55078# ctopp 0.39fF
C12568 a_23395_53135# a_18243_28327# 3.18fF
C12569 a_49286_23548# a_49286_22544# 1.00fF
C12570 VDD m2_27972_54946# 0.62fF
C12571 a_3615_71631# a_12604_47080# 0.40fF
C12572 VDD a_34768_47375# 0.44fF
C12573 a_48282_60146# a_49286_60146# 0.97fF
C12574 m2_51064_71010# m3_51196_71142# 2.76fF
C12575 a_18546_69224# a_39154_69182# 0.35fF
C12576 pmat.col_n[11] ctopp 2.02fF
C12577 VDD pmat.col[6] 4.63fF
C12578 a_32218_11500# a_32218_10496# 1.00fF
C12579 VDD a_37146_72194# 0.32fF
C12580 _1154_.A a_41731_49525# 0.93fF
C12581 VDD nmat.rowoff_n[8] 2.39fF
C12582 cgen.dlycontrol4_in[5] a_11041_39860# 1.24fF
C12583 a_9405_66627# a_1586_63927# 0.41fF
C12584 a_11497_38543# a_14773_38306# 0.48fF
C12585 pmat.row_n[1] a_13091_52047# 0.78fF
C12586 pmat.rowoff_n[12] a_9963_13967# 0.52fF
C12587 a_36234_22544# vcm 0.65fF
C12588 a_37238_61150# a_38242_61150# 0.97fF
C12589 a_34226_68178# ctopp 3.58fF
C12590 VDD a_43262_68178# 0.52fF
C12591 a_13503_37981# a_14773_38306# 0.60fF
C12592 a_22178_12504# a_22178_11500# 1.00fF
C12593 a_50290_63158# vcm 0.62fF
C12594 a_11115_71285# a_11203_62037# 1.09fF
C12595 pmat.en_bit_n[2] a_2007_25597# 0.68fF
C12596 a_14287_69455# pmat.rowoff_n[8] 0.46fF
C12597 a_1823_76181# a_1823_74557# 1.56fF
C12598 a_10239_14183# a_6634_26133# 0.31fF
C12599 a_18546_20534# a_45178_20942# 0.35fF
C12600 a_31214_20536# a_32218_20536# 0.97fF
C12601 VDD a_2163_69821# 0.48fF
C12602 a_41254_16520# ctopn 3.58fF
C12603 a_12447_16143# a_4075_31591# 0.66fF
C12604 a_34226_24552# m2_32992_24282# 0.96fF
C12605 VDD a_2847_28095# 0.62fF
C12606 VDD m2_19940_7214# 1.09fF
C12607 a_18546_62196# a_30118_62154# 0.35fF
C12608 _1224_.X a_21215_48071# 0.34fF
C12609 _1183_.A2 a_29937_31055# 1.17fF
C12610 a_44266_67174# a_44266_66170# 1.00fF
C12611 a_18546_66212# a_26102_66170# 0.35fF
C12612 a_30210_9492# a_30210_8488# 1.00fF
C12613 VDD a_48282_23548# 0.55fF
C12614 VDD a_50290_9492# 0.54fF
C12615 a_1895_36666# a_1757_36501# 0.55fF
C12616 a_18546_11498# a_48190_11906# 0.35fF
C12617 VDD a_11317_36924# 7.46fF
C12618 VDD a_82787_14709# 0.31fF
C12619 pmat.rowoff_n[7] cgen.dlycontrol1_in[1] 0.59fF
C12620 m2_48052_7214# m3_48184_7346# 2.79fF
C12621 VDD a_20170_19532# 0.52fF
C12622 a_43262_17524# a_44266_17524# 0.97fF
C12623 a_3576_17143# a_4865_12533# 0.61fF
C12624 m2_25964_54946# m3_26096_55078# 2.79fF
C12625 a_41254_57134# a_42258_57134# 0.97fF
C12626 a_14641_57711# pmat.rowoff_n[9] 0.71fF
C12627 a_46274_20536# a_46274_19532# 1.00fF
C12628 a_40250_71190# a_41254_71190# 0.97fF
C12629 ANTENNA__1197__B.DIODE nmat.col[12] 1.24fF
C12630 a_27198_58138# a_28202_58138# 0.97fF
C12631 a_44266_14512# vcm 0.65fF
C12632 a_43262_64162# vcm 0.62fF
C12633 a_40837_46261# a_43533_30761# 0.33fF
C12634 _1196_.B1 nmat.col_n[31] 0.52fF
C12635 a_44266_8488# a_45270_8488# 0.97fF
C12636 m2_51064_67998# m3_51196_68130# 2.76fF
C12637 VDD a_36919_31849# 0.41fF
C12638 a_10873_36341# a_11921_35286# 0.33fF
C12639 VDD a_4227_34293# 0.42fF
C12640 VDD a_46274_13508# 0.52fF
C12641 pmat.rowon_n[8] a_6467_29415# 1.00fF
C12642 a_39246_22544# ctopn 3.57fF
C12643 a_20170_16520# vcm 0.65fF
C12644 VDD a_44266_18528# 0.52fF
C12645 a_15667_27239# _1183_.A2 1.61fF
C12646 VDD a_33281_49551# 0.63fF
C12647 a_9675_10396# comp_latch 0.39fF
C12648 a_27198_61150# a_27198_60146# 1.00fF
C12649 pmat.row_n[12] nmat.sample 0.35fF
C12650 a_35230_19532# a_35230_18528# 1.00fF
C12651 m2_17932_23278# m2_17932_22274# 0.99fF
C12652 a_18546_70228# a_28110_70186# 0.35fF
C12653 ANTENNA__1190__A2.DIODE nmat.col[18] 6.60fF
C12654 VDD a_12585_40443# 1.56fF
C12655 m2_51064_70006# m2_51064_69002# 0.99fF
C12656 a_2007_25597# a_4068_25615# 0.54fF
C12657 _1194_.A2 ANTENNA__1395__B1.DIODE 1.27fF
C12658 VDD a_12047_14165# 0.56fF
C12659 a_18546_14510# a_46182_14918# 0.35fF
C12660 a_27198_62154# vcm 0.62fF
C12661 a_18546_17522# a_23090_17930# 0.35fF
C12662 a_18546_64204# a_44174_64162# 0.35fF
C12663 ANTENNA__1187__B1.DIODE a_10883_3303# 0.74fF
C12664 a_6927_30503# a_2411_43301# 0.94fF
C12665 VDD a_14471_3561# 0.39fF
C12666 a_28202_59142# a_28202_58138# 1.00fF
C12667 a_3615_71631# a_12719_69367# 0.56fF
C12668 a_1739_47893# cgen.dlycontrol3_in[1] 1.04fF
C12669 nmat.col[7] a_7026_24527# 1.26fF
C12670 VDD a_6323_26409# 0.60fF
C12671 VDD m3_18064_64114# 0.33fF
C12672 VDD dummypin[1] 1.15fF
C12673 a_18546_15514# a_23090_15922# 0.35fF
C12674 a_46274_65166# vcm 0.62fF
C12675 a_26194_63158# pmat.col[7] 0.31fF
C12676 a_42258_60146# ctopp 3.58fF
C12677 m2_40020_72014# m3_40152_72146# 2.79fF
C12678 VDD a_17959_36649# 0.60fF
C12679 VDD _0467_ 0.96fF
C12680 a_3866_57399# a_5779_71285# 0.44fF
C12681 a_26194_70186# vcm 0.62fF
C12682 VDD pmat.col_n[4] 5.21fF
C12683 a_1899_35051# a_4985_51433# 0.30fF
C12684 pmat.col[7] vcm 5.88fF
C12685 a_34226_56130# a_34226_55126# 1.00fF
C12686 a_33222_17524# a_33222_16520# 1.00fF
C12687 VDD a_6564_24527# 0.40fF
C12688 a_47278_14512# ctopn 3.58fF
C12689 pmat.en_bit_n[0] a_17139_30503# 0.36fF
C12690 a_39246_12504# a_40250_12504# 0.97fF
C12691 a_10873_38517# a_10873_36341# 0.73fF
C12692 a_15667_27239# a_34204_27765# 0.78fF
C12693 a_11711_50959# a_11455_50237# 0.50fF
C12694 _1179_.X clk_ena 4.05fF
C12695 m2_51064_9222# m2_51064_8218# 0.99fF
C12696 a_13091_52047# a_25839_49783# 0.69fF
C12697 pmat.col_n[0] pmat.col[0] 0.73fF
C12698 VDD a_41443_28879# 0.34fF
C12699 VDD a_8305_20871# 6.22fF
C12700 a_18546_59184# a_39154_59142# 0.35fF
C12701 a_28202_59142# a_29206_59142# 0.97fF
C12702 m2_51064_64986# m3_51196_65118# 2.76fF
C12703 a_35230_57134# ctopp 3.58fF
C12704 VDD a_38851_30761# 0.44fF
C12705 a_8031_76757# a_8197_76757# 0.42fF
C12706 a_6975_76823# a_2149_45717# 0.41fF
C12707 a_34226_71190# ctopp 3.40fF
C12708 VDD a_44266_57134# 0.52fF
C12709 a_21174_58138# ctopp 3.58fF
C12710 VDD a_43262_71190# 0.55fF
C12711 a_30111_47911# a_35786_47893# 0.75fF
C12712 VDD a_30210_58138# 0.52fF
C12713 a_38851_28327# nmat.col[30] 0.55fF
C12714 VDD a_9871_48463# 0.48fF
C12715 m2_51064_19262# vcm 0.51fF
C12716 VDD a_5053_59575# 1.17fF
C12717 cgen.dlycontrol2_in[0] a_12934_35823# 0.52fF
C12718 VDD a_7355_37013# 0.38fF
C12719 a_11067_16359# a_11711_50959# 0.99fF
C12720 a_19166_12504# vcm 0.65fF
C12721 a_1899_35051# a_1586_50247# 0.62fF
C12722 a_31214_56130# m2_30984_54946# 0.99fF
C12723 a_12447_16143# a_7644_16341# 0.59fF
C12724 a_18546_24550# a_44174_24958# 0.35fF
C12725 a_2007_25597# a_35559_30209# 0.33fF
C12726 a_17139_30503# a_44573_45173# 0.95fF
C12727 nmat.col[15] vcm 5.76fF
C12728 a_24186_68178# a_24186_67174# 1.00fF
C12729 _1154_.A vcm 0.76fF
C12730 a_22178_23548# vcm 0.65fF
C12731 a_24186_9492# vcm 0.65fF
C12732 VDD a_22178_69182# 0.52fF
C12733 a_46274_61150# vcm 0.62fF
C12734 a_12263_50959# a_6283_31591# 0.39fF
C12735 ANTENNA__1395__A1.DIODE a_15667_27239# 0.37fF
C12736 VDD m3_18064_11362# 0.32fF
C12737 a_18546_22542# a_41162_22950# 0.35fF
C12738 a_40250_20536# vcm 0.65fF
C12739 a_22178_59142# ctopp 3.58fF
C12740 ANTENNA__1190__A1.DIODE a_43533_30761# 0.36fF
C12741 VDD a_2422_29575# 0.58fF
C12742 a_2419_53351# a_3746_58487# 1.21fF
C12743 VDD a_31214_59142# 0.52fF
C12744 a_20170_21540# a_20170_20536# 1.00fF
C12745 pmat.row_n[7] a_13091_52047# 0.73fF
C12746 VDD pmat.row_n[5] 19.70fF
C12747 VDD m2_17932_14242# 1.00fF
C12748 a_18546_23546# a_18162_23548# 2.61fF
C12749 nmat.rowoff_n[6] a_11897_21263# 0.60fF
C12750 a_22178_16520# a_23182_16520# 0.97fF
C12751 a_18546_16518# a_27106_16926# 0.35fF
C12752 m2_32992_54946# vcm 0.42fF
C12753 a_2935_38279# a_6369_39465# 0.47fF
C12754 pmat.rowon_n[8] a_9135_60967# 0.66fF
C12755 pmat.row_n[4] a_18546_60188# 0.35fF
C12756 a_1781_9308# a_32827_46805# 0.54fF
C12757 a_3305_27791# a_4712_27023# 0.42fF
C12758 nmat.rowon_n[14] cgen.dlycontrol1_in[1] 1.88fF
C12759 m2_36004_7214# m2_37008_7214# 0.96fF
C12760 a_24374_29941# a_22628_30485# 0.42fF
C12761 m2_51064_61974# m3_51196_62106# 2.76fF
C12762 a_30111_47911# a_46968_45743# 0.32fF
C12763 a_29206_15516# vcm 0.65fF
C12764 VDD a_9319_50639# 0.52fF
C12765 a_3063_14741# a_3229_14741# 0.61fF
C12766 VDD a_46487_47919# 0.53fF
C12767 a_31214_70186# a_31214_69182# 1.00fF
C12768 VDD a_4043_33535# 0.53fF
C12769 _1194_.B1 a_11711_50959# 0.70fF
C12770 pmat.rowoff_n[4] nmat.en_bit_n[1] 0.38fF
C12771 a_18546_56172# vcm 0.40fF
C12772 VDD a_16890_36911# 0.90fF
C12773 a_48282_12504# vcm 0.65fF
C12774 a_22459_28879# nmat.col[12] 0.33fF
C12775 a_13641_23439# a_10147_29415# 0.43fF
C12776 a_25190_23548# ctopn 3.40fF
C12777 VDD a_31214_19532# 0.52fF
C12778 a_24407_31375# nmat.col[21] 0.52fF
C12779 a_27198_9492# ctopn 3.57fF
C12780 VDD m2_37008_72014# 0.98fF
C12781 a_24186_57134# a_24186_56130# 1.00fF
C12782 ANTENNA__1195__A1.DIODE a_24407_31375# 1.17fF
C12783 a_28202_19532# a_29206_19532# 0.97fF
C12784 a_25190_60146# vcm 0.62fF
C12785 VDD a_30210_10496# 0.52fF
C12786 a_43262_20536# ctopn 3.58fF
C12787 VDD a_33489_44219# 1.24fF
C12788 a_32957_30287# a_33684_32143# 0.35fF
C12789 a_6283_31591# clk_ena 1.72fF
C12790 VDD a_13739_51701# 0.53fF
C12791 a_19166_59142# a_20170_59142# 0.97fF
C12792 a_30543_40721# a_20221_40835# 1.74fF
C12793 a_2215_47375# a_4979_38127# 0.61fF
C12794 a_18546_58180# a_37146_58138# 0.35fF
C12795 VDD a_1957_43567# 8.18fF
C12796 a_12934_35823# cgen.dlycontrol1_in[2] 0.44fF
C12797 a_27198_10496# a_28202_10496# 0.97fF
C12798 a_18546_10494# a_37146_10902# 0.35fF
C12799 ANTENNA__1395__A2.DIODE a_15667_27239# 0.39fF
C12800 a_37238_62154# ctopp 3.58fF
C12801 VDD a_46274_62154# 0.52fF
C12802 a_31214_16520# vcm 0.65fF
C12803 VDD a_23815_48981# 0.30fF
C12804 a_38242_56130# a_39246_56130# 0.97fF
C12805 a_10878_58487# a_11007_58229# 0.45fF
C12806 a_18162_67214# ctopp 1.49fF
C12807 a_23182_13508# ctopn 3.58fF
C12808 VDD a_11731_8751# 0.38fF
C12809 VDD a_29772_40517# 1.28fF
C12810 a_2935_38279# cgen.dlycontrol2_in[2] 0.75fF
C12811 _1154_.A _1154_.X 3.05fF
C12812 VDD a_10867_38007# 0.59fF
C12813 pmat.sw _1179_.X 0.39fF
C12814 nmat.sw a_4516_21531# 1.64fF
C12815 a_21174_18528# ctopn 3.58fF
C12816 pmat.sw a_33423_47695# 1.04fF
C12817 a_24374_29941# a_23021_29199# 0.48fF
C12818 m2_51064_58962# m3_51196_59094# 2.76fF
C12819 a_4128_46983# cgen.dlycontrol4_in[5] 0.93fF
C12820 a_2419_69455# a_3746_58487# 0.72fF
C12821 ANTENNA__1196__A2.DIODE a_29937_31055# 1.07fF
C12822 a_36234_70186# ctopp 3.57fF
C12823 VDD a_45270_70186# 0.52fF
C12824 a_32218_15516# ctopn 3.58fF
C12825 VDD a_32218_11500# 0.52fF
C12826 a_30210_23548# m2_29980_24282# 0.99fF
C12827 a_6467_29415# a_9307_31068# 0.95fF
C12828 cgen.enable_dlycontrol_in a_25755_34343# 0.86fF
C12829 pmat.col_n[21] _1179_.X 0.40fF
C12830 VDD a_44628_45717# 0.45fF
C12831 pmat.rowoff_n[12] a_18162_20536# 1.33fF
C12832 a_43262_62154# a_44266_62154# 0.97fF
C12833 a_50290_16520# a_50290_15516# 1.00fF
C12834 a_41254_66170# a_42258_66170# 0.97fF
C12835 VDD a_6803_77269# 0.35fF
C12836 a_18546_69224# a_32126_69182# 0.35fF
C12837 nmat.col_n[29] ctopn 2.05fF
C12838 a_47278_56130# vcm 0.62fF
C12839 VDD a_47035_36495# 0.38fF
C12840 pmat.col[31] vcm 6.48fF
C12841 cgen.dlycontrol1_in[2] config_2_in[3] 0.31fF
C12842 a_2263_43719# cgen.dlycontrol3_in[2] 1.87fF
C12843 a_34226_63158# a_35230_63158# 0.97fF
C12844 a_18546_63200# a_51202_63158# 0.35fF
C12845 a_9411_2215# a_32405_32463# 0.44fF
C12846 a_29206_22544# vcm 0.65fF
C12847 a_27198_68178# ctopp 3.58fF
C12848 VDD config_2_in[7] 1.05fF
C12849 a_50290_66170# vcm 0.62fF
C12850 VDD a_36234_68178# 0.52fF
C12851 a_23821_35279# clk_dig 0.54fF
C12852 a_37820_30485# a_35312_31599# 1.29fF
C12853 a_10767_39087# a_11773_39087# 0.94fF
C12854 pmat.col_n[6] vcm 2.80fF
C12855 VDD a_19166_15516# 0.56fF
C12856 a_43262_63158# vcm 0.62fF
C12857 VDD a_18162_65206# 2.73fF
C12858 VDD nmat.col[12] 7.61fF
C12859 pmat.col[31] _1194_.B1 0.50fF
C12860 ANTENNA__1196__A2.DIODE a_15667_27239# 1.67fF
C12861 VDD a_10287_29941# 0.44fF
C12862 nmat.sample_n clk_ena 0.38fF
C12863 pmat.col_n[26] ANTENNA__1190__B1.DIODE 0.48fF
C12864 ANTENNA__1187__B1.DIODE clk_vcm 0.39fF
C12865 a_18546_20534# a_38150_20942# 0.35fF
C12866 a_13275_48783# a_13643_29415# 1.33fF
C12867 a_34226_16520# ctopn 3.58fF
C12868 VDD pmat.row_n[13] 21.01fF
C12869 a_5687_71829# a_3615_71631# 0.36fF
C12870 VDD cgen.enable_dlycontrol_in 10.99fF
C12871 a_18546_62196# a_23090_62154# 0.35fF
C12872 VDD a_30409_48463# 0.40fF
C12873 VDD a_41254_23548# 0.55fF
C12874 a_42258_70186# a_43262_70186# 0.97fF
C12875 VDD a_3410_66003# 0.32fF
C12876 VDD a_43262_9492# 0.52fF
C12877 a_29206_11500# a_30210_11500# 0.97fF
C12878 a_18546_11498# a_41162_11906# 0.35fF
C12879 a_4075_50087# a_4985_51433# 0.51fF
C12880 pmat.col_n[16] pmat.col[16] 0.64fF
C12881 nmat.col[31] a_31263_28309# 0.77fF
C12882 ANTENNA__1197__A.DIODE nmat.col[29] 0.57fF
C12883 a_30571_50959# a_30663_50087# 3.07fF
C12884 a_22628_30485# a_22459_28879# 0.31fF
C12885 VDD a_4135_19391# 0.39fF
C12886 a_31214_64162# a_31214_63158# 1.00fF
C12887 a_34226_10496# a_34226_9492# 1.00fF
C12888 nmat.col_n[22] nmat.col[22] 0.70fF
C12889 a_48282_67174# vcm 0.62fF
C12890 a_31214_58138# a_31214_57134# 1.00fF
C12891 a_16083_50069# a_13275_48783# 0.51fF
C12892 ANTENNA__1195__A1.DIODE a_17842_27497# 0.38fF
C12893 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[29] 2.48fF
C12894 a_37238_14512# vcm 0.65fF
C12895 a_7840_27247# _0467_ 0.38fF
C12896 a_5687_71829# a_3339_70759# 0.60fF
C12897 inp_analog ANTENNA__1197__B.DIODE 0.65fF
C12898 a_36234_64162# vcm 0.62fF
C12899 VDD m2_41024_24282# 0.62fF
C12900 a_35230_60146# a_35230_59142# 1.00fF
C12901 a_23182_18528# a_23182_17524# 1.00fF
C12902 a_14287_69455# pmat.rowon_n[12] 0.33fF
C12903 pmat.row_n[12] a_18162_68218# 25.57fF
C12904 a_11041_36596# cgen.dlycontrol1_in[1] 1.22fF
C12905 VDD a_5211_57172# 1.27fF
C12906 VDD a_4991_69831# 7.98fF
C12907 VDD a_39246_13508# 0.52fF
C12908 a_19166_62154# ctopp 3.43fF
C12909 a_35312_31599# a_34204_27765# 0.99fF
C12910 a_32218_22544# ctopn 3.57fF
C12911 a_13459_28111# a_25879_31591# 0.98fF
C12912 VDD a_37238_18528# 0.52fF
C12913 a_23182_63158# a_23182_62154# 1.00fF
C12914 m2_22952_24282# vcm 0.42fF
C12915 VDD a_15839_49525# 0.43fF
C12916 a_39246_67174# a_40250_67174# 0.97fF
C12917 a_2149_45717# pmat.rowoff_n[7] 0.55fF
C12918 a_18546_70228# a_21082_70186# 0.35fF
C12919 VDD pmat.row_n[11] 13.48fF
C12920 m2_51064_19262# m3_51196_19394# 2.76fF
C12921 a_3339_59879# a_10049_60663# 0.37fF
C12922 VDD a_18162_61190# 2.73fF
C12923 a_14773_38306# a_14712_37429# 0.73fF
C12924 a_3339_70759# a_4583_68021# 1.63fF
C12925 pmat.rowon_n[8] nmat.rowon_n[7] 20.80fF
C12926 pmat.row_n[10] pmat.rowoff_n[10] 0.42fF
C12927 a_36234_66170# a_36234_65166# 1.00fF
C12928 a_29206_22544# a_29206_21540# 1.00fF
C12929 VDD a_48282_15516# 0.52fF
C12930 a_28202_14512# a_29206_14512# 0.97fF
C12931 a_18546_14510# a_39154_14918# 0.35fF
C12932 a_20170_62154# vcm 0.62fF
C12933 a_18546_55168# a_20078_55126# 0.39fF
C12934 a_18546_64204# a_37146_64162# 0.35fF
C12935 a_27198_64162# a_28202_64162# 0.97fF
C12936 VDD a_1761_2767# 1.04fF
C12937 a_33222_68178# a_34226_68178# 0.97fF
C12938 a_3663_9269# a_4865_8181# 0.33fF
C12939 a_18546_70228# ctopp 1.57fF
C12940 a_19166_20536# a_19166_19532# 1.00fF
C12941 VDD a_5445_11177# 0.42fF
C12942 a_22178_13508# a_22178_12504# 1.00fF
C12943 _1154_.X pmat.col[31] 0.47fF
C12944 VDD a_5931_74183# 0.50fF
C12945 a_39246_65166# vcm 0.62fF
C12946 ANTENNA__1395__A1.DIODE a_11067_27239# 0.43fF
C12947 a_46274_21540# vcm 0.65fF
C12948 a_1781_9308# a_2199_13887# 1.08fF
C12949 VDD nmat.rowon_n[1] 4.20fF
C12950 a_35230_60146# ctopp 3.58fF
C12951 VDD a_44266_60146# 0.52fF
C12952 VDD a_14833_72049# 0.38fF
C12953 a_7415_29397# a_10814_29111# 0.51fF
C12954 a_21739_29415# ANTENNA__1183__B1.DIODE 3.58fF
C12955 cgen.dlycontrol3_in[4] cgen.dlycontrol2_in[0] 0.68fF
C12956 m2_21948_24282# m3_22080_24414# 2.79fF
C12957 a_13432_62581# a_13973_66933# 0.30fF
C12958 ANTENNA__1197__A.DIODE _1187_.A2 4.41fF
C12959 ANTENNA__1196__A2.DIODE a_14943_26703# 0.33fF
C12960 a_18546_19530# a_50198_19938# 0.35fF
C12961 a_40250_14512# ctopn 3.58fF
C12962 VDD a_18546_68220# 32.63fF
C12963 a_13091_28327# a_10147_29415# 0.98fF
C12964 a_4075_50087# a_1674_57711# 1.76fF
C12965 pmat.rowon_n[12] pmat.rowoff_n[10] 0.31fF
C12966 a_14641_57711# pmat.row_n[6] 0.67fF
C12967 a_28131_50069# a_22199_30287# 1.41fF
C12968 VDD a_12069_38517# 8.82fF
C12969 VDD a_50290_16520# 0.56fF
C12970 a_27947_41245# a_12116_40871# 0.34fF
C12971 _1187_.A2 clk_comp 0.38fF
C12972 VDD a_6179_65479# 0.54fF
C12973 a_23933_32143# a_20616_27791# 0.45fF
C12974 pmat.row_n[15] a_2389_45859# 0.81fF
C12975 VDD a_6579_21583# 0.39fF
C12976 a_18546_59184# a_32126_59142# 0.35fF
C12977 a_29206_65166# a_29206_64162# 1.00fF
C12978 a_28202_57134# ctopp 3.57fF
C12979 VDD a_22628_30485# 1.60fF
C12980 a_27198_71190# ctopp 3.40fF
C12981 VDD a_37238_57134# 0.52fF
C12982 VDD a_36234_71190# 0.55fF
C12983 a_18546_62196# pmat.rowoff_n[6] 4.09fF
C12984 VDD a_23182_58138# 0.52fF
C12985 a_38242_23548# a_39246_23548# 0.97fF
C12986 a_12069_38517# a_14773_39394# 2.35fF
C12987 a_33222_71190# m2_32992_72014# 1.00fF
C12988 a_12993_66415# a_10921_64786# 0.76fF
C12989 pmat.row_n[4] a_2007_25597# 0.98fF
C12990 a_40250_9492# a_41254_9492# 0.97fF
C12991 cgen.dlycontrol4_in[3] a_2743_28853# 0.52fF
C12992 VDD a_36167_38825# 0.62fF
C12993 a_12309_38659# a_22537_36911# 0.88fF
C12994 a_47278_12504# a_47278_11500# 1.00fF
C12995 a_20170_11500# a_21174_11500# 0.97fF
C12996 VDD a_39469_38053# 1.26fF
C12997 VDD a_2411_33749# 4.86fF
C12998 a_18243_28327# a_10883_3303# 3.26fF
C12999 a_18546_55168# a_48190_55126# 0.35fF
C13000 a_18546_24550# a_37146_24958# 0.35fF
C13001 a_17842_27497# a_7415_29397# 0.61fF
C13002 VDD a_12228_39605# 3.84fF
C13003 a_15667_27239# a_12053_27497# 2.31fF
C13004 a_13459_28111# nmat.col_n[9] 0.91fF
C13005 nmat.col[15] a_40837_46261# 0.64fF
C13006 a_39246_61150# vcm 0.62fF
C13007 a_18546_22542# a_34134_22950# 0.35fF
C13008 a_49286_21540# ctopn 3.57fF
C13009 VDD a_2659_35015# 2.83fF
C13010 VDD a_7387_16367# 0.40fF
C13011 a_11497_40719# a_12116_40871# 0.37fF
C13012 pmat.col_n[24] pmat.col[24] 0.78fF
C13013 VDD m2_37008_54946# 0.61fF
C13014 VDD a_45943_47375# 0.43fF
C13015 VDD a_12895_53359# 0.87fF
C13016 a_33222_20536# vcm 0.65fF
C13017 pmat.row_n[7] nmat.rowon_n[7] 4.53fF
C13018 VDD a_48282_22544# 0.52fF
C13019 a_30210_65166# a_31214_65166# 0.97fF
C13020 VDD a_40903_32375# 0.33fF
C13021 VDD a_9195_7423# 0.40fF
C13022 VDD a_24186_59142# 0.52fF
C13023 pmat.col_n[14] ctopp 2.02fF
C13024 a_37238_21540# a_38242_21540# 0.97fF
C13025 VDD a_23479_35831# 0.66fF
C13026 a_44870_48437# a_44774_48695# 0.38fF
C13027 nmat.rowon_n[6] ctopn 1.40fF
C13028 VDD a_40158_72194# 0.32fF
C13029 a_41731_49525# a_45866_38279# 0.84fF
C13030 a_3866_57399# a_4025_54965# 0.92fF
C13031 a_7693_22365# a_11159_23145# 0.45fF
C13032 a_11067_27239# ANTENNA__1395__A2.DIODE 0.63fF
C13033 nmat.en_bit_n[1] _1194_.B1 1.08fF
C13034 a_45270_17524# vcm 0.65fF
C13035 a_6283_31591# a_5687_38279# 0.54fF
C13036 a_14839_20871# a_9528_20407# 0.40fF
C13037 a_18546_16518# a_19074_16926# 0.35fF
C13038 ANTENNA__1197__B.DIODE a_44389_40553# 0.59fF
C13039 _1196_.B1 a_12463_22351# 0.64fF
C13040 a_38242_71190# a_38242_70186# 1.00fF
C13041 a_46274_8488# vcm 0.64fF
C13042 a_17139_30503# a_10147_29415# 0.81fF
C13043 VDD _1519_.A 1.77fF
C13044 a_20438_35431# a_15049_36374# 1.27fF
C13045 VDD a_24667_43177# 0.55fF
C13046 a_18546_14510# a_21082_14918# 0.35fF
C13047 m2_28976_7214# m2_29980_7214# 0.96fF
C13048 a_7717_14735# a_25575_31055# 1.93fF
C13049 VDD a_12437_28585# 1.38fF
C13050 a_18546_64204# a_18162_64202# 2.62fF
C13051 pmat.rowoff_n[12] config_2_in[10] 0.87fF
C13052 VDD a_23021_29199# 1.81fF
C13053 a_35312_31599# a_44382_40847# 1.26fF
C13054 a_33467_46261# a_35186_47375# 0.47fF
C13055 a_36234_13508# a_37238_13508# 0.97fF
C13056 a_6292_65479# a_5595_65301# 0.82fF
C13057 a_22178_15516# vcm 0.65fF
C13058 VDD a_6787_47607# 11.71fF
C13059 a_18546_18526# a_51202_18934# 0.35fF
C13060 a_34226_18528# a_35230_18528# 0.97fF
C13061 ANTENNA__1197__B.DIODE a_28915_50959# 0.42fF
C13062 VDD a_2847_36799# 0.40fF
C13063 pmat.row_n[3] a_16800_47213# 1.20fF
C13064 a_12116_39783# a_11681_35823# 1.98fF
C13065 a_21174_62154# a_21174_61150# 1.00fF
C13066 a_41254_12504# vcm 0.65fF
C13067 a_46274_64162# ctopp 3.58fF
C13068 VDD a_4509_62037# 0.38fF
C13069 a_1683_45205# a_1849_45205# 0.75fF
C13070 a_19166_58138# ctopp 3.42fF
C13071 VDD a_24186_19532# 0.52fF
C13072 m2_30984_54946# m3_31116_55078# 2.79fF
C13073 VDD m2_22952_72014# 1.33fF
C13074 pmat.en_bit_n[2] clk_ena 2.62fF
C13075 a_3688_17179# clk_dig 0.31fF
C13076 VDD a_23182_10496# 0.52fF
C13077 a_29937_31055# a_2007_25597# 0.89fF
C13078 a_36234_20536# ctopn 3.58fF
C13079 a_6451_67655# a_13349_72405# 0.58fF
C13080 a_5521_72373# a_5257_69679# 0.32fF
C13081 a_11435_58791# a_4976_16091# 1.27fF
C13082 pmat.col[13] ctopp 1.97fF
C13083 a_45270_15516# a_46274_15516# 0.97fF
C13084 a_21174_15516# a_21174_14512# 1.00fF
C13085 a_18546_58180# a_30118_58138# 0.35fF
C13086 a_44266_69182# a_45270_69182# 0.97fF
C13087 a_23182_69182# a_23182_68178# 1.00fF
C13088 ANTENNA__1187__B1.DIODE nmat.col[21] 0.44fF
C13089 VDD a_77980_38962# 0.32fF
C13090 VDD pmat.row_n[2] 18.18fF
C13091 a_18546_10494# a_30118_10902# 0.35fF
C13092 VDD a_19166_57134# 0.56fF
C13093 _1196_.B1 ANTENNA__1395__A1.DIODE 0.58fF
C13094 a_31214_21540# a_31214_20536# 1.00fF
C13095 VDD a_13529_34951# 1.01fF
C13096 ANTENNA__1197__A.DIODE pmat.col[4] 0.32fF
C13097 ANTENNA__1197__B.DIODE ANTENNA__1395__B1.DIODE 3.56fF
C13098 ANTENNA__1187__B1.DIODE ANTENNA__1195__A1.DIODE 18.22fF
C13099 a_24591_28327# a_13459_28111# 0.33fF
C13100 a_48282_17524# ctopn 3.58fF
C13101 pmat.rowoff_n[4] a_9963_13967# 0.84fF
C13102 a_30210_62154# ctopp 3.58fF
C13103 VDD a_39246_62154# 0.52fF
C13104 a_24186_16520# vcm 0.65fF
C13105 cgen.dlycontrol4_in[3] cgen.start_conv_in 0.52fF
C13106 m2_46044_24282# vcm 0.42fF
C13107 a_49286_8488# ctopn 3.39fF
C13108 pmat.row_n[6] ANTENNA__1395__B1.DIODE 0.46fF
C13109 a_25695_28111# nmat.en_bit_n[0] 0.42fF
C13110 ANTENNA__1196__A2.DIODE a_35312_31599# 0.37fF
C13111 VDD a_5654_9527# 1.54fF
C13112 pmat.rowon_n[8] nmat.rowoff_n[9] 0.38fF
C13113 nmat.col_n[21] nmat.col_n[18] 9.10fF
C13114 a_49286_65166# ctopp 3.57fF
C13115 a_18546_55168# a_31122_55126# 0.35fF
C13116 a_32957_30287# a_10147_29415# 0.57fF
C13117 a_1781_9308# a_1979_12342# 0.31fF
C13118 pmat.row_n[12] pmat.row_n[3] 0.55fF
C13119 VDD nmat.col_n[4] 5.23fF
C13120 a_29206_70186# ctopp 3.57fF
C13121 a_5363_33551# clk_ena 0.34fF
C13122 VDD a_2163_53057# 0.48fF
C13123 a_19541_28879# a_18083_47593# 0.36fF
C13124 VDD a_38242_70186# 0.52fF
C13125 a_25190_15516# ctopn 3.58fF
C13126 VDD a_25190_11500# 0.52fF
C13127 a_42258_23548# a_42258_22544# 1.00fF
C13128 ANTENNA__1190__A1.DIODE nmat.col[15] 0.54fF
C13129 a_6007_42479# a_6173_42479# 0.66fF
C13130 _1154_.A ANTENNA__1190__A1.DIODE 0.39fF
C13131 pmat.col_n[12] pmat.col[12] 1.44fF
C13132 VDD nmat.col_n[13] 11.87fF
C13133 m2_17932_12234# m2_17932_11230# 0.99fF
C13134 VDD m2_17932_55950# 1.02fF
C13135 a_41254_60146# a_42258_60146# 0.97fF
C13136 a_43720_32143# a_44444_32233# 0.72fF
C13137 m2_45040_72014# m3_45172_72146# 2.79fF
C13138 a_44266_12504# ctopn 3.58fF
C13139 a_18546_69224# a_25098_69182# 0.35fF
C13140 VDD nmat.rowoff_n[6] 4.16fF
C13141 a_22537_36911# cgen.dlycontrol1_in[4] 0.50fF
C13142 a_25190_11500# a_25190_10496# 1.00fF
C13143 a_40250_56130# vcm 0.62fF
C13144 a_8491_47911# a_9405_66627# 0.43fF
C13145 VDD pmat.col_n[7] 5.54fF
C13146 a_10239_14183# a_4843_54826# 1.40fF
C13147 a_11435_58791# a_6283_31591# 0.31fF
C13148 VDD a_2467_18517# 0.50fF
C13149 a_18546_63200# a_44174_63158# 0.35fF
C13150 a_1591_15829# a_1757_15829# 0.55fF
C13151 nmat.col_n[31] nmat.col_n[30] 1.71fF
C13152 a_10883_3303# a_11948_49783# 0.67fF
C13153 a_49286_68178# a_49286_67174# 1.00fF
C13154 a_4351_55527# pmat.row_n[7] 0.56fF
C13155 a_22178_22544# vcm 0.65fF
C13156 a_30210_61150# a_31214_61150# 0.97fF
C13157 a_20170_68178# ctopp 3.57fF
C13158 a_43262_66170# vcm 0.62fF
C13159 VDD a_29206_68178# 0.52fF
C13160 a_18162_72234# vcm 7.34fF
C13161 a_18162_19532# ctopn 1.49fF
C13162 VDD a_24833_40719# 2.94fF
C13163 ANTENNA__1190__B1.DIODE a_29937_31055# 1.49fF
C13164 VDD a_4319_15039# 0.44fF
C13165 pmat.rowon_n[3] a_2389_45859# 0.35fF
C13166 a_36234_63158# vcm 0.62fF
C13167 VDD a_8443_20719# 2.99fF
C13168 VDD a_18162_21540# 2.74fF
C13169 a_7658_71543# a_7663_71317# 0.32fF
C13170 VDD inp_analog 5.75fF
C13171 pmat.col[23] ctopp 1.97fF
C13172 VDD a_4167_30511# 0.43fF
C13173 a_6292_69831# a_2149_45717# 0.47fF
C13174 a_13459_28111# a_33423_47695# 0.48fF
C13175 a_24186_20536# a_25190_20536# 0.97fF
C13176 a_18546_20534# a_31122_20942# 0.35fF
C13177 a_27198_16520# ctopn 3.58fF
C13178 pmat.row_n[4] cgen.dlycontrol4_in[5] 0.52fF
C13179 nmat.col[8] vcm 5.76fF
C13180 a_47278_16520# a_48282_16520# 0.97fF
C13181 VDD a_28901_48437# 1.26fF
C13182 a_37238_67174# a_37238_66170# 1.00fF
C13183 a_23182_9492# a_23182_8488# 1.00fF
C13184 VDD a_34226_23548# 0.54fF
C13185 a_49286_61150# ctopp 3.57fF
C13186 a_5351_19913# a_6821_18543# 0.95fF
C13187 _1196_.B1 ANTENNA__1395__A2.DIODE 8.34fF
C13188 VDD a_36234_9492# 0.52fF
C13189 a_18546_11498# a_34134_11906# 0.35fF
C13190 VDD a_14600_37607# 2.39fF
C13191 a_38851_28327# nmat.col[28] 0.56fF
C13192 a_10883_3303# ANTENNA__1190__A2.DIODE 1.96fF
C13193 VDD comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top 4.45fF
C13194 VDD a_25671_40719# 0.47fF
C13195 a_36234_17524# a_37238_17524# 0.97fF
C13196 VDD a_33949_39867# 1.27fF
C13197 m2_51064_62978# vcm 0.51fF
C13198 a_10515_15055# a_4383_7093# 1.05fF
C13199 a_34226_57134# a_35230_57134# 0.97fF
C13200 nmat.col_n[16] nmat.col[16] 0.64fF
C13201 a_39246_20536# a_39246_19532# 1.00fF
C13202 pmat.sample_n pmat.row_n[2] 3.60fF
C13203 a_41254_67174# vcm 0.62fF
C13204 a_18546_71232# a_49194_71190# 0.35fF
C13205 a_33222_71190# a_34226_71190# 0.97fF
C13206 a_33423_47695# a_45432_46983# 0.30fF
C13207 ANTENNA__1190__B1.DIODE a_15667_27239# 0.66fF
C13208 a_20170_58138# a_21174_58138# 0.97fF
C13209 VDD config_1_in[5] 1.24fF
C13210 VDD a_16657_42567# 1.28fF
C13211 a_30210_14512# vcm 0.65fF
C13212 a_15049_42902# a_14497_42658# 2.48fF
C13213 ANTENNA__1187__B1.DIODE a_7415_29397# 2.25fF
C13214 a_29206_64162# vcm 0.62fF
C13215 a_13909_39605# a_13503_39069# 0.71fF
C13216 a_37238_8488# a_38242_8488# 0.97fF
C13217 pmat.row_n[8] pmat.row_n[6] 0.60fF
C13218 VDD a_16635_31573# 0.45fF
C13219 VDD a_32218_13508# 0.52fF
C13220 a_45270_14512# a_45270_13508# 1.00fF
C13221 a_25190_22544# ctopn 3.57fF
C13222 VDD a_30210_18528# 0.52fF
C13223 pmat.sw pmat.en_bit_n[2] 0.55fF
C13224 m2_42028_54946# vcm 0.42fF
C13225 a_1586_18231# a_1591_26159# 0.64fF
C13226 a_49286_57134# a_49286_56130# 1.00fF
C13227 a_20170_61150# a_20170_60146# 1.00fF
C13228 a_4339_27804# a_5351_19913# 0.81fF
C13229 a_28202_19532# a_28202_18528# 1.00fF
C13230 VDD a_14641_57711# 1.41fF
C13231 a_7521_47081# a_11067_64015# 0.75fF
C13232 a_14773_38306# a_13597_37571# 0.47fF
C13233 a_1957_43567# cgen.dlycontrol4_in[4] 0.46fF
C13234 a_5768_9527# a_2021_11043# 0.52fF
C13235 cgen.start_conv_in a_11297_36091# 0.69fF
C13236 VDD a_41254_15516# 0.52fF
C13237 a_18546_14510# a_32126_14918# 0.35fF
C13238 a_14691_27399# a_8568_26703# 1.19fF
C13239 a_13091_52047# a_11067_30287# 1.69fF
C13240 pmat.row_n[2] pmat.rowoff_n[1] 0.34fF
C13241 a_18546_64204# a_30118_64162# 0.35fF
C13242 ANTENNA__1187__B1.DIODE pmat.col[21] 0.73fF
C13243 a_21174_59142# a_21174_58138# 1.00fF
C13244 a_5823_40303# a_5989_40303# 0.63fF
C13245 a_23182_8488# m2_22952_7214# 1.00fF
C13246 VDD m2_49056_7214# 0.91fF
C13247 pmat.col_n[1] _1179_.X 1.32fF
C13248 VDD a_17559_51157# 0.35fF
C13249 a_32218_65166# vcm 0.62fF
C13250 _1196_.B1 ANTENNA__1196__A2.DIODE 14.99fF
C13251 a_39246_21540# vcm 0.65fF
C13252 a_28202_60146# ctopp 3.58fF
C13253 a_3615_71631# pmat.rowon_n[8] 2.12fF
C13254 VDD a_45287_33231# 0.38fF
C13255 VDD a_18546_8486# 32.69fF
C13256 VDD a_37238_60146# 0.52fF
C13257 a_32405_32463# a_37637_32149# 0.60fF
C13258 a_19166_21540# a_20170_21540# 0.97fF
C13259 a_10515_61839# nmat.rowoff_n[1] 1.22fF
C13260 pmat.rowoff_n[10] ctopp 0.60fF
C13261 nmat.col_n[6] m2_24960_24282# 0.37fF
C13262 a_26194_17524# a_26194_16520# 1.00fF
C13263 a_18546_19530# a_43170_19938# 0.35fF
C13264 m2_29980_54946# m2_30984_54946# 0.96fF
C13265 a_33222_14512# ctopn 3.58fF
C13266 VDD a_4075_68583# 2.94fF
C13267 a_32218_12504# a_33222_12504# 0.97fF
C13268 a_18546_12502# a_47186_12910# 0.35fF
C13269 a_8491_47911# a_5363_70543# 0.38fF
C13270 nmat.en_bit_n[1] nmat.col_n[7] 1.26fF
C13271 a_45270_22544# a_46274_22544# 0.97fF
C13272 VDD a_43262_16520# 0.52fF
C13273 a_7717_14735# a_28704_29568# 0.57fF
C13274 a_21174_59142# a_22178_59142# 0.97fF
C13275 a_18546_59184# a_25098_59142# 0.35fF
C13276 a_10883_3303# nmat.col_n[1] 4.33fF
C13277 VDD a_33130_55126# 0.42fF
C13278 a_21174_57134# ctopp 3.57fF
C13279 a_20170_71190# ctopp 3.39fF
C13280 VDD a_30210_57134# 0.52fF
C13281 a_46274_69182# vcm 0.62fF
C13282 VDD a_29206_71190# 0.55fF
C13283 nmat.col[13] ctopn 1.97fF
C13284 pmat.sw a_4068_25615# 1.34fF
C13285 pmat.sw a_28336_29967# 0.84fF
C13286 VDD a_45238_49007# 0.48fF
C13287 a_10239_14183# nmat.rowon_n[13] 0.71fF
C13288 a_11435_58791# pmat.rowon_n[3] 0.45fF
C13289 a_11067_16359# a_9963_13967# 0.40fF
C13290 VDD a_17536_38567# 1.03fF
C13291 VDD a_44389_40553# 1.10fF
C13292 VDD a_22725_38053# 1.36fF
C13293 a_34942_51701# a_28131_50069# 0.56fF
C13294 nmat.col_n[18] clk_ena 0.53fF
C13295 a_2791_57703# pmat.rowoff_n[7] 0.94fF
C13296 a_18546_55168# a_41162_55126# 0.35fF
C13297 a_18546_24550# a_30118_24958# 0.35fF
C13298 a_10515_15055# a_4259_31375# 4.59fF
C13299 nmat.col[24] nmat.col_n[24] 1.42fF
C13300 a_11711_58261# a_11877_58261# 0.69fF
C13301 a_50290_56130# ctopp 3.37fF
C13302 a_42258_8488# m2_42028_7214# 1.00fF
C13303 a_32218_61150# vcm 0.62fF
C13304 a_16311_28327# a_18597_31599# 0.45fF
C13305 a_18546_22542# a_27106_22950# 0.35fF
C13306 a_42258_21540# ctopn 3.58fF
C13307 VDD a_2939_45503# 0.68fF
C13308 a_4707_32156# a_7939_31591# 1.33fF
C13309 a_26194_20536# vcm 0.65fF
C13310 VDD a_6799_75637# 1.26fF
C13311 VDD a_41254_22544# 0.52fF
C13312 VDD a_6927_30503# 8.01fF
C13313 nmat.col_n[27] ctopn 2.02fF
C13314 a_2199_13887# a_3413_6037# 0.36fF
C13315 VDD a_5227_13077# 0.31fF
C13316 a_46274_63158# ctopp 3.58fF
C13317 VDD a_28915_50959# 12.29fF
C13318 a_38242_17524# vcm 0.65fF
C13319 a_12309_38659# a_11113_38659# 1.37fF
C13320 VDD a_3325_20175# 1.58fF
C13321 a_11067_64015# a_6467_29415# 1.29fF
C13322 m2_26968_24282# m2_27972_24282# 0.96fF
C13323 a_39246_8488# vcm 0.64fF
C13324 nmat.rowon_n[12] a_13091_7655# 3.60fF
C13325 pmat.col_n[9] vcm 2.80fF
C13326 a_6787_47607# a_10595_53361# 1.95fF
C13327 VDD a_7263_42453# 0.45fF
C13328 nmat.col[28] nmat.col_n[19] 2.78fF
C13329 a_14149_39747# a_10767_39087# 1.96fF
C13330 pmat.row_n[15] pmat.row_n[9] 0.50fF
C13331 m2_21948_7214# m2_22952_7214# 0.96fF
C13332 a_9441_20189# a_9528_20407# 1.82fF
C13333 a_4409_74183# a_5257_69679# 0.35fF
C13334 a_48282_18528# a_48282_17524# 1.00fF
C13335 a_11921_35286# a_17996_35303# 0.42fF
C13336 VDD a_5402_56079# 0.32fF
C13337 ANTENNA__1187__B1.DIODE nmat.col_n[28] 0.48fF
C13338 a_18546_13506# a_48190_13914# 0.35fF
C13339 VDD ANTENNA__1395__B1.DIODE 17.82fF
C13340 a_11067_27239# a_2007_25597# 0.67fF
C13341 a_48282_63158# a_48282_62154# 1.00fF
C13342 a_18546_18526# a_44174_18934# 0.35fF
C13343 pmat.row_n[7] a_2952_25045# 0.47fF
C13344 a_24186_70186# a_24186_69182# 1.00fF
C13345 VDD a_19166_60146# 0.56fF
C13346 a_4075_50087# a_7435_68021# 0.49fF
C13347 VDD a_37739_37737# 0.62fF
C13348 a_34226_12504# vcm 0.65fF
C13349 a_39246_64162# ctopp 3.58fF
C13350 a_7415_29397# a_2952_25045# 0.73fF
C13351 VDD a_49286_14512# 0.52fF
C13352 a_2199_13887# a_5579_12394# 1.04fF
C13353 pmat.sample vcm 12.60fF
C13354 VDD a_48282_64162# 0.52fF
C13355 nmat.col_n[5] nmat.col[6] 6.77fF
C13356 nmat.col_n[25] nmat.col[26] 6.92fF
C13357 a_21174_19532# a_22178_19532# 0.97fF
C13358 pmat.row_n[15] pmat.rowon_n[13] 0.49fF
C13359 a_2389_45859# a_4128_46983# 0.68fF
C13360 VDD a_4611_9839# 0.51fF
C13361 a_47278_13508# a_47278_12504# 1.00fF
C13362 a_29206_20536# ctopn 3.58fF
C13363 VDD a_36854_44527# 0.31fF
C13364 pmat.rowoff_n[3] ctopp 0.60fF
C13365 VDD a_8568_26703# 1.70fF
C13366 a_2046_30184# a_7717_14735# 0.67fF
C13367 a_18546_58180# a_23090_58138# 0.35fF
C13368 pmat.col_n[6] pmat.col[6] 0.77fF
C13369 cgen.dlycontrol2_in[0] cgen.dlycontrol1_in[3] 0.46fF
C13370 a_18546_10494# a_23090_10902# 0.35fF
C13371 VDD a_12613_57141# 0.78fF
C13372 a_41254_17524# ctopn 3.58fF
C13373 nmat.col[24] ctopn 1.99fF
C13374 a_23182_62154# ctopp 3.58fF
C13375 pmat.col_n[9] pmat.col[10] 6.41fF
C13376 a_25879_31591# nmat.col[11] 0.52fF
C13377 VDD a_32218_62154# 0.52fF
C13378 a_2007_25597# a_3387_22869# 0.73fF
C13379 a_42258_8488# ctopn 3.40fF
C13380 m2_51064_21270# m3_51196_21402# 2.76fF
C13381 a_19166_67174# a_19166_66170# 1.00fF
C13382 a_22153_37179# cgen.dlycontrol2_in[0] 2.80fF
C13383 a_31214_56130# a_32218_56130# 0.97fF
C13384 a_18546_56172# a_45178_56130# 0.35fF
C13385 VDD a_44174_24958# 0.44fF
C13386 a_1591_18005# a_1757_18005# 0.47fF
C13387 a_13459_28111# nmat.col_n[6] 0.33fF
C13388 _1192_.A2 nmat.col_n[26] 4.20fF
C13389 ANTENNA__1395__A2.DIODE a_45019_38645# 0.39fF
C13390 nmat.rowon_n[13] ctopn 1.40fF
C13391 a_42258_65166# ctopp 3.58fF
C13392 VDD a_10873_40693# 6.00fF
C13393 ANTENNA__1197__B.DIODE _1192_.B1 1.13fF
C13394 a_18546_55168# a_24094_55126# 0.35fF
C13395 a_1674_68047# a_1591_67503# 0.32fF
C13396 a_18546_17522# a_19074_17930# 0.35fF
C13397 m2_17932_65990# vcm 0.44fF
C13398 a_2648_29397# a_5131_13255# 0.43fF
C13399 a_35230_24552# vcm 0.62fF
C13400 a_22178_70186# ctopp 3.57fF
C13401 a_3615_71631# a_12152_66415# 0.43fF
C13402 VDD a_31214_70186# 0.52fF
C13403 a_1923_31743# clk_dig 0.54fF
C13404 a_1586_33927# a_4149_41941# 0.37fF
C13405 pmat.row_n[4] a_12263_50959# 0.36fF
C13406 pmat.sample_n a_28915_50959# 0.48fF
C13407 a_18546_15514# a_18162_15516# 2.61fF
C13408 a_36234_62154# a_37238_62154# 0.97fF
C13409 a_43262_16520# a_43262_15516# 1.00fF
C13410 ANTENNA__1190__B1.DIODE a_11067_27239# 0.78fF
C13411 _1187_.A2 ANTENNA__1184__B1.DIODE 4.71fF
C13412 a_34226_66170# a_35230_66170# 0.97fF
C13413 pmat.rowon_n[0] ctopn 0.42fF
C13414 pmat.row_n[3] a_18546_59184# 0.35fF
C13415 nmat.col_n[7] nmat.col[8] 6.65fF
C13416 a_37238_12504# ctopn 3.58fF
C13417 _1194_.A2 a_10883_3303# 1.99fF
C13418 ANTENNA__1197__A.DIODE a_25695_28111# 0.49fF
C13419 a_33222_56130# vcm 0.62fF
C13420 _1192_.B1 a_31675_47695# 1.29fF
C13421 VDD a_20078_72194# 0.32fF
C13422 pmat.sw nmat.col_n[18] 0.32fF
C13423 nmat.en_bit_n[0] comp_latch 4.18fF
C13424 a_20170_17524# vcm 0.65fF
C13425 pmat.col[21] m2_40020_54946# 0.39fF
C13426 nmat.sample_n a_9528_20407# 0.97fF
C13427 a_27198_63158# a_28202_63158# 0.97fF
C13428 a_18546_63200# a_37146_63158# 0.35fF
C13429 m2_26968_24282# m3_27100_24414# 2.79fF
C13430 a_2411_43301# a_7847_56085# 0.40fF
C13431 a_13479_26935# a_13145_26935# 0.56fF
C13432 a_36234_66170# vcm 0.62fF
C13433 VDD a_22178_68178# 0.52fF
C13434 a_5363_12015# a_5223_11079# 0.31fF
C13435 a_8583_29199# nmat.col_n[13] 0.52fF
C13436 m2_46044_72014# m2_47048_72014# 0.96fF
C13437 a_29206_63158# vcm 0.62fF
C13438 VDD pmat.row_n[8] 33.06fF
C13439 a_26479_32117# a_39939_29967# 0.47fF
C13440 nmat.rowoff_n[6] a_8583_29199# 0.69fF
C13441 VDD a_12437_28879# 4.08fF
C13442 a_34226_55126# ctopp 1.01fF
C13443 pmat.rowon_n[7] pmat.rowoff_n[10] 0.37fF
C13444 a_18243_28327# ANTENNA__1195__A1.DIODE 0.71fF
C13445 VDD a_43170_55126# 0.42fF
C13446 a_19166_63158# pmat.col[0] 0.31fF
C13447 a_18546_20534# a_24094_20942# 0.35fF
C13448 a_6283_31591# a_19541_28879# 2.10fF
C13449 VDD pmat.rowoff_n[15] 19.62fF
C13450 a_10515_13967# a_14887_46377# 2.09fF
C13451 nmat.col_n[22] ctopn 2.02fF
C13452 a_10286_60405# a_10190_60663# 1.05fF
C13453 VDD nmat.col[5] 4.31fF
C13454 VDD a_30111_47911# 15.31fF
C13455 a_19166_9492# a_19166_8488# 1.00fF
C13456 VDD a_27198_23548# 0.55fF
C13457 a_11435_58791# a_5363_33551# 0.58fF
C13458 a_42258_61150# ctopp 3.58fF
C13459 ANTENNA__1196__A2.DIODE a_45019_38645# 2.29fF
C13460 a_35230_70186# a_36234_70186# 0.97fF
C13461 VDD a_29206_9492# 0.52fF
C13462 a_22178_11500# a_23182_11500# 0.97fF
C13463 a_18546_11498# a_27106_11906# 0.35fF
C13464 VDD a_13357_37429# 3.17fF
C13465 ANTENNA__1190__A2.DIODE a_9668_10651# 0.64fF
C13466 a_8583_29199# a_8443_20719# 0.66fF
C13467 m2_19940_7214# m3_20072_7346# 2.79fF
C13468 VDD a_45270_20536# 0.52fF
C13469 a_24186_64162# a_24186_63158# 1.00fF
C13470 a_18546_23546# vcm 0.41fF
C13471 a_27198_10496# a_27198_9492# 1.00fF
C13472 cgen.dlycontrol1_in[2] cgen.dlycontrol1_in[3] 1.23fF
C13473 a_4516_21531# clk_dig 0.97fF
C13474 a_34226_67174# vcm 0.62fF
C13475 a_18546_71232# a_42166_71190# 0.35fF
C13476 VDD a_18162_69222# 2.75fF
C13477 a_24186_58138# a_24186_57134# 1.00fF
C13478 ANTENNA__1195__A1.DIODE a_28704_29568# 0.53fF
C13479 a_40837_46261# a_45866_38279# 0.78fF
C13480 a_11067_27239# a_7109_29423# 1.84fF
C13481 a_4075_50087# a_5081_53135# 0.46fF
C13482 a_24867_53135# a_21739_29415# 0.33fF
C13483 a_23182_14512# vcm 0.65fF
C13484 nmat.col_n[3] nmat.col[4] 6.61fF
C13485 a_22178_64162# vcm 0.62fF
C13486 a_18546_8486# a_50198_8894# 0.35fF
C13487 a_28202_60146# a_28202_59142# 1.00fF
C13488 a_18546_65208# a_47186_65166# 0.35fF
C13489 a_18162_59182# ctopp 1.49fF
C13490 pmat.col_n[17] ctopp 2.01fF
C13491 VDD a_35799_35831# 0.61fF
C13492 VDD a_43170_72194# 0.33fF
C13493 a_46274_62154# a_46274_61150# 1.00fF
C13494 VDD a_25190_13508# 0.52fF
C13495 a_30699_29397# a_19405_28853# 0.76fF
C13496 a_2791_57703# a_1591_61519# 0.42fF
C13497 cgen.dlycontrol4_in[5] cgen.dlycontrol4_in[1] 4.35fF
C13498 VDD a_23182_18528# 0.52fF
C13499 a_29206_63158# pmat.col[10] 0.31fF
C13500 VDD m2_51064_67998# 1.06fF
C13501 a_32218_67174# a_33222_67174# 0.97fF
C13502 a_18546_67216# a_47186_67174# 0.35fF
C13503 a_18546_9490# a_20078_9898# 0.35fF
C13504 a_26155_46831# a_26321_46831# 0.39fF
C13505 nmat.col[23] m2_42028_24282# 0.39fF
C13506 a_29206_66170# a_29206_65166# 1.00fF
C13507 a_22178_22544# a_22178_21540# 1.00fF
C13508 VDD a_36617_43131# 1.33fF
C13509 VDD a_34226_15516# 0.52fF
C13510 a_18546_14510# a_25098_14918# 0.35fF
C13511 a_21174_14512# a_22178_14512# 0.97fF
C13512 a_46274_15516# a_46274_14512# 1.00fF
C13513 a_14653_53458# a_11067_30287# 0.54fF
C13514 VDD a_18795_28882# 0.39fF
C13515 a_15667_27239# nmat.col[26] 0.88fF
C13516 a_18546_7482# a_47186_7890# 0.35fF
C13517 a_20170_64162# a_21174_64162# 0.97fF
C13518 a_18546_64204# a_23090_64162# 0.35fF
C13519 a_4399_51157# a_2983_48071# 0.67fF
C13520 a_48282_69182# a_48282_68178# 1.00fF
C13521 a_26194_68178# a_27198_68178# 0.97fF
C13522 pmat.rowoff_n[14] ctopp 0.60fF
C13523 ANTENNA__1197__B.DIODE a_43720_32143# 0.45fF
C13524 VDD a_10864_68565# 0.87fF
C13525 VDD a_2493_11477# 0.62fF
C13526 a_11892_21959# a_8305_20871# 0.33fF
C13527 VDD m2_35000_7214# 1.30fF
C13528 VDD a_6979_51157# 1.07fF
C13529 _1183_.A2 nmat.col_n[30] 2.66fF
C13530 a_25190_65166# vcm 0.62fF
C13531 VDD a_15899_47939# 4.09fF
C13532 a_32218_21540# vcm 0.65fF
C13533 a_21174_60146# ctopp 3.58fF
C13534 a_5363_70543# a_3923_68021# 1.59fF
C13535 VDD a_44533_33749# 1.35fF
C13536 VDD a_12815_8213# 0.48fF
C13537 VDD a_30210_60146# 0.52fF
C13538 ANTENNA__1395__A1.DIODE a_22199_30287# 1.07fF
C13539 VDD a_12934_35823# 1.06fF
C13540 a_47278_58138# vcm 0.62fF
C13541 a_20475_49783# a_13643_29415# 0.46fF
C13542 a_18546_63200# a_18162_63198# 2.62fF
C13543 m2_37008_54946# m3_37140_55078# 2.79fF
C13544 ANTENNA__1195__A1.DIODE a_18547_51565# 0.40fF
C13545 a_18546_19530# a_36142_19938# 0.35fF
C13546 m2_22952_54946# m2_23956_54946# 0.96fF
C13547 a_18546_66212# vcm 0.40fF
C13548 a_26194_14512# ctopn 3.58fF
C13549 pmat.en_bit_n[0] _1179_.X 0.64fF
C13550 a_18546_12502# a_40158_12910# 0.35fF
C13551 a_50290_12504# m2_51064_12234# 0.96fF
C13552 VDD a_14773_43746# 1.34fF
C13553 VDD a_36234_16520# 0.52fF
C13554 pmat.col[22] ctopp 1.97fF
C13555 pmat.col_n[13] m2_31988_54946# 0.38fF
C13556 VDD m2_17932_22274# 1.01fF
C13557 VDD a_9463_50877# 0.96fF
C13558 nmat.rowon_n[4] vcm 0.54fF
C13559 a_22178_65166# a_22178_64162# 1.00fF
C13560 a_30571_50959# a_38391_47381# 0.62fF
C13561 VDD a_26102_55126# 0.42fF
C13562 VDD a_46182_7890# 0.33fF
C13563 a_50290_11500# a_50290_10496# 1.00fF
C13564 VDD a_23182_57134# 0.52fF
C13565 _1196_.B1 ANTENNA__1190__B1.DIODE 0.56fF
C13566 a_39246_69182# vcm 0.62fF
C13567 VDD a_22178_71190# 0.55fF
C13568 a_18546_23546# a_45178_23954# 0.35fF
C13569 a_31214_23548# a_32218_23548# 0.97fF
C13570 a_38851_28327# nmat.col[31] 2.16fF
C13571 a_18546_9490# a_49194_9898# 0.35fF
C13572 a_33222_9492# a_34226_9492# 0.97fF
C13573 pmat.rowoff_n[7] a_1769_13103# 0.90fF
C13574 a_19166_58138# a_20170_58138# 0.97fF
C13575 VDD a_6412_8725# 0.38fF
C13576 a_48282_59142# vcm 0.62fF
C13577 VDD a_17441_40482# 1.25fF
C13578 a_40250_12504# a_40250_11500# 1.00fF
C13579 a_34204_27765# nmat.col_n[30] 1.20fF
C13580 ANTENNA__1190__A1.DIODE nmat.col[8] 0.45fF
C13581 pmat.rowon_n[0] a_4257_34319# 2.41fF
C13582 a_9217_23983# a_8013_25615# 0.58fF
C13583 VDD a_8656_63811# 0.65fF
C13584 VDD config_2_in[3] 1.19fF
C13585 a_18546_24550# a_23090_24958# 0.35fF
C13586 a_28704_29568# a_7415_29397# 1.12fF
C13587 a_20170_24552# ctopn 0.57fF
C13588 nmat.col[29] nmat.col_n[29] 1.06fF
C13589 ANTENNA__1190__B1.DIODE a_9785_28879# 1.73fF
C13590 a_7658_71543# a_1674_57711# 0.91fF
C13591 _1187_.A2 pmat.col[23] 0.47fF
C13592 a_43262_56130# ctopp 3.40fF
C13593 VDD nmat.col[18] 10.17fF
C13594 a_49286_20536# a_50290_20536# 0.97fF
C13595 ANTENNA__1196__A2.DIODE nmat.sw 1.27fF
C13596 a_25190_61150# vcm 0.62fF
C13597 a_6283_31591# a_33869_31599# 0.39fF
C13598 a_35230_21540# ctopn 3.58fF
C13599 pmat.row_n[2] a_18359_49140# 0.64fF
C13600 a_18162_20536# vcm 6.95fF
C13601 a_48282_9492# a_48282_8488# 1.00fF
C13602 a_23182_65166# a_24186_65166# 0.97fF
C13603 VDD a_34226_22544# 0.52fF
C13604 a_46274_66170# ctopp 3.58fF
C13605 m2_50060_72014# m3_50192_72146# 2.79fF
C13606 pmat.rowon_n[8] a_2046_30184# 1.08fF
C13607 a_30210_21540# a_31214_21540# 0.97fF
C13608 VDD a_34611_36649# 0.64fF
C13609 VDD pmat.col_n[10] 5.17fF
C13610 a_39246_63158# ctopp 3.58fF
C13611 VDD a_48282_63158# 0.52fF
C13612 pmat.row_n[9] nmat.rowoff_n[5] 0.54fF
C13613 a_14653_53458# _1192_.A2 0.78fF
C13614 a_31214_17524# vcm 0.65fF
C13615 a_34705_51959# a_34942_51701# 1.72fF
C13616 cgen.dlycontrol4_in[4] a_16657_42567# 0.63fF
C13617 VDD a_10975_18231# 0.41fF
C13618 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot vcm 673.52fF
C13619 a_18546_61192# a_47186_61150# 0.35fF
C13620 a_31214_71190# a_31214_70186# 1.00fF
C13621 a_32218_8488# vcm 0.64fF
C13622 a_7840_27247# a_8568_26703# 0.62fF
C13623 a_45270_58138# a_46274_58138# 0.97fF
C13624 nmat.col[21] ANTENNA__1190__A2.DIODE 7.85fF
C13625 a_2199_13887# a_1717_13647# 0.59fF
C13626 ANTENNA__1195__A1.DIODE ANTENNA__1190__A2.DIODE 0.97fF
C13627 pmat.col_n[18] pmat.col[18] 0.78fF
C13628 a_48282_19532# vcm 0.65fF
C13629 _1196_.B1 a_7109_29423# 0.34fF
C13630 nmat.rowon_n[7] a_11067_64015# 1.41fF
C13631 VDD a_9761_30511# 0.53fF
C13632 a_47278_10496# vcm 0.65fF
C13633 VDD result_out[13] 0.63fF
C13634 a_10055_31591# a_6559_33767# 0.88fF
C13635 a_18546_13506# a_41162_13914# 0.35fF
C13636 a_29206_13508# a_30210_13508# 0.97fF
C13637 a_11948_49783# a_25839_49783# 0.62fF
C13638 a_4991_69831# a_11711_50959# 0.44fF
C13639 a_2263_43719# a_5173_45993# 0.33fF
C13640 a_30663_50087# a_31675_47695# 0.80fF
C13641 a_45270_61150# a_45270_60146# 1.00fF
C13642 a_44266_67174# ctopp 3.58fF
C13643 a_18546_18526# a_37146_18934# 0.35fF
C13644 a_27198_18528# a_28202_18528# 0.97fF
C13645 VDD a_19817_37692# 1.18fF
C13646 m2_51064_67998# m2_51064_66994# 0.99fF
C13647 a_27198_12504# vcm 0.65fF
C13648 a_32218_64162# ctopp 3.58fF
C13649 VDD a_42258_14512# 0.52fF
C13650 a_13459_28111# a_19283_49783# 0.35fF
C13651 VDD a_41254_64162# 0.52fF
C13652 VDD a_39413_40956# 1.33fF
C13653 a_10055_31591# a_2215_47375# 0.63fF
C13654 VDD comp.adc_nor_latch_0.NOR_1/A 1.16fF
C13655 VDD _1192_.B1 14.44fF
C13656 a_18546_58180# vcm 0.41fF
C13657 a_46274_59142# a_46274_58138# 1.00fF
C13658 _1187_.A2 nmat.col_n[29] 1.66fF
C13659 VDD a_12705_10389# 0.33fF
C13660 ANTENNA__1395__B1.DIODE a_8583_29199# 0.32fF
C13661 ANTENNA__1184__B1.DIODE a_47212_29673# 0.36fF
C13662 a_22178_20536# ctopn 3.58fF
C13663 VDD a_23663_44535# 0.60fF
C13664 a_38242_15516# a_39246_15516# 0.97fF
C13665 VDD m2_32992_24282# 0.61fF
C13666 a_2419_53351# a_3199_53877# 0.54fF
C13667 a_2046_30184# a_9944_32259# 0.49fF
C13668 a_37238_69182# a_38242_69182# 0.97fF
C13669 nmat.col[17] a_36234_24552# 0.39fF
C13670 VDD a_23395_53135# 4.46fF
C13671 a_24186_21540# a_24186_20536# 1.00fF
C13672 a_4075_31591# a_4707_32156# 0.48fF
C13673 a_34226_17524# ctopn 3.58fF
C13674 a_33467_46261# a_13275_48783# 0.39fF
C13675 a_49286_11500# vcm 0.65fF
C13676 a_35312_31599# nmat.col_n[21] 0.93fF
C13677 pmat.row_n[6] nmat.sample 0.34fF
C13678 ANTENNA__1187__B1.DIODE a_11067_30287# 0.78fF
C13679 VDD a_25190_62154# 0.52fF
C13680 a_2051_29973# a_2217_29973# 0.41fF
C13681 a_24937_43655# a_11041_39860# 0.49fF
C13682 nmat.col_n[31] vcm 3.97fF
C13683 a_9963_28111# nmat.col_n[1] 0.92fF
C13684 a_35230_8488# ctopn 3.40fF
C13685 a_6283_31591# a_32405_32463# 0.57fF
C13686 a_18546_56172# a_38150_56130# 0.35fF
C13687 VDD a_37146_24958# 0.44fF
C13688 a_4339_27804# a_9075_28023# 0.73fF
C13689 VDD a_10195_59861# 0.40fF
C13690 a_4128_64391# a_6927_30503# 0.35fF
C13691 a_12345_39100# a_11497_38543# 0.34fF
C13692 a_35230_65166# ctopp 3.58fF
C13693 a_9963_28111# a_15667_28111# 0.38fF
C13694 a_1895_41018# a_1757_40853# 0.70fF
C13695 VDD a_44266_65166# 0.52fF
C13696 a_46274_59142# a_47278_59142# 0.97fF
C13697 a_4843_54826# a_1586_50247# 0.41fF
C13698 a_50290_10496# ctopn 3.43fF
C13699 a_18546_68220# a_46182_68178# 0.35fF
C13700 VDD a_10441_21263# 4.89fF
C13701 VDD a_24186_70186# 0.52fF
C13702 nmat.col[4] vcm 5.76fF
C13703 VDD a_5012_10927# 0.48fF
C13704 VDD a_4627_26703# 0.37fF
C13705 a_35230_23548# a_35230_22544# 1.00fF
C13706 a_1781_9308# a_1949_9308# 0.48fF
C13707 a_3339_59879# a_8841_60405# 0.40fF
C13708 a_34226_60146# a_35230_60146# 0.97fF
C13709 a_18546_60188# a_51202_60146# 0.35fF
C13710 pmat.row_n[7] a_1586_18231# 0.55fF
C13711 a_30210_12504# ctopn 3.58fF
C13712 a_7674_69135# a_4583_68021# 0.55fF
C13713 pmat.row_n[5] nmat.en_bit_n[1] 1.36fF
C13714 _1154_.X vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.65fF
C13715 a_26194_56130# vcm 0.62fF
C13716 VDD a_31425_37218# 1.20fF
C13717 VDD a_3111_53333# 0.46fF
C13718 pmat.sw a_29937_31055# 0.31fF
C13719 nmat.en_bit_n[0] ANTENNA__1183__B1.DIODE 1.43fF
C13720 a_17842_27497# a_24747_29967# 0.38fF
C13721 a_12197_38306# ndecision_finish 0.74fF
C13722 a_18546_63200# a_30118_63158# 0.35fF
C13723 a_4339_27804# a_2564_21959# 0.34fF
C13724 _1154_.A _1519_.A 0.33fF
C13725 VDD m2_17932_71010# 1.03fF
C13726 a_42258_68178# a_42258_67174# 1.00fF
C13727 a_23182_61150# a_24186_61150# 0.97fF
C13728 a_49286_69182# ctopp 3.57fF
C13729 a_7415_29397# ANTENNA__1190__A2.DIODE 1.29fF
C13730 a_29206_66170# vcm 0.62fF
C13731 VDD a_5651_66975# 8.37fF
C13732 m2_39016_72014# m2_40020_72014# 0.96fF
C13733 a_10515_13967# a_7533_19087# 0.70fF
C13734 a_22178_63158# vcm 0.62fF
C13735 VDD a_1643_65301# 0.39fF
C13736 pmat.en_bit_n[0] nmat.sample_n 1.63fF
C13737 VDD a_46027_44905# 0.73fF
C13738 VDD a_36142_55126# 0.38fF
C13739 nmat.rowon_n[7] a_4613_19087# 0.41fF
C13740 VDD a_8399_6037# 0.52fF
C13741 a_2419_53351# a_1823_58237# 2.14fF
C13742 a_20170_13508# a_21174_13508# 0.97fF
C13743 a_27603_34191# a_29159_37607# 0.49fF
C13744 VDD m2_17932_10226# 1.01fF
C13745 a_10781_42869# a_12228_40693# 1.86fF
C13746 cgen.dlycontrol4_in[0] cgen.dlycontrol4_in[2] 2.13fF
C13747 nmat.col_n[9] ctopn 2.02fF
C13748 pmat.col[0] pmat.col[8] 0.41fF
C13749 a_40250_16520# a_41254_16520# 0.97fF
C13750 a_30210_67174# a_30210_66170# 1.00fF
C13751 VDD a_26957_38779# 1.27fF
C13752 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 1285.92fF
C13753 a_35230_61150# ctopp 3.58fF
C13754 m2_17932_22274# m2_17932_21270# 0.99fF
C13755 pmat.row_n[15] pmat.rowoff_n[8] 3.59fF
C13756 VDD a_22178_9492# 0.52fF
C13757 VDD a_44266_61150# 0.52fF
C13758 a_18546_11498# a_19074_11906# 0.35fF
C13759 VDD a_31701_37462# 1.20fF
C13760 nmat.col[30] nmat.col[19] 4.52fF
C13761 a_2411_33749# a_1591_36501# 0.34fF
C13762 pmat.sw a_15667_27239# 2.78fF
C13763 VDD a_38242_20536# 0.52fF
C13764 a_29206_17524# a_30210_17524# 0.97fF
C13765 ANTENNA__1196__A2.DIODE nmat.col_n[30] 1.32fF
C13766 a_27198_57134# a_28202_57134# 0.97fF
C13767 a_22085_38550# a_22541_38779# 0.47fF
C13768 a_32218_20536# a_32218_19532# 1.00fF
C13769 a_26194_71190# a_27198_71190# 0.97fF
C13770 a_18546_71232# a_35138_71190# 0.35fF
C13771 a_27198_67174# vcm 0.62fF
C13772 m3_36136_55078# ctopp 0.36fF
C13773 _1187_.A2 a_13091_28327# 1.29fF
C13774 ANTENNA__1187__B1.DIODE _1192_.A2 0.75fF
C13775 a_10049_60663# a_9135_60967# 0.33fF
C13776 pmat.col_n[27] _1179_.X 0.39fF
C13777 VDD a_43720_32143# 5.45fF
C13778 pmat.rowoff_n[8] pmat.col[0] 0.33fF
C13779 VDD a_50290_17524# 0.54fF
C13780 pmat.col_n[7] pmat.col[7] 0.76fF
C13781 VDD a_5991_23983# 3.36fF
C13782 pmat.col_n[0] m2_18936_54946# 0.37fF
C13783 VDD m2_28976_54946# 0.62fF
C13784 a_9983_32385# a_7939_31591# 0.33fF
C13785 a_30210_8488# a_31214_8488# 0.97fF
C13786 a_18546_8486# a_43170_8894# 0.35fF
C13787 a_18546_65208# a_40158_65166# 0.35fF
C13788 _1154_.X nmat.col_n[31] 0.75fF
C13789 a_49286_70186# a_49286_69182# 1.00fF
C13790 a_13503_36893# a_15144_36165# 0.52fF
C13791 pmat.col[16] pmat.col[15] 0.48fF
C13792 a_8305_20871# a_3688_17179# 0.61fF
C13793 VDD a_15107_35831# 0.62fF
C13794 a_38242_14512# a_38242_13508# 1.00fF
C13795 VDD cgen.dlycontrol3_in[4] 9.55fF
C13796 a_11497_38543# a_12693_38543# 0.45fF
C13797 a_18546_67216# a_40158_67174# 0.35fF
C13798 a_18546_56172# a_20078_56130# 0.35fF
C13799 a_42258_57134# a_42258_56130# 1.00fF
C13800 a_21174_19532# a_21174_18528# 1.00fF
C13801 a_46274_19532# a_47278_19532# 0.97fF
C13802 a_12309_38659# a_12197_38306# 0.57fF
C13803 a_16311_28327# a_45915_29941# 0.57fF
C13804 pmat.col_n[12] vcm 2.80fF
C13805 VDD a_16355_43123# 1.44fF
C13806 VDD a_27198_15516# 0.52fF
C13807 nmat.col_n[11] nmat.col_n[29] 0.32fF
C13808 m2_51064_17254# vcm 0.50fF
C13809 nmat.rowon_n[7] a_3325_40847# 0.40fF
C13810 a_31210_31751# a_31339_31787# 0.42fF
C13811 a_18546_7482# a_40158_7890# 0.35fF
C13812 pmat.rowon_n[0] ctopp 1.34fF
C13813 a_45270_10496# a_46274_10496# 0.97fF
C13814 VDD pmat.row_n[0] 20.11fF
C13815 a_6283_31591# a_13830_47607# 0.30fF
C13816 a_4128_46983# a_19541_28879# 1.29fF
C13817 VDD a_46274_12504# 0.52fF
C13818 VDD m2_20944_7214# 0.91fF
C13819 a_18546_15514# vcm 0.41fF
C13820 a_11113_39747# cgen.dlycontrol2_in[4] 2.68fF
C13821 VDD pmat.col[14] 4.71fF
C13822 VDD a_11397_76457# 0.34fF
C13823 a_3615_71631# a_11067_30287# 1.05fF
C13824 VDD a_11547_48061# 0.45fF
C13825 nmat.rowon_n[7] a_3571_13627# 0.90fF
C13826 a_25190_21540# vcm 0.65fF
C13827 a_1591_8213# a_1757_8213# 0.75fF
C13828 VDD a_23182_60146# 0.52fF
C13829 VDD a_12345_36924# 4.24fF
C13830 a_40250_58138# vcm 0.62fF
C13831 a_18563_27791# a_34204_27765# 0.30fF
C13832 nmat.rowon_n[6] a_14457_15823# 0.68fF
C13833 a_1923_31743# a_9595_30511# 0.60fF
C13834 a_5363_70543# a_1957_43567# 0.38fF
C13835 a_11435_58791# pmat.row_n[4] 2.00fF
C13836 a_18546_19530# a_29114_19938# 0.35fF
C13837 a_18162_14512# ctopn 1.49fF
C13838 a_25190_12504# a_26194_12504# 0.97fF
C13839 a_18546_12502# a_33130_12910# 0.35fF
C13840 a_2215_47375# a_6559_33767# 1.72fF
C13841 ANTENNA__1184__B1.DIODE nmat.col[30] 1.64fF
C13842 _1187_.A2 a_17139_30503# 0.74fF
C13843 a_3339_59879# a_10811_77437# 0.34fF
C13844 a_38242_22544# a_39246_22544# 0.97fF
C13845 VDD a_10591_44265# 0.57fF
C13846 VDD a_29206_16520# 0.52fF
C13847 a_11497_40719# a_12197_41570# 0.34fF
C13848 a_10515_13967# a_12263_50959# 0.49fF
C13849 a_40837_46261# a_35244_32411# 0.58fF
C13850 pmat.col_n[9] m2_27972_54946# 0.38fF
C13851 a_4707_32156# a_14287_31599# 0.73fF
C13852 VDD a_19074_55126# 0.43fF
C13853 VDD a_39154_7890# 0.34fF
C13854 _1519_.A pmat.col[31] 5.26fF
C13855 VDD a_4831_34561# 0.40fF
C13856 a_32218_69182# vcm 0.62fF
C13857 VDD a_6087_70919# 0.52fF
C13858 a_18546_23546# a_38150_23954# 0.35fF
C13859 pmat.rowon_n[0] a_1586_50247# 0.84fF
C13860 a_18546_9490# a_42166_9898# 0.35fF
C13861 a_41254_59142# vcm 0.62fF
C13862 a_10949_43124# a_11297_36091# 1.62fF
C13863 VDD a_30663_50087# 10.45fF
C13864 _1194_.A2 ANTENNA__1195__A1.DIODE 0.71fF
C13865 vcm.sky130_fd_sc_hd__buf_4_0.X vcm.sky130_fd_sc_hd__buf_4_1.X 0.72fF
C13866 nmat.col_n[28] ANTENNA__1190__A2.DIODE 0.53fF
C13867 VDD a_20170_20536# 0.52fF
C13868 a_20170_17524# a_21174_17524# 0.97fF
C13869 a_36234_56130# ctopp 3.44fF
C13870 VDD a_22979_29967# 0.60fF
C13871 a_18546_57176# a_19074_57134# 0.35fF
C13872 pmat.rowon_n[1] a_18162_57174# 1.19fF
C13873 VDD a_45270_56130# 0.55fF
C13874 a_33467_46261# a_1781_9308# 2.34fF
C13875 a_19965_39867# a_19509_39638# 0.33fF
C13876 a_28202_21540# ctopn 3.58fF
C13877 _1196_.B1 nmat.col[26] 6.45fF
C13878 VDD a_12604_47080# 0.47fF
C13879 VDD a_27198_22544# 0.52fF
C13880 a_39246_66170# ctopp 3.58fF
C13881 VDD a_48282_66170# 0.52fF
C13882 a_47278_11500# a_48282_11500# 0.97fF
C13883 VDD a_21124_36391# 1.14fF
C13884 a_37820_30485# a_41731_49525# 1.20fF
C13885 a_32218_63158# ctopp 3.58fF
C13886 VDD a_41254_63158# 0.52fF
C13887 a_6664_26159# ANTENNA__1183__B1.DIODE 0.37fF
C13888 a_24186_17524# vcm 0.65fF
C13889 pmat.col_n[12] _1154_.X 0.37fF
C13890 pmat.row_n[11] a_3305_17999# 0.53fF
C13891 a_49286_64162# a_49286_63158# 1.00fF
C13892 m2_31988_24282# m3_32120_24414# 2.79fF
C13893 pmat.rowon_n[11] nmat.rowoff_n[3] 2.46fF
C13894 a_18162_22544# vcm 6.95fF
C13895 a_18546_61192# a_40158_61150# 0.35fF
C13896 VDD a_8307_23439# 0.57fF
C13897 m2_46044_54946# m2_47048_54946# 0.96fF
C13898 a_25190_8488# vcm 0.64fF
C13899 a_49286_58138# a_49286_57134# 1.00fF
C13900 pmat.col_n[25] pmat.col[26] 5.88fF
C13901 pmat.sample_n pmat.row_n[0] 0.40fF
C13902 a_10873_38517# a_11041_36596# 0.69fF
C13903 _1187_.A2 a_11927_27399# 0.37fF
C13904 cgen.start_conv_in a_17675_37001# 0.37fF
C13905 VDD a_28525_43655# 1.20fF
C13906 VDD a_9287_65087# 0.39fF
C13907 ANTENNA__1190__B1.DIODE nmat.sw 3.74fF
C13908 a_41254_19532# vcm 0.65fF
C13909 _1192_.A2 a_16800_47213# 0.56fF
C13910 a_41254_18528# a_41254_17524# 1.00fF
C13911 pmat.rowoff_n[4] nmat.rowon_n[12] 0.42fF
C13912 VDD a_40125_31029# 0.33fF
C13913 a_6975_76823# a_8539_76181# 0.37fF
C13914 a_6795_76989# a_9183_76359# 0.34fF
C13915 a_35230_24552# m3_35132_24990# 1.39fF
C13916 VDD nmat.sample 6.91fF
C13917 a_40250_10496# vcm 0.65fF
C13918 a_18546_13506# a_34134_13914# 0.35fF
C13919 _1183_.A2 nmat.col[1] 0.42fF
C13920 a_24937_36039# clk_dig 0.52fF
C13921 cgen.dlycontrol4_in[0] a_12228_40693# 0.34fF
C13922 a_41254_63158# a_41254_62154# 1.00fF
C13923 pmat.sw a_3622_29967# 0.35fF
C13924 a_38242_71190# m2_38012_72014# 1.00fF
C13925 a_37238_67174# ctopp 3.58fF
C13926 a_18546_18526# a_30118_18934# 0.35fF
C13927 nmat.col[10] vcm 5.77fF
C13928 VDD a_46274_67174# 0.52fF
C13929 m2_17932_18258# vcm 0.44fF
C13930 nmat.rowon_n[12] nmat.col_n[3] 0.34fF
C13931 a_9411_2215# a_4383_7093# 1.08fF
C13932 a_47278_22544# a_47278_21540# 1.00fF
C13933 a_2021_26677# a_1923_31743# 1.43fF
C13934 a_25190_64162# ctopp 3.58fF
C13935 VDD a_35230_14512# 0.52fF
C13936 a_23182_62154# pmat.col[4] 0.31fF
C13937 a_46274_14512# a_47278_14512# 0.97fF
C13938 m2_24960_7214# m3_25092_7346# 2.79fF
C13939 VDD a_34226_64162# 0.52fF
C13940 pmat.en_bit_n[2] pmat.en_bit_n[0] 12.10fF
C13941 nmat.en_bit_n[0] a_20310_28029# 0.65fF
C13942 a_45270_64162# a_46274_64162# 0.97fF
C13943 nmat.col[11] m2_29980_24282# 0.39fF
C13944 a_18546_57176# a_48190_57134# 0.35fF
C13945 a_2411_16101# a_9319_15279# 0.49fF
C13946 VDD a_51202_11906# 0.30fF
C13947 VDD a_1895_50308# 0.43fF
C13948 a_40250_13508# a_40250_12504# 1.00fF
C13949 _1187_.A2 _1184_.A2 2.93fF
C13950 VDD a_3911_44431# 0.36fF
C13951 _1194_.B1 nmat.col[10] 0.37fF
C13952 a_6283_31591# cgen.dlycontrol1_in[0] 1.11fF
C13953 a_3339_59879# a_3615_71631# 0.31fF
C13954 a_10515_15055# nmat.rowon_n[2] 0.90fF
C13955 VDD a_21082_7890# 0.33fF
C13956 pmat.col_n[20] ctopp 2.02fF
C13957 VDD a_10651_35507# 1.06fF
C13958 VDD a_46182_72194# 0.32fF
C13959 a_27198_17524# ctopn 3.58fF
C13960 a_42258_11500# vcm 0.65fF
C13961 a_50290_14512# m2_51064_14242# 0.96fF
C13962 nmat.rowoff_n[6] a_11892_21959# 0.76fF
C13963 a_28202_8488# ctopn 3.40fF
C13964 a_24186_56130# a_25190_56130# 0.97fF
C13965 a_18546_56172# a_31122_56130# 0.35fF
C13966 VDD a_30118_24958# 0.44fF
C13967 pmat.row_n[15] ctopn 1.39fF
C13968 m2_43032_24282# m2_44036_24282# 0.96fF
C13969 nmat.sw a_7109_29423# 0.94fF
C13970 a_44266_19532# ctopn 3.58fF
C13971 a_28202_65166# ctopp 3.58fF
C13972 VDD a_10781_42364# 7.99fF
C13973 a_40837_46261# a_44763_34293# 0.87fF
C13974 VDD a_37238_65166# 0.52fF
C13975 a_1761_7119# a_1761_6031# 0.47fF
C13976 VDD a_44266_21540# 0.52fF
C13977 a_47278_65166# a_47278_64162# 1.00fF
C13978 a_43262_10496# ctopn 3.58fF
C13979 a_18546_68220# a_39154_68178# 0.35fF
C13980 a_6787_47607# a_6292_65479# 0.77fF
C13981 a_10697_75218# a_12981_74581# 0.60fF
C13982 a_11225_35836# clk_ena 1.48fF
C13983 a_50290_58138# ctopp 3.43fF
C13984 a_46274_68178# vcm 0.62fF
C13985 VDD a_12719_69367# 1.38fF
C13986 VDD a_8472_11739# 1.12fF
C13987 a_18546_72236# a_23090_72194# 0.35fF
C13988 pmat.col[24] ctopp 1.97fF
C13989 ANTENNA__1395__A1.DIODE a_41731_49525# 0.37fF
C13990 _1187_.A2 a_9411_2215# 0.35fF
C13991 a_2149_45717# a_2791_57703# 2.09fF
C13992 a_6292_69831# a_3615_71631# 0.37fF
C13993 a_36234_16520# a_36234_15516# 1.00fF
C13994 a_29206_62154# a_30210_62154# 0.97fF
C13995 a_27198_66170# a_28202_66170# 0.97fF
C13996 a_18546_60188# a_44174_60146# 0.35fF
C13997 a_25879_31591# nmat.col[14] 0.33fF
C13998 a_28915_50959# nmat.col[15] 0.42fF
C13999 a_23182_12504# ctopn 3.58fF
C14000 _1154_.A a_28915_50959# 0.31fF
C14001 a_5497_62839# a_4075_68583# 3.29fF
C14002 a_2419_69455# cgen.dlycontrol4_in[2] 0.92fF
C14003 nmat.col_n[4] m2_22952_24282# 0.38fF
C14004 pmat.row_n[7] a_2411_43301# 1.32fF
C14005 a_20170_14512# a_20170_13508# 1.00fF
C14006 a_18546_63200# a_23090_63158# 0.35fF
C14007 a_20170_63158# a_21174_63158# 0.97fF
C14008 nmat.rowon_n[14] a_2683_22089# 1.31fF
C14009 m2_42028_54946# m3_42160_55078# 2.79fF
C14010 pmat.row_n[1] pmat.rowoff_n[0] 0.75fF
C14011 VDD m2_38012_72014# 1.00fF
C14012 a_9785_28879# clk_ena 2.99fF
C14013 a_42258_69182# ctopp 3.58fF
C14014 a_22178_66170# vcm 0.62fF
C14015 m2_31988_72014# m2_32992_72014# 0.96fF
C14016 VDD a_13091_18535# 3.19fF
C14017 VDD a_14491_51969# 0.41fF
C14018 a_48282_65166# a_49286_65166# 0.97fF
C14019 a_45270_11500# ctopn 3.58fF
C14020 VDD a_5535_29980# 1.53fF
C14021 ANTENNA__1190__B1.DIODE a_14947_26159# 0.53fF
C14022 VDD a_12967_58559# 0.52fF
C14023 _1154_.A ANTENNA__1395__B1.DIODE 0.99fF
C14024 VDD a_46779_35113# 0.39fF
C14025 a_21279_48999# a_33423_47695# 3.28fF
C14026 a_10239_14183# pmat.rowon_n[3] 0.53fF
C14027 a_4383_7093# a_9459_5461# 0.55fF
C14028 nmat.rowon_n[13] nmat.rowoff_n[1] 0.89fF
C14029 a_2215_47375# a_4413_62037# 0.44fF
C14030 a_19166_67174# ctopp 3.43fF
C14031 VDD a_11497_38543# 3.80fF
C14032 a_28202_61150# ctopp 3.58fF
C14033 a_30210_63158# pmat.col[11] 0.31fF
C14034 a_28202_70186# a_29206_70186# 0.97fF
C14035 VDD a_37238_61150# 0.52fF
C14036 VDD a_26423_40183# 0.63fF
C14037 a_36161_37462# a_36617_37691# 0.33fF
C14038 a_2935_38279# a_2839_38101# 1.06fF
C14039 pmat.rowon_n[1] vcm 0.62fF
C14040 VDD a_13503_37981# 2.11fF
C14041 a_49286_13508# vcm 0.65fF
C14042 VDD a_25209_42043# 1.15fF
C14043 a_4719_30287# a_13091_18535# 2.85fF
C14044 nmat.col[24] nmat.col_n[23] 7.03fF
C14045 a_4719_30287# a_5535_29980# 0.40fF
C14046 a_47278_18528# vcm 0.65fF
C14047 VDD a_31214_20536# 0.52fF
C14048 a_18546_71232# a_28110_71190# 0.35fF
C14049 a_20170_67174# vcm 0.62fF
C14050 a_5403_67655# a_5081_53135# 1.20fF
C14051 _1183_.A2 vcm 0.46fF
C14052 VDD a_43262_17524# 0.52fF
C14053 a_12658_42895# a_16355_43123# 0.69fF
C14054 pmat.sample pmat.row_n[5] 0.46fF
C14055 a_22199_30287# a_7109_29423# 3.90fF
C14056 a_18546_8486# a_36142_8894# 0.35fF
C14057 VDD a_10291_77269# 0.38fF
C14058 a_21174_60146# a_21174_59142# 1.00fF
C14059 a_18546_65208# a_33130_65166# 0.35fF
C14060 a_10055_31591# a_16083_50069# 0.49fF
C14061 VDD a_44266_8488# 0.55fF
C14062 nmat.col[7] ctopn 1.97fF
C14063 nmat.col[17] ctopn 2.01fF
C14064 a_11416_50363# a_11455_50237# 0.53fF
C14065 a_18546_21538# a_47186_21946# 0.35fF
C14066 VDD pmat.col_n[13] 5.23fF
C14067 a_39246_62154# a_39246_61150# 1.00fF
C14068 pmat.rowoff_n[4] a_18546_60188# 4.09fF
C14069 a_12461_29673# a_16478_29423# 0.68fF
C14070 a_7521_47081# a_9135_60967# 0.71fF
C14071 nmat.col[30] nmat.col_n[29] 6.77fF
C14072 a_25190_67174# a_26194_67174# 0.97fF
C14073 a_18546_67216# a_33130_67174# 0.35fF
C14074 a_4081_61127# a_5053_59575# 0.37fF
C14075 ANTENNA__1196__A2.DIODE nmat.col_n[3] 2.97fF
C14076 _1194_.B1 _1183_.A2 3.78fF
C14077 pmat.row_n[15] pmat.rowon_n[12] 0.41fF
C14078 ANTENNA__1190__A1.DIODE nmat.col_n[31] 1.70fF
C14079 m2_17932_71010# m2_17932_70006# 0.99fF
C14080 a_22178_66170# a_22178_65166# 1.00fF
C14081 a_39246_15516# a_39246_14512# 1.00fF
C14082 VDD a_19166_65166# 0.56fF
C14083 a_14839_20871# a_13479_26935# 1.72fF
C14084 a_18546_7482# a_33130_7890# 0.35fF
C14085 a_13459_28111# a_15667_27239# 1.63fF
C14086 a_41254_69182# a_41254_68178# 1.00fF
C14087 VDD a_7847_56085# 0.50fF
C14088 a_49286_21540# a_49286_20536# 1.00fF
C14089 VDD a_1591_67503# 1.67fF
C14090 VDD a_39246_12504# 0.52fF
C14091 a_9441_20189# a_10498_19631# 0.61fF
C14092 a_6283_31591# a_4707_32156# 0.39fF
C14093 VDD a_5785_48463# 0.96fF
C14094 ANTENNA__1197__B.DIODE a_7717_14735# 1.14fF
C14095 pmat.rowon_n[10] a_18162_66210# 1.19fF
C14096 a_18546_66212# a_19074_66170# 0.35fF
C14097 _1224_.X ANTENNA__1184__B1.DIODE 0.51fF
C14098 VDD a_3688_65987# 0.65fF
C14099 a_47278_57134# vcm 0.62fF
C14100 a_46274_71190# vcm 0.60fF
C14101 a_25695_28111# nmat.col_n[29] 0.43fF
C14102 a_50290_18528# ctopn 3.43fF
C14103 a_33222_58138# vcm 0.62fF
C14104 a_39246_56130# m2_39016_54946# 0.99fF
C14105 nmat.col[19] comp_latch 0.84fF
C14106 cgen.dlycontrol1_in[0] a_2648_29397# 0.71fF
C14107 m2_51064_55950# m3_51196_56082# 2.76fF
C14108 _1192_.A2 a_18243_28327# 1.75fF
C14109 a_18546_19530# a_22086_19938# 0.35fF
C14110 VDD a_10883_3303# 15.95fF
C14111 a_18546_12502# a_26102_12910# 0.35fF
C14112 a_4719_30287# a_5785_48463# 0.64fF
C14113 a_2215_47375# a_2315_44124# 0.42fF
C14114 pmat.row_n[15] a_4257_34319# 1.33fF
C14115 VDD a_22178_16520# 0.52fF
C14116 a_2411_43301# a_8907_48437# 0.33fF
C14117 m2_17932_10226# m2_17932_9222# 0.99fF
C14118 pmat.col_n[5] m2_23956_54946# 0.37fF
C14119 VDD m2_42028_24282# 0.62fF
C14120 VDD a_27236_46831# 0.31fF
C14121 a_5179_31591# a_18597_31599# 8.88fF
C14122 nmat.col_n[6] ctopn 2.02fF
C14123 a_10515_13967# a_12447_16143# 1.53fF
C14124 pmat.rowoff_n[7] a_1586_18231# 1.80fF
C14125 VDD a_32126_7890# 0.33fF
C14126 a_24833_34191# a_11057_35836# 0.63fF
C14127 a_43262_11500# a_43262_10496# 1.00fF
C14128 a_18546_10494# a_18162_10496# 2.61fF
C14129 VDD a_23655_35279# 0.50fF
C14130 a_25190_69182# vcm 0.62fF
C14131 VDD a_7829_71317# 0.67fF
C14132 a_12585_39355# a_12513_39100# 2.69fF
C14133 a_24186_23548# a_25190_23548# 0.97fF
C14134 a_18546_23546# a_31122_23954# 0.35fF
C14135 a_34002_44527# a_11149_40188# 0.31fF
C14136 cgen.dlycontrol4_in[3] cgen.dlycontrol4_in[2] 1.06fF
C14137 m2_23956_24282# vcm 0.42fF
C14138 nmat.rowon_n[12] vcm 0.55fF
C14139 pmat.rowon_n[3] ctopn 0.60fF
C14140 VDD a_17139_49551# 0.35fF
C14141 a_26194_9492# a_27198_9492# 0.97fF
C14142 a_18546_9490# a_35138_9898# 0.35fF
C14143 a_48282_61150# a_49286_61150# 0.97fF
C14144 a_19166_70186# a_20170_70186# 0.97fF
C14145 a_34226_59142# vcm 0.62fF
C14146 VDD a_19166_61150# 0.56fF
C14147 a_1586_8439# a_6559_6031# 0.53fF
C14148 a_33222_12504# a_33222_11500# 1.00fF
C14149 VDD a_21815_42351# 0.37fF
C14150 ANTENNA__1196__A2.DIODE nmat.col[1] 1.31fF
C14151 _1154_.X _1183_.A2 1.82fF
C14152 pmat.rowon_n[7] a_4075_31591# 1.04fF
C14153 a_29206_56130# ctopp 3.40fF
C14154 a_2124_56891# a_2163_56765# 0.76fF
C14155 a_9668_10651# a_10378_7637# 1.06fF
C14156 a_3663_9269# a_5654_9527# 0.68fF
C14157 a_18162_70226# ctopp 1.49fF
C14158 VDD a_38242_56130# 0.55fF
C14159 a_42258_20536# a_43262_20536# 0.97fF
C14160 a_28202_8488# m2_27972_7214# 1.00fF
C14161 VDD a_1591_26159# 0.37fF
C14162 VDD m3_40152_72146# 0.33fF
C14163 a_21174_21540# ctopn 3.58fF
C14164 _1224_.X ANTENNA_fanout52_A.DIODE 12.75fF
C14165 ANTENNA__1395__A1.DIODE _1194_.B1 0.55fF
C14166 VDD a_1775_47375# 0.61fF
C14167 a_18546_66212# a_48190_66170# 0.35fF
C14168 a_41254_9492# a_41254_8488# 1.00fF
C14169 a_32218_66170# ctopp 3.58fF
C14170 VDD a_41254_66170# 0.52fF
C14171 a_23182_21540# a_24186_21540# 0.97fF
C14172 VDD a_10873_36341# 5.71fF
C14173 a_25190_63158# ctopp 3.58fF
C14174 a_6664_26159# a_9741_28585# 0.62fF
C14175 VDD a_34226_63158# 0.52fF
C14176 a_1769_13103# a_1586_33927# 1.91fF
C14177 m2_51064_58962# vcm 0.54fF
C14178 a_18546_61192# a_33130_61150# 0.35fF
C14179 m2_39016_54946# m2_40020_54946# 0.96fF
C14180 a_24186_71190# a_24186_70186# 1.00fF
C14181 VDD a_18162_68218# 2.73fF
C14182 nmat.sw inn_analog 0.91fF
C14183 pmat.sample pmat.row_n[13] 0.51fF
C14184 a_2411_16101# a_1591_20181# 0.33fF
C14185 a_38242_58138# a_39246_58138# 0.97fF
C14186 a_44774_40821# a_32405_32463# 0.62fF
C14187 nmat.rowoff_n[6] a_11235_26159# 0.36fF
C14188 VDD a_45861_29967# 1.10fF
C14189 a_34226_19532# vcm 0.65fF
C14190 a_18546_7482# a_19074_7890# 0.35fF
C14191 VDD cgen.dlycontrol1_in[3] 6.24fF
C14192 pmat.row_n[15] a_18546_71232# 0.35fF
C14193 a_33222_10496# vcm 0.65fF
C14194 a_10239_14183# a_5363_33551# 0.89fF
C14195 a_22178_13508# a_23182_13508# 0.97fF
C14196 a_18546_13506# a_27106_13914# 0.35fF
C14197 _1154_.X a_34204_27765# 0.90fF
C14198 VDD a_5687_71829# 5.19fF
C14199 pmat.row_n[10] pmat.rowon_n[3] 1.79fF
C14200 a_38242_61150# a_38242_60146# 1.00fF
C14201 a_30210_67174# ctopp 3.58fF
C14202 VDD a_22153_37179# 7.75fF
C14203 pmat.col_n[8] pmat.col[9] 6.42fF
C14204 a_46274_19532# a_46274_18528# 1.00fF
C14205 a_18546_18526# a_23090_18934# 0.35fF
C14206 a_18546_70228# a_50198_70186# 0.35fF
C14207 VDD a_39246_67174# 0.52fF
C14208 VDD a_37463_38007# 0.64fF
C14209 VDD a_2847_41151# 0.38fF
C14210 VDD a_28202_14512# 0.52fF
C14211 a_13091_28327# a_25695_28111# 3.67fF
C14212 a_49286_62154# vcm 0.62fF
C14213 VDD a_27198_64162# 0.52fF
C14214 a_18546_17522# a_45178_17930# 0.35fF
C14215 a_2046_30184# a_2051_29973# 0.56fF
C14216 a_18546_57176# a_41162_57134# 0.35fF
C14217 nmat.col[28] nmat.col[19] 2.80fF
C14218 a_13091_28327# a_1781_9308# 0.40fF
C14219 a_39246_59142# a_39246_58138# 1.00fF
C14220 VDD a_4583_68021# 2.65fF
C14221 a_47278_8488# m2_47048_7214# 1.00fF
C14222 m3_50768_55078# ctopp 0.38fF
C14223 a_38242_23548# m2_38012_24282# 0.99fF
C14224 VDD a_5597_44807# 0.44fF
C14225 a_12658_42895# a_10781_42364# 1.31fF
C14226 a_31214_15516# a_32218_15516# 0.97fF
C14227 a_18546_15514# a_45178_15922# 0.35fF
C14228 a_18162_64202# vcm 6.95fF
C14229 VDD m2_38012_54946# 0.62fF
C14230 nmat.sw a_14773_37218# 1.02fF
C14231 a_8305_20871# a_10957_14191# 0.59fF
C14232 nmat.rowoff_n[5] ctopn 0.60fF
C14233 a_30210_69182# a_31214_69182# 0.97fF
C14234 VDD a_41427_32143# 0.40fF
C14235 VDD a_27789_36039# 1.26fF
C14236 pmat.sample pmat.row_n[11] 0.42fF
C14237 a_11067_64015# a_12851_28853# 0.54fF
C14238 a_48282_70186# vcm 0.62fF
C14239 a_44774_48695# a_45370_48169# 0.31fF
C14240 pmat.row_n[6] pmat.row_n[1] 0.33fF
C14241 a_35230_11500# vcm 0.65fF
C14242 _1154_.X ANTENNA__1395__A1.DIODE 1.05fF
C14243 VDD a_13205_62607# 0.41fF
C14244 ANTENNA__1197__A.DIODE nmat.col[31] 1.10fF
C14245 ANTENNA__1395__A2.DIODE _1194_.B1 4.00fF
C14246 a_44266_17524# a_44266_16520# 1.00fF
C14247 a_18546_16518# a_20078_16926# 0.35fF
C14248 a_21174_8488# ctopn 3.40fF
C14249 a_18546_56172# a_24094_56130# 0.35fF
C14250 a_11435_58791# a_10515_13967# 0.72fF
C14251 VDD a_23090_24958# 0.44fF
C14252 pmat.row_n[14] a_18546_70228# 0.36fF
C14253 VDD a_17845_27791# 0.34fF
C14254 nmat.col[31] clk_comp 1.05fF
C14255 a_27603_34191# a_11681_35823# 0.31fF
C14256 pmat.col_n[15] vcm 2.79fF
C14257 a_1781_9308# a_27155_31599# 0.62fF
C14258 a_37238_19532# ctopn 3.58fF
C14259 a_21174_65166# ctopp 3.58fF
C14260 a_19166_14512# a_20170_14512# 0.97fF
C14261 VDD a_30210_65166# 0.52fF
C14262 a_7717_14735# a_22459_28879# 0.53fF
C14263 VDD a_10589_22351# 2.85fF
C14264 ANTENNA__1190__B1.DIODE a_47039_31599# 0.50fF
C14265 VDD a_37238_21540# 0.52fF
C14266 a_39246_59142# a_40250_59142# 0.97fF
C14267 _1192_.A2 a_30571_50959# 0.31fF
C14268 a_36234_10496# ctopn 3.58fF
C14269 a_18546_68220# a_32126_68178# 0.35fF
C14270 a_43262_58138# ctopp 3.58fF
C14271 a_39246_68178# vcm 0.62fF
C14272 cgen.dlycontrol3_in[2] a_14379_6567# 0.43fF
C14273 a_2411_43301# a_6553_53047# 0.42fF
C14274 VDD a_7140_27805# 1.25fF
C14275 a_28202_23548# a_28202_22544# 1.00fF
C14276 VDD a_5731_17455# 0.32fF
C14277 a_22199_30287# inn_analog 2.35fF
C14278 a_27198_60146# a_28202_60146# 0.97fF
C14279 a_18546_60188# a_37146_60146# 0.35fF
C14280 a_5462_62215# a_12889_64789# 0.30fF
C14281 a_8031_64789# a_8197_64789# 0.42fF
C14282 nmat.rowon_n[14] a_1586_18231# 2.50fF
C14283 a_14691_29575# a_8443_20719# 0.60fF
C14284 a_11067_64015# a_2046_30184# 1.26fF
C14285 a_1923_61759# a_2124_65595# 0.40fF
C14286 a_17139_30503# a_25695_28111# 0.96fF
C14287 nmat.rowoff_n[0] ctopn 0.51fF
C14288 VDD m2_23956_72014# 1.15fF
C14289 a_35230_68178# a_35230_67174# 1.00fF
C14290 a_44266_23548# vcm 0.65fF
C14291 a_35230_69182# ctopp 3.58fF
C14292 a_2389_45859# a_4399_51157# 0.58fF
C14293 VDD a_44266_69182# 0.52fF
C14294 a_46274_9492# vcm 0.65fF
C14295 a_18546_60188# vcm 0.40fF
C14296 m2_24960_72014# m2_25964_72014# 0.96fF
C14297 VDD a_13503_39069# 1.25fF
C14298 VDD a_22449_44219# 1.32fF
C14299 a_43262_62154# pmat.col[24] 0.31fF
C14300 a_44266_59142# ctopp 3.58fF
C14301 a_38242_11500# ctopn 3.58fF
C14302 pmat.row_n[10] nmat.rowoff_n[5] 0.32fF
C14303 VDD a_15144_35077# 1.10fF
C14304 _1194_.B1 ANTENNA__1196__A2.DIODE 3.13fF
C14305 ANTENNA__1197__B.DIODE ANTENNA__1195__A1.DIODE 0.46fF
C14306 a_11067_27239# a_13459_28111# 1.15fF
C14307 a_8491_47911# a_11007_58229# 0.34fF
C14308 a_5351_19913# a_13768_22325# 0.30fF
C14309 VDD a_18162_71230# 2.78fF
C14310 a_22199_30287# nmat.col[26] 0.54fF
C14311 pmat.rowon_n[2] a_18162_58178# 1.19fF
C14312 a_18546_58180# a_19074_58138# 0.35fF
C14313 a_18546_16518# a_49194_16926# 0.35fF
C14314 a_33222_16520# a_34226_16520# 0.97fF
C14315 m2_47048_24282# vcm 0.42fF
C14316 VDD a_41335_49551# 0.47fF
C14317 a_23182_67174# a_23182_66170# 1.00fF
C14318 a_9581_56079# a_6559_33767# 0.35fF
C14319 a_21174_61150# ctopp 3.58fF
C14320 a_13459_28111# a_35312_31599# 0.39fF
C14321 a_2419_53351# a_2263_43719# 1.15fF
C14322 VDD a_30210_61150# 0.52fF
C14323 _1154_.X ANTENNA__1395__A2.DIODE 0.51fF
C14324 a_42258_13508# vcm 0.65fF
C14325 a_18546_15514# nmat.rowoff_n[8] 4.09fF
C14326 a_14917_23983# a_13479_26935# 0.38fF
C14327 a_40250_18528# vcm 0.65fF
C14328 VDD a_24186_20536# 0.52fF
C14329 a_5363_33551# a_10147_29415# 0.93fF
C14330 a_22178_17524# a_23182_17524# 0.97fF
C14331 nmat.sw clk_ena 1.95fF
C14332 VDD a_83217_4649# 0.35fF
C14333 a_20170_57134# a_21174_57134# 0.97fF
C14334 ANTENNA__1195__A1.DIODE a_31675_47695# 0.73fF
C14335 VDD a_17323_27791# 0.33fF
C14336 a_25190_20536# a_25190_19532# 1.00fF
C14337 a_18546_71232# a_21082_71190# 0.35fF
C14338 VDD clk_vcm 2.78fF
C14339 VDD a_36234_17524# 0.52fF
C14340 VDD m2_18936_55950# 0.57fF
C14341 VDD a_22276_46831# 0.59fF
C14342 _1183_.A2 a_40837_46261# 0.32fF
C14343 a_23182_8488# a_24186_8488# 0.97fF
C14344 a_18546_8486# a_29114_8894# 0.35fF
C14345 a_13432_62581# a_1957_43567# 0.53fF
C14346 a_18546_65208# a_26102_65166# 0.35fF
C14347 cgen.dlycontrol3_in[0] a_13909_39605# 2.27fF
C14348 pmat.row_n[11] a_1923_31743# 0.39fF
C14349 a_42258_70186# a_42258_69182# 1.00fF
C14350 VDD a_7717_14735# 17.36fF
C14351 VDD a_37238_8488# 0.55fF
C14352 pmat.row_n[15] ctopp 1.37fF
C14353 a_43776_30287# a_40951_31599# 0.68fF
C14354 a_18546_21538# a_40158_21946# 0.35fF
C14355 VDD a_27619_36649# 0.62fF
C14356 VDD a_82863_64213# 0.98fF
C14357 a_31214_14512# a_31214_13508# 1.00fF
C14358 a_10147_29415# a_28336_29967# 0.67fF
C14359 a_47278_23548# ctopn 3.40fF
C14360 VDD a_5087_18543# 0.45fF
C14361 a_49286_9492# ctopn 3.56fF
C14362 m2_38012_24282# m3_38144_24414# 2.79fF
C14363 nmat.col[3] ctopn 1.97fF
C14364 a_18546_67216# a_26102_67174# 0.35fF
C14365 a_35230_57134# a_35230_56130# 1.00fF
C14366 a_39246_19532# a_40250_19532# 0.97fF
C14367 m2_50060_54946# m2_51064_54946# 0.59fF
C14368 a_47278_60146# vcm 0.62fF
C14369 a_1591_31599# cgen.dlycontrol4_in[0] 1.51fF
C14370 a_14917_23983# a_5351_19913# 1.06fF
C14371 pmat.rowon_n[10] pmat.rowon_n[9] 0.78fF
C14372 a_19166_19532# ctopn 3.43fF
C14373 a_26891_28327# a_25695_28111# 1.32fF
C14374 VDD a_30103_43447# 0.62fF
C14375 VDD a_5589_14967# 0.39fF
C14376 a_2149_45717# a_3936_70197# 0.68fF
C14377 pmat.col[0] ctopp 1.55fF
C14378 a_2163_31741# a_2422_29575# 0.39fF
C14379 a_9963_28111# a_14691_27399# 0.31fF
C14380 a_18546_7482# a_26102_7890# 0.35fF
C14381 VDD a_19166_21540# 0.58fF
C14382 a_9963_13967# pmat.row_n[2] 0.40fF
C14383 a_6007_33767# a_5179_31591# 0.87fF
C14384 a_38242_10496# a_39246_10496# 0.97fF
C14385 VDD a_32218_12504# 0.52fF
C14386 nmat.col_n[12] ctopn 2.02fF
C14387 VDD a_30189_48437# 0.60fF
C14388 a_49286_56130# a_50290_56130# 0.97fF
C14389 a_18546_60188# a_18162_60186# 2.62fF
C14390 _1154_.X ANTENNA__1196__A2.DIODE 4.31fF
C14391 a_45270_13508# ctopn 3.58fF
C14392 a_14653_53458# a_13091_52047# 0.40fF
C14393 VDD pmat.row_n[3] 18.14fF
C14394 a_40250_57134# vcm 0.62fF
C14395 VDD a_14712_37429# 2.24fF
C14396 a_39246_71190# vcm 0.60fF
C14397 pmat.rowoff_n[7] a_1923_53055# 0.83fF
C14398 a_43262_18528# ctopn 3.58fF
C14399 a_26194_58138# vcm 0.62fF
C14400 ANTENNA__1183__B1.DIODE nmat.col[19] 3.71fF
C14401 m2_29980_7214# m3_30112_7346# 2.79fF
C14402 pmat.en_bit_n[2] a_15101_29423# 0.92fF
C14403 nmat.col_n[12] a_10147_29415# 2.37fF
C14404 VDD a_7521_19631# 0.63fF
C14405 nmat.col[7] m2_25964_24282# 0.40fF
C14406 VDD a_33007_38771# 1.12fF
C14407 m2_17932_61974# vcm 0.44fF
C14408 _1184_.A2 a_1781_9308# 0.40fF
C14409 a_10883_3303# a_4523_21276# 0.56fF
C14410 pmat.sample pmat.row_n[2] 0.92fF
C14411 a_82818_69135# _1154_.X 1.16fF
C14412 pmat.row_n[8] nmat.en_bit_n[1] 5.89fF
C14413 VDD a_9668_10651# 1.55fF
C14414 cgen.start_conv_in a_12309_38659# 0.97fF
C14415 a_9963_13967# nmat.col_n[13] 1.53fF
C14416 VDD m3_27100_7346# 0.36fF
C14417 a_31214_22544# a_32218_22544# 0.97fF
C14418 VDD config_1_in[3] 0.97fF
C14419 a_18546_20534# ctopn 1.59fF
C14420 VDD a_25090_46831# 0.46fF
C14421 a_9963_13967# nmat.rowoff_n[6] 1.23fF
C14422 a_5363_33551# a_4707_32156# 0.42fF
C14423 pmat.row_n[7] pmat.row_n[6] 0.36fF
C14424 a_20170_11500# ctopn 3.57fF
C14425 VDD a_21279_31599# 0.46fF
C14426 VDD a_25098_7890# 0.33fF
C14427 pmat.col_n[23] ctopp 2.02fF
C14428 a_10883_3303# a_22499_49783# 1.05fF
C14429 VDD a_7079_34837# 0.56fF
C14430 a_12987_26159# a_13145_26935# 0.36fF
C14431 a_5351_19913# a_9441_20189# 1.13fF
C14432 VDD a_49194_72194# 0.32fF
C14433 a_1923_61759# pmat.rowoff_n[7] 1.06fF
C14434 a_18546_23546# a_24094_23954# 0.35fF
C14435 a_10147_29415# a_35559_30209# 0.62fF
C14436 a_4259_31375# a_4075_31591# 0.31fF
C14437 a_45270_63158# a_46274_63158# 0.97fF
C14438 m2_43032_54946# vcm 0.42fF
C14439 a_1586_18231# a_1757_26159# 0.42fF
C14440 a_18546_9490# a_28110_9898# 0.35fF
C14441 a_49286_68178# ctopp 3.57fF
C14442 a_6830_22895# a_5351_19913# 0.74fF
C14443 a_41926_46983# a_42024_46805# 0.56fF
C14444 a_27198_59142# vcm 0.62fF
C14445 a_18180_38341# a_13597_37571# 0.31fF
C14446 ANTENNA__1195__A1.DIODE a_28812_29575# 0.74fF
C14447 a_2021_9563# a_2021_11043# 0.69fF
C14448 a_12228_40693# a_11297_36091# 0.43fF
C14449 VDD cgen.dlycontrol2_in[3] 7.37fF
C14450 ANTENNA__1395__A1.DIODE a_40837_46261# 0.51fF
C14451 pmat.row_n[11] nmat.rowon_n[4] 20.98fF
C14452 a_13909_39605# a_12969_40175# 0.96fF
C14453 a_24374_29941# a_7415_29397# 0.43fF
C14454 a_25695_28111# a_9411_2215# 2.36fF
C14455 a_22178_56130# ctopp 3.40fF
C14456 a_13319_35507# cgen.dlycontrol1_in[3] 0.35fF
C14457 VDD a_31214_56130# 0.55fF
C14458 a_7644_16341# a_4383_7093# 0.38fF
C14459 a_18546_72236# a_26102_72194# 0.35fF
C14460 VDD a_8031_26703# 0.32fF
C14461 VDD m2_50060_7214# 0.96fF
C14462 ANTENNA__1190__B1.DIODE a_41731_49525# 1.50fF
C14463 ANTENNA__1190__A1.DIODE a_37820_30485# 0.57fF
C14464 _1224_.X a_13091_28327# 1.72fF
C14465 a_2199_13887# config_1_in[0] 0.36fF
C14466 a_18546_62196# a_45178_62154# 0.35fF
C14467 _1196_.B1 a_13459_28111# 0.85fF
C14468 VDD a_25384_48169# 0.44fF
C14469 a_18546_66212# a_41162_66170# 0.35fF
C14470 a_25190_66170# ctopp 3.58fF
C14471 m2_21948_72014# m3_22080_72146# 2.79fF
C14472 a_2215_47375# a_1739_47893# 0.46fF
C14473 VDD a_34226_66170# 0.52fF
C14474 ANTENNA__1190__A1.DIODE _1183_.A2 2.32fF
C14475 a_40250_11500# a_41254_11500# 0.97fF
C14476 VDD a_8283_71829# 0.39fF
C14477 nmat.col_n[17] vcm 2.79fF
C14478 VDD a_27198_63158# 0.52fF
C14479 a_20170_24552# a_20170_23548# 1.00fF
C14480 a_42258_64162# a_42258_63158# 1.00fF
C14481 m2_47048_54946# m3_47180_55078# 2.79fF
C14482 a_29937_31055# a_44573_45173# 1.05fF
C14483 a_45270_10496# a_45270_9492# 1.00fF
C14484 a_18546_61192# a_26102_61150# 0.35fF
C14485 VDD a_11837_68591# 0.51fF
C14486 a_42258_58138# a_42258_57134# 1.00fF
C14487 a_1586_63927# a_8197_64789# 0.60fF
C14488 VDD a_37463_39095# 0.64fF
C14489 a_1781_9308# a_7939_31591# 2.66fF
C14490 ANTENNA__1184__B1.DIODE ANTENNA__1183__B1.DIODE 1.46fF
C14491 a_18162_63198# vcm 6.95fF
C14492 a_27198_19532# vcm 0.65fF
C14493 a_46274_60146# a_46274_59142# 1.00fF
C14494 a_34226_18528# a_34226_17524# 1.00fF
C14495 a_37238_63158# pmat.col[18] 0.31fF
C14496 VDD a_15259_31029# 0.50fF
C14497 VDD a_3247_6037# 0.52fF
C14498 VDD pmat.row_n[1] 18.29fF
C14499 a_26194_10496# vcm 0.65fF
C14500 nmat.col_n[18] ctopn 2.03fF
C14501 VDD a_10839_11989# 1.10fF
C14502 a_18546_13506# a_19074_13914# 0.35fF
C14503 a_11927_27399# a_12987_26159# 0.65fF
C14504 a_34226_63158# a_34226_62154# 1.00fF
C14505 VDD m2_51064_63982# 1.18fF
C14506 a_2935_38279# a_2411_33749# 0.35fF
C14507 a_14641_57711# a_9963_13967# 0.32fF
C14508 pmat.rowoff_n[12] a_12447_16143# 2.96fF
C14509 a_1769_13103# start_conversion_in 0.42fF
C14510 a_1899_35051# a_10055_31591# 0.67fF
C14511 VDD a_11159_23145# 0.48fF
C14512 a_23182_67174# ctopp 3.58fF
C14513 VDD a_17499_38825# 0.63fF
C14514 a_18546_70228# a_43170_70186# 0.35fF
C14515 VDD a_32218_67174# 0.52fF
C14516 VDD a_18546_9490# 32.63fF
C14517 VDD a_20811_38007# 0.60fF
C14518 a_47278_66170# a_47278_65166# 1.00fF
C14519 a_40250_22544# a_40250_21540# 1.00fF
C14520 nmat.col_n[21] m2_40020_24282# 0.37fF
C14521 VDD a_33489_42043# 1.14fF
C14522 VDD a_21174_14512# 0.52fF
C14523 a_22178_56130# m2_21948_54946# 0.99fF
C14524 a_39246_14512# a_40250_14512# 0.97fF
C14525 a_42258_62154# vcm 0.62fF
C14526 VDD a_20170_64162# 0.52fF
C14527 ANTENNA__1190__A2.DIODE a_3571_13627# 0.42fF
C14528 m2_50060_54946# clk_ena 0.58fF
C14529 a_19283_49783# a_21279_48999# 2.08fF
C14530 a_11711_58261# a_1957_43567# 0.31fF
C14531 a_18546_17522# a_38150_17930# 0.35fF
C14532 a_38242_64162# a_39246_64162# 0.97fF
C14533 a_44266_68178# a_45270_68178# 0.97fF
C14534 a_18546_57176# a_34134_57134# 0.35fF
C14535 pmat.col[14] m2_32992_54946# 0.39fF
C14536 VDD a_1643_54965# 0.38fF
C14537 a_33222_13508# a_33222_12504# 1.00fF
C14538 ANTENNA__1395__A2.DIODE a_40837_46261# 0.53fF
C14539 a_1899_35051# a_1591_31599# 0.49fF
C14540 pmat.rowon_n[8] a_4955_40277# 0.60fF
C14541 VDD a_9339_28335# 0.37fF
C14542 a_18546_15514# a_38150_15922# 0.35fF
C14543 VDD a_38391_47381# 0.43fF
C14544 a_4259_73807# a_4025_54965# 0.39fF
C14545 pmat.rowon_n[3] ctopp 1.57fF
C14546 VDD a_2099_49525# 0.50fF
C14547 a_1591_67503# a_2124_67771# 0.61fF
C14548 VDD a_9963_28111# 4.09fF
C14549 a_41254_70186# vcm 0.62fF
C14550 VDD pmat.col_n[16] 5.31fF
C14551 a_28202_11500# vcm 0.65fF
C14552 VDD a_5173_9839# 1.25fF
C14553 a_24747_29967# a_15667_28111# 1.80fF
C14554 VDD pmat.col[19] 4.88fF
C14555 _1194_.A2 _1192_.A2 11.76fF
C14556 pmat.row_n[0] a_18546_56172# 0.35fF
C14557 _1154_.A a_30663_50087# 2.96fF
C14558 a_19166_64162# m2_17932_63982# 0.96fF
C14559 a_19166_19532# a_19166_18528# 1.00fF
C14560 ANTENNA_fanout52_A.DIODE ANTENNA__1183__B1.DIODE 2.83fF
C14561 a_13091_28327# comp_latch 0.33fF
C14562 a_30210_19532# ctopn 3.58fF
C14563 a_1586_50247# a_5639_49007# 0.33fF
C14564 VDD a_23182_65166# 0.52fF
C14565 VDD a_3944_28853# 0.32fF
C14566 a_2407_49289# a_6451_67655# 0.77fF
C14567 VDD a_30210_21540# 0.52fF
C14568 ANTENNA__1197__A.DIODE a_24867_53135# 1.53fF
C14569 ANTENNA__1395__A1.DIODE ANTENNA__1190__A1.DIODE 2.74fF
C14570 a_40250_65166# a_40250_64162# 1.00fF
C14571 a_29206_10496# ctopn 3.58fF
C14572 a_18546_68220# a_25098_68178# 0.35fF
C14573 a_50290_57134# ctopp 3.42fF
C14574 VDD a_31323_29967# 0.33fF
C14575 a_49286_71190# ctopp 3.39fF
C14576 a_36234_58138# ctopp 3.58fF
C14577 a_32218_68178# vcm 0.62fF
C14578 a_11067_30287# a_32687_46607# 0.43fF
C14579 VDD a_45270_58138# 0.52fF
C14580 VDD nmat.col[21] 7.22fF
C14581 a_49286_23548# a_50290_23548# 0.97fF
C14582 a_10515_13967# a_19541_28879# 0.38fF
C14583 VDD ANTENNA__1195__A1.DIODE 17.39fF
C14584 cgen.dlycontrol4_in[2] a_30543_40721# 1.84fF
C14585 a_22178_62154# a_23182_62154# 0.97fF
C14586 a_29206_16520# a_29206_15516# 1.00fF
C14587 VDD a_40897_48463# 0.40fF
C14588 a_20170_66170# a_21174_66170# 0.97fF
C14589 a_18546_60188# a_30118_60146# 0.35fF
C14590 VDD pmat.rowon_n[8] 16.00fF
C14591 a_19166_21540# m2_17932_21270# 0.96fF
C14592 cgen.dlycontrol2_in[0] a_11041_36596# 3.22fF
C14593 VDD a_38651_37737# 0.60fF
C14594 a_10239_14183# pmat.row_n[4] 0.80fF
C14595 a_8583_29199# a_10589_22351# 1.32fF
C14596 a_13641_23439# a_31263_28309# 1.76fF
C14597 pmat.col[25] vcm 5.88fF
C14598 a_1923_31743# a_4167_30511# 0.35fF
C14599 pmat.rowon_n[3] a_1586_50247# 1.46fF
C14600 a_37238_23548# vcm 0.65fF
C14601 a_28202_69182# ctopp 3.58fF
C14602 a_39246_9492# vcm 0.65fF
C14603 VDD a_37238_69182# 0.52fF
C14604 VDD a_9583_10121# 1.22fF
C14605 VDD a_16879_50345# 0.39fF
C14606 a_1586_18231# a_1591_23445# 0.54fF
C14607 m2_17932_72014# m2_18936_72014# 0.96fF
C14608 a_1674_68047# a_3339_59879# 0.33fF
C14609 VDD a_29367_44535# 0.59fF
C14610 pmat.rowon_n[8] a_4719_30287# 0.42fF
C14611 a_9963_13967# a_6927_30503# 6.00fF
C14612 a_41254_65166# a_42258_65166# 0.97fF
C14613 pmat.rowoff_n[2] ctopp 0.60fF
C14614 a_37238_59142# ctopp 3.58fF
C14615 a_31214_11500# ctopn 3.58fF
C14616 VDD a_46274_59142# 0.52fF
C14617 a_48282_21540# a_49286_21540# 0.97fF
C14618 VDD a_45829_35407# 0.71fF
C14619 a_4583_68021# a_4128_64391# 0.64fF
C14620 a_10781_42869# a_11317_40188# 1.52fF
C14621 a_18546_16518# a_42166_16926# 0.35fF
C14622 _1519_.A vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot 0.81fF
C14623 VDD a_25839_49783# 1.75fF
C14624 nmat.col[30] nmat.col[24] 1.78fF
C14625 a_49286_71190# a_49286_70186# 1.00fF
C14626 a_21174_70186# a_22178_70186# 0.97fF
C14627 VDD a_23182_61150# 0.52fF
C14628 a_14773_38306# a_22059_37683# 0.48fF
C14629 a_35230_13508# vcm 0.65fF
C14630 nmat.en_bit_n[1] _1192_.B1 0.77fF
C14631 a_33222_18528# vcm 0.65fF
C14632 VDD a_32865_30199# 0.41fF
C14633 a_4259_73807# a_2407_49289# 2.08fF
C14634 pmat.rowoff_n[12] a_11435_58791# 0.60fF
C14635 a_4075_68583# a_4081_61127# 1.19fF
C14636 a_6200_70919# a_6795_76989# 0.45fF
C14637 nmat.rowoff_n[10] ctopn 0.60fF
C14638 a_21174_23548# m2_20944_24282# 0.99fF
C14639 a_47278_13508# a_48282_13508# 0.97fF
C14640 a_44266_15516# vcm 0.65fF
C14641 _1224_.X _1184_.A2 5.90fF
C14642 VDD a_29206_17524# 0.52fF
C14643 a_13503_43421# a_10781_42364# 0.44fF
C14644 _1194_.B1 a_31339_31787# 1.16fF
C14645 ANTENNA__1190__A1.DIODE ANTENNA__1395__A2.DIODE 0.32fF
C14646 ANTENNA__1190__B1.DIODE _1194_.B1 15.79fF
C14647 a_5087_32687# a_5253_32687# 0.39fF
C14648 a_18546_8486# a_22086_8894# 0.35fF
C14649 a_45270_18528# a_46274_18528# 0.97fF
C14650 a_3305_27791# a_4703_24527# 0.99fF
C14651 VDD a_30210_8488# 0.55fF
C14652 cgen.dlycontrol2_in[0] cgen.dlycontrol1_in[1] 1.54fF
C14653 a_18546_21538# a_33130_21946# 0.35fF
C14654 m2_51064_65990# m2_51064_64986# 0.99fF
C14655 a_32218_62154# a_32218_61150# 1.00fF
C14656 a_6175_60039# a_5682_56311# 0.99fF
C14657 pmat.sw m2_50060_54946# 0.33fF
C14658 a_40250_23548# ctopn 3.40fF
C14659 VDD a_46274_19532# 0.52fF
C14660 a_42258_9492# ctopn 3.57fF
C14661 a_11784_47099# a_11823_46973# 0.46fF
C14662 a_40250_60146# vcm 0.62fF
C14663 VDD a_45270_10496# 0.52fF
C14664 a_32218_15516# a_32218_14512# 1.00fF
C14665 VDD pmat.row_n[7] 17.75fF
C14666 a_7717_14735# a_8583_29199# 0.81fF
C14667 VDD a_16966_29673# 1.03fF
C14668 a_10055_31591# a_10515_15055# 1.34fF
C14669 a_18243_28327# a_16311_28327# 5.08fF
C14670 cgen.dlycontrol4_in[5] clk_dig 1.60fF
C14671 a_34226_69182# a_34226_68178# 1.00fF
C14672 VDD a_7415_29397# 10.32fF
C14673 a_11041_36596# cgen.dlycontrol1_in[2] 2.33fF
C14674 _1154_.X a_19405_28853# 0.39fF
C14675 a_42258_21540# a_42258_20536# 1.00fF
C14676 a_38391_48469# a_33423_47695# 0.62fF
C14677 VDD a_25190_12504# 0.52fF
C14678 a_20170_24552# m2_18936_24282# 0.96fF
C14679 a_46274_16520# vcm 0.65fF
C14680 a_11149_40188# a_12228_40693# 1.52fF
C14681 nmat.col_n[25] ctopn 2.02fF
C14682 a_35230_55126# vcm 0.58fF
C14683 a_38242_13508# ctopn 3.58fF
C14684 a_13459_28111# a_45019_38645# 0.33fF
C14685 a_12513_36924# a_11149_36924# 1.07fF
C14686 a_21219_36885# a_24015_36911# 0.31fF
C14687 a_11927_27399# comp_latch 1.89fF
C14688 a_33222_57134# vcm 0.62fF
C14689 VDD a_13597_37571# 0.73fF
C14690 a_32218_71190# vcm 0.60fF
C14691 a_36234_18528# ctopn 3.58fF
C14692 VDD a_15107_41271# 0.62fF
C14693 VDD a_16837_40955# 1.14fF
C14694 pmat.row_n[4] ctopn 1.65fF
C14695 pmat.col[28] m2_47048_54946# 0.39fF
C14696 a_4976_16091# a_4383_7093# 0.72fF
C14697 a_47278_15516# ctopn 3.58fF
C14698 VDD a_19166_69182# 0.58fF
C14699 ANTENNA_fanout52_A.DIODE a_38913_31055# 0.56fF
C14700 VDD a_47278_11500# 0.52fF
C14701 VDD pmat.col[21] 4.68fF
C14702 _1179_.X _1187_.A2 0.60fF
C14703 ANTENNA__1190__A1.DIODE ANTENNA__1196__A2.DIODE 1.03fF
C14704 a_13091_52047# a_16800_47213# 1.49fF
C14705 ANTENNA__1184__B1.DIODE a_21739_29415# 0.85fF
C14706 pmat.en_bit_n[0] a_11067_27239# 0.99fF
C14707 a_18546_58180# pmat.row_n[2] 0.36fF
C14708 a_14839_66103# pmat.rowoff_n[3] 2.73fF
C14709 a_19166_59142# ctopp 3.43fF
C14710 a_18546_69224# a_47186_69182# 0.35fF
C14711 a_36234_11500# a_36234_10496# 1.00fF
C14712 VDD vcm.sky130_fd_sc_hd__buf_4_3.A 1.00fF
C14713 _1154_.X ANTENNA__1190__B1.DIODE 1.97fF
C14714 a_2791_57703# a_3345_62839# 0.89fF
C14715 a_18546_22542# ctopn 1.58fF
C14716 VDD m2_17932_66994# 1.00fF
C14717 a_40837_46261# a_44966_43255# 1.52fF
C14718 a_44266_22544# vcm 0.65fF
C14719 a_41254_61150# a_42258_61150# 0.97fF
C14720 a_42258_68178# ctopp 3.58fF
C14721 a_20170_59142# vcm 0.62fF
C14722 _1184_.A2 comp_latch 0.74fF
C14723 a_26194_12504# a_26194_11500# 1.00fF
C14724 a_9441_20189# a_4383_7093# 0.38fF
C14725 pmat.col_n[18] vcm 2.80fF
C14726 a_14533_39631# a_12969_40175# 1.14fF
C14727 a_2315_44124# a_1739_47893# 1.29fF
C14728 VDD a_45212_30761# 0.37fF
C14729 cgen.dlycontrol1_in[1] cgen.dlycontrol1_in[2] 4.63fF
C14730 a_2046_30184# a_6007_33767# 0.42fF
C14731 a_41731_49525# inn_analog 0.38fF
C14732 VDD a_24186_56130# 0.55fF
C14733 a_4257_34319# a_2563_34837# 1.16fF
C14734 a_35230_20536# a_36234_20536# 0.97fF
C14735 a_2419_53351# a_3838_70455# 0.72fF
C14736 a_49286_16520# ctopn 3.57fF
C14737 VDD a_12152_66415# 1.09fF
C14738 VDD m2_36004_7214# 1.05fF
C14739 VDD a_1644_74549# 0.32fF
C14740 a_18546_62196# a_38150_62154# 0.35fF
C14741 VDD a_30687_48071# 0.60fF
C14742 a_18546_66212# a_34134_66170# 0.35fF
C14743 a_48282_67174# a_48282_66170# 1.00fF
C14744 a_34226_9492# a_34226_8488# 1.00fF
C14745 m2_17932_20266# m2_17932_19262# 0.99fF
C14746 a_5363_70543# a_5651_66975# 0.94fF
C14747 VDD a_27198_66170# 0.52fF
C14748 VDD a_12981_8213# 0.48fF
C14749 nmat.col_n[8] vcm 2.80fF
C14750 a_3746_58487# a_4705_39759# 0.32fF
C14751 VDD a_20170_63158# 0.52fF
C14752 a_4985_51433# a_4128_46983# 0.48fF
C14753 pmat.sample pmat.row_n[8] 0.58fF
C14754 a_47278_17524# a_48282_17524# 0.97fF
C14755 a_45270_57134# a_46274_57134# 0.97fF
C14756 a_18563_27791# clk_ena 0.46fF
C14757 a_38851_28327# a_45119_32661# 0.77fF
C14758 a_13091_28327# a_22307_27791# 0.96fF
C14759 a_50290_20536# a_50290_19532# 1.00fF
C14760 a_18162_66210# vcm 6.95fF
C14761 a_44266_71190# a_45270_71190# 0.97fF
C14762 a_10814_29111# a_7693_22365# 0.59fF
C14763 VDD a_22085_38550# 1.49fF
C14764 a_31214_58138# a_32218_58138# 0.97fF
C14765 a_9411_2215# comp_latch 0.32fF
C14766 VDD a_12197_43746# 1.41fF
C14767 pmat.rowoff_n[15] pmat.sample 0.38fF
C14768 a_48282_8488# a_49286_8488# 0.97fF
C14769 nmat.col[4] nmat.col_n[4] 0.75fF
C14770 a_30571_50959# a_38557_47381# 0.62fF
C14771 VDD a_9307_31068# 2.81fF
C14772 a_18162_10496# vcm 6.95fF
C14773 a_13091_7655# a_9528_20407# 0.95fF
C14774 a_47278_22544# ctopn 3.57fF
C14775 a_11317_40188# cgen.dlycontrol4_in[0] 0.30fF
C14776 pmat.col[11] ctopp 1.97fF
C14777 a_24186_71190# m2_23956_72014# 1.00fF
C14778 VDD a_8907_48437# 0.64fF
C14779 a_12693_38543# a_12585_37179# 0.71fF
C14780 a_31214_61150# a_31214_60146# 1.00fF
C14781 a_50290_64162# m2_51064_63982# 0.96fF
C14782 a_39246_19532# a_39246_18528# 1.00fF
C14783 a_20170_13508# ctopn 3.57fF
C14784 a_18546_70228# a_36142_70186# 0.35fF
C14785 VDD a_25190_67174# 0.52fF
C14786 VDD a_6956_8965# 0.31fF
C14787 VDD a_47357_38127# 0.60fF
C14788 a_8861_24527# a_8013_25615# 0.72fF
C14789 a_35230_62154# vcm 0.62fF
C14790 m2_51064_13238# vcm 0.51fF
C14791 VDD config_2_in[1] 0.96fF
C14792 _1154_.A a_10883_3303# 0.50fF
C14793 a_18546_17522# a_31122_17930# 0.35fF
C14794 a_18546_57176# a_27106_57134# 0.35fF
C14795 a_14641_57167# pmat.rowoff_n[6] 0.43fF
C14796 VDD nmat.col[9] 4.50fF
C14797 a_32218_59142# a_32218_58138# 1.00fF
C14798 a_13459_28111# nmat.sw 2.03fF
C14799 a_5351_19913# nmat.col[3] 0.48fF
C14800 a_18162_22544# nmat.rowon_n[1] 1.33fF
C14801 a_18546_22542# a_20078_22950# 0.35fF
C14802 VDD nmat.col_n[28] 10.90fF
C14803 a_24186_15516# a_25190_15516# 0.97fF
C14804 a_18546_15514# a_31122_15922# 0.35fF
C14805 a_16311_28327# a_30571_50959# 0.39fF
C14806 a_19166_20536# vcm 0.65fF
C14807 a_50290_60146# ctopp 3.43fF
C14808 a_23182_69182# a_24186_69182# 0.97fF
C14809 a_50290_21540# m2_51064_21270# 0.96fF
C14810 nmat.col_n[10] nmat.col_n[3] 1.29fF
C14811 VDD a_37129_36130# 1.09fF
C14812 a_4075_50087# a_5535_57993# 0.72fF
C14813 a_34226_70186# vcm 0.62fF
C14814 a_2791_57703# a_3615_71631# 0.42fF
C14815 a_21174_11500# vcm 0.65fF
C14816 a_10441_21263# a_14691_29575# 0.80fF
C14817 a_37238_17524# a_37238_16520# 1.00fF
C14818 m2_43032_24282# m3_43164_24414# 2.79fF
C14819 nmat.rowon_n[15] ctopn 1.19fF
C14820 pmat.row_n[14] pmat.rowoff_n[14] 0.49fF
C14821 a_43262_12504# a_44266_12504# 0.97fF
C14822 pmat.rowoff_n[8] a_18546_64204# 4.09fF
C14823 a_23182_19532# ctopn 3.58fF
C14824 a_11711_50959# a_10883_3303# 1.17fF
C14825 pmat.col_n[30] m2_49056_54946# 0.45fF
C14826 a_16311_28327# ANTENNA__1190__A2.DIODE 1.54fF
C14827 VDD a_36459_29673# 0.91fF
C14828 VDD a_23182_21540# 0.52fF
C14829 _1196_.B1 a_46582_46519# 1.09fF
C14830 a_32218_59142# a_33222_59142# 0.97fF
C14831 a_18546_59184# a_47186_59142# 0.35fF
C14832 pmat.rowoff_n[7] pmat.row_n[6] 0.34fF
C14833 a_22178_10496# ctopn 3.58fF
C14834 a_43262_57134# ctopp 3.57fF
C14835 pmat.en_bit_n[0] _1196_.B1 1.46fF
C14836 a_42258_71190# ctopp 3.40fF
C14837 VDD a_11902_56775# 0.49fF
C14838 a_29206_58138# ctopp 3.58fF
C14839 a_25190_68178# vcm 0.62fF
C14840 VDD result_out[11] 0.78fF
C14841 pmat.row_n[4] a_4257_34319# 2.06fF
C14842 VDD a_38242_58138# 0.52fF
C14843 a_21174_23548# a_21174_22544# 1.00fF
C14844 nmat.col[2] ctopn 1.97fF
C14845 VDD a_6975_76823# 1.37fF
C14846 a_18546_62196# a_20078_62154# 0.35fF
C14847 a_43262_71190# m2_43032_72014# 1.00fF
C14848 pmat.rowon_n[8] a_4523_21276# 0.57fF
C14849 a_20170_60146# a_21174_60146# 0.97fF
C14850 a_18546_60188# a_23090_60146# 0.35fF
C14851 nmat.col_n[21] vcm 3.39fF
C14852 VDD a_13919_65871# 0.58fF
C14853 VDD a_11842_59887# 0.53fF
C14854 a_6451_67655# pmat.rowoff_n[12] 0.66fF
C14855 VDD a_19928_37253# 1.01fF
C14856 nmat.col[31] a_13641_23439# 0.45fF
C14857 ANTENNA__1190__B1.DIODE nmat.col_n[7] 8.19fF
C14858 _1196_.B1 a_32405_32463# 1.57fF
C14859 m2_35000_7214# m3_35132_7346# 2.79fF
C14860 VDD a_39019_41001# 0.61fF
C14861 a_28202_68178# a_28202_67174# 1.00fF
C14862 a_30210_23548# vcm 0.65fF
C14863 a_21174_69182# ctopp 3.58fF
C14864 a_18162_58178# vcm 6.95fF
C14865 nmat.rowon_n[9] ctopn 1.40fF
C14866 a_32218_9492# vcm 0.65fF
C14867 VDD a_30210_69182# 0.52fF
C14868 a_18546_22542# a_49194_22950# 0.35fF
C14869 VDD a_27789_44743# 1.11fF
C14870 VDD a_18546_16518# 32.65fF
C14871 a_11232_73211# a_11271_73085# 0.46fF
C14872 _1194_.B1 nmat.col_n[21] 0.36fF
C14873 a_7717_14735# a_18241_31698# 0.37fF
C14874 _1183_.A2 nmat.col[12] 0.38fF
C14875 a_48282_20536# vcm 0.65fF
C14876 a_11007_58229# a_1957_43567# 0.43fF
C14877 a_30210_59142# ctopp 3.58fF
C14878 VDD nmat.col_n[20] 5.30fF
C14879 a_24186_11500# ctopn 3.58fF
C14880 VDD a_39939_29967# 0.71fF
C14881 VDD a_39246_59142# 0.52fF
C14882 pmat.col_n[26] ctopp 2.02fF
C14883 VDD a_17996_35303# 1.23fF
C14884 a_9075_28023# a_9441_20189# 0.49fF
C14885 ANTENNA__1197__B.DIODE a_11067_30287# 0.53fF
C14886 a_26194_16520# a_27198_16520# 0.97fF
C14887 a_18546_16518# a_35138_16926# 0.35fF
C14888 pmat.sw a_18563_27791# 1.02fF
C14889 m2_51064_54946# vcm 0.48fF
C14890 a_18546_67216# pmat.rowoff_n[11] 4.09fF
C14891 a_7415_29397# a_7840_27247# 0.55fF
C14892 a_28202_13508# vcm 0.65fF
C14893 m2_44036_7214# m2_45040_7214# 0.96fF
C14894 a_26194_18528# vcm 0.65fF
C14895 a_20475_49783# a_9411_2215# 0.77fF
C14896 a_2411_33749# a_4533_38279# 0.43fF
C14897 a_3339_59879# a_13183_72405# 0.71fF
C14898 a_2727_58470# a_1823_58237# 0.33fF
C14899 VDD a_11207_11079# 0.82fF
C14900 a_25879_31591# a_25695_28111# 3.80fF
C14901 a_18546_72236# a_29114_72194# 0.35fF
C14902 VDD m3_27100_72146# 0.40fF
C14903 a_37238_15516# vcm 0.65fF
C14904 VDD a_22178_17524# 0.52fF
C14905 a_4075_50087# a_2215_47375# 1.01fF
C14906 VDD a_2163_74173# 0.53fF
C14907 a_25879_31591# a_1781_9308# 0.66fF
C14908 m2_26968_72014# m3_27100_72146# 2.79fF
C14909 a_35230_70186# a_35230_69182# 1.00fF
C14910 VDD a_23182_8488# 0.55fF
C14911 a_19405_28853# a_21365_27247# 1.02fF
C14912 a_11317_36924# a_12069_36341# 1.15fF
C14913 a_18546_21538# a_26102_21946# 0.35fF
C14914 a_10239_14183# nmat.rowoff_n[3] 0.39fF
C14915 VDD a_6553_53047# 1.19fF
C14916 a_24186_14512# a_24186_13508# 1.00fF
C14917 nmat.col[26] vcm 8.88fF
C14918 pmat.rowon_n[0] nmat.rowon_n[2] 0.48fF
C14919 a_33222_23548# ctopn 3.40fF
C14920 VDD a_39246_19532# 0.52fF
C14921 pmat.row_n[6] pmat.rowon_n[6] 20.69fF
C14922 m2_17932_24282# m3_18064_24414# 2.79fF
C14923 a_35230_9492# ctopn 3.57fF
C14924 a_28202_57134# a_28202_56130# 1.00fF
C14925 ANTENNA__1197__A.DIODE a_19579_52789# 0.33fF
C14926 a_32218_19532# a_33222_19532# 0.97fF
C14927 VDD a_6970_67191# 0.71fF
C14928 a_33222_60146# vcm 0.62fF
C14929 VDD a_38242_10496# 0.52fF
C14930 a_2879_57487# a_2419_69455# 2.34fF
C14931 pmat.col_n[0] vcm 2.80fF
C14932 a_33423_47695# a_33515_31055# 0.57fF
C14933 VDD a_2124_65595# 0.67fF
C14934 VDD a_36234_55126# 0.58fF
C14935 a_18546_58180# a_45178_58138# 0.35fF
C14936 a_4951_76983# a_5047_76983# 0.33fF
C14937 pmat.row_n[8] nmat.rowon_n[4] 0.56fF
C14938 VDD a_8565_6037# 0.66fF
C14939 _1194_.B1 nmat.col[26] 3.50fF
C14940 a_31214_10496# a_32218_10496# 0.97fF
C14941 a_18546_10494# a_45178_10902# 0.35fF
C14942 a_2149_45717# a_1769_14735# 0.42fF
C14943 a_4719_30287# a_6553_53047# 0.56fF
C14944 a_45270_62154# ctopp 3.58fF
C14945 a_39246_16520# vcm 0.65fF
C14946 a_42258_56130# a_43262_56130# 0.97fF
C14947 a_18546_18526# a_18162_18528# 2.61fF
C14948 a_31214_13508# ctopn 3.58fF
C14949 a_40837_46261# a_7109_29423# 0.77fF
C14950 a_11921_37462# a_11149_36924# 0.37fF
C14951 a_18546_11498# a_20078_11906# 0.35fF
C14952 a_26194_57134# vcm 0.62fF
C14953 VDD a_30431_37683# 1.83fF
C14954 a_25190_71190# vcm 0.60fF
C14955 a_10949_42364# a_11297_36091# 0.69fF
C14956 a_1586_33927# cgen.dlycontrol1_in[2] 0.48fF
C14957 a_29206_18528# ctopn 3.58fF
C14958 a_35230_63158# pmat.col[16] 0.31fF
C14959 a_17842_27497# a_25575_31055# 0.43fF
C14960 a_8583_29199# a_7415_29397# 0.57fF
C14961 VDD a_5823_40303# 0.43fF
C14962 a_13459_28111# nmat.col_n[30] 0.89fF
C14963 _1187_.A2 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top 0.89fF
C14964 a_44266_70186# ctopp 3.57fF
C14965 a_26891_28327# ANTENNA__1183__B1.DIODE 1.19fF
C14966 a_30571_50959# a_45915_29941# 0.48fF
C14967 a_18243_28327# nmat.col_n[26] 0.91fF
C14968 a_40250_15516# ctopn 3.58fF
C14969 VDD a_3508_69135# 0.39fF
C14970 a_9411_2215# a_22307_27791# 0.47fF
C14971 VDD a_40250_11500# 0.52fF
C14972 a_14653_53458# a_16800_47213# 2.89fF
C14973 _1194_.B1 a_12263_50959# 0.74fF
C14974 a_13432_62581# pmat.row_n[8] 0.41fF
C14975 a_24186_22544# a_25190_22544# 0.97fF
C14976 pmat.rowon_n[11] nmat.rowoff_n[14] 0.32fF
C14977 a_47278_62154# a_48282_62154# 0.97fF
C14978 VDD m2_29980_54946# 0.62fF
C14979 a_45270_66170# a_46274_66170# 0.97fF
C14980 a_4351_55527# a_3345_62839# 0.65fF
C14981 _1154_.X inn_analog 0.47fF
C14982 a_18546_69224# a_40158_69182# 0.35fF
C14983 VDD a_27890_32143# 0.37fF
C14984 VDD a_18272_35077# 1.23fF
C14985 VDD pmat.col_n[19] 5.29fF
C14986 a_36265_48981# a_33467_46261# 0.35fF
C14987 a_10239_14183# a_10515_13967# 0.77fF
C14988 a_24867_53135# ANTENNA__1184__B1.DIODE 1.26fF
C14989 a_38242_63158# a_39246_63158# 0.97fF
C14990 a_1781_9308# config_1_in[15] 0.42fF
C14991 a_37238_22544# vcm 0.65fF
C14992 pmat.row_n[15] a_6173_22895# 2.51fF
C14993 pmat.row_n[4] pmat.rowon_n[4] 20.85fF
C14994 a_35230_68178# ctopp 3.58fF
C14995 VDD a_44266_68178# 0.52fF
C14996 a_13091_7655# a_12079_9615# 5.89fF
C14997 _1192_.A2 a_31675_47695# 1.29fF
C14998 a_4991_69831# a_11416_50363# 0.49fF
C14999 a_13091_28327# a_12461_29673# 1.22fF
C15000 a_30819_40191# a_11297_36091# 0.62fF
C15001 VDD a_16295_43177# 0.60fF
C15002 nmat.col[28] nmat.col_n[27] 6.58fF
C15003 nmat.col[20] nmat.col_n[20] 0.77fF
C15004 pmat.sw a_41731_49525# 1.84fF
C15005 m2_17932_16250# vcm 0.44fF
C15006 VDD a_9395_27791# 0.39fF
C15007 ANTENNA__1190__B1.DIODE ANTENNA__1190__A1.DIODE 0.56fF
C15008 a_9581_73487# a_10697_75218# 0.42fF
C15009 a_18546_20534# a_46182_20942# 0.35fF
C15010 a_42258_16520# ctopn 3.58fF
C15011 pmat.rowoff_n[4] a_12447_16143# 0.56fF
C15012 a_6830_22895# a_6173_22895# 0.71fF
C15013 a_14287_69455# a_10055_31591# 0.38fF
C15014 VDD m2_21948_7214# 0.93fF
C15015 VDD pmat.col[17] 4.51fF
C15016 pmat.rowon_n[8] a_3305_15823# 1.82fF
C15017 a_18546_62196# a_31122_62154# 0.35fF
C15018 pmat.rowon_n[9] vcm 0.58fF
C15019 a_3746_58487# a_2563_34837# 1.34fF
C15020 nmat.col_n[10] vcm 2.82fF
C15021 _1154_.A a_82863_64213# 0.40fF
C15022 a_18546_66212# a_27106_66170# 0.35fF
C15023 VDD a_49286_23548# 0.55fF
C15024 a_46274_70186# a_47278_70186# 0.97fF
C15025 VDD a_20170_66170# 0.52fF
C15026 a_33222_11500# a_34226_11500# 0.97fF
C15027 a_18546_11498# a_49194_11906# 0.35fF
C15028 VDD a_12585_37179# 1.13fF
C15029 vcm clk_ena 0.63fF
C15030 a_44266_56130# m2_44036_54946# 0.99fF
C15031 VDD nmat.col_n[5] 5.06fF
C15032 a_35230_64162# a_35230_63158# 1.00fF
C15033 a_13091_52047# a_11948_49783# 1.44fF
C15034 nmat.rowoff_n[3] ctopn 0.60fF
C15035 a_1923_53055# a_2163_55233# 0.35fF
C15036 VDD m2_17246_73620# 0.60fF
C15037 a_38242_10496# a_38242_9492# 1.00fF
C15038 a_18243_28327# a_24407_31375# 1.02fF
C15039 a_13091_28327# a_21739_29415# 0.77fF
C15040 a_19166_14512# ctopn 3.43fF
C15041 a_35230_58138# a_35230_57134# 1.00fF
C15042 VDD a_20170_10496# 0.52fF
C15043 VDD a_1757_38677# 0.62fF
C15044 a_9411_2215# ANTENNA__1183__B1.DIODE 0.70fF
C15045 VDD a_1927_43541# 0.42fF
C15046 a_45270_14512# vcm 0.65fF
C15047 cgen.dlycontrol2_in[4] a_10767_39087# 1.59fF
C15048 a_44266_64162# vcm 0.62fF
C15049 a_18241_31698# a_9963_28111# 0.64fF
C15050 a_39246_60146# a_39246_59142# 1.00fF
C15051 a_27198_18528# a_27198_17524# 1.00fF
C15052 _1194_.B1 clk_ena 0.71fF
C15053 ANTENNA_fanout52_A.DIODE a_24867_53135# 0.39fF
C15054 a_6283_31591# a_13275_48783# 1.49fF
C15055 VDD a_47278_13508# 0.52fF
C15056 pmat.rowon_n[11] nmat.rowoff_n[13] 0.36fF
C15057 a_40250_22544# ctopn 3.57fF
C15058 VDD a_45270_18528# 0.52fF
C15059 a_12263_50959# a_11067_49871# 0.37fF
C15060 a_27198_63158# a_27198_62154# 1.00fF
C15061 a_43262_67174# a_44266_67174# 0.97fF
C15062 pmat.row_n[4] ctopp 1.65fF
C15063 a_18546_70228# a_29114_70186# 0.35fF
C15064 cgen.dlycontrol3_in[3] a_14533_39631# 0.65fF
C15065 VDD vcm.sky130_fd_sc_hd__nand2_1_0.Y 0.42fF
C15066 m2_17932_69002# m2_17932_67998# 0.99fF
C15067 a_40250_66170# a_40250_65166# 1.00fF
C15068 a_33222_22544# a_33222_21540# 1.00fF
C15069 a_18546_14510# a_47186_14918# 0.35fF
C15070 a_32218_14512# a_33222_14512# 0.97fF
C15071 a_28202_62154# vcm 0.62fF
C15072 VDD pmat.rowoff_n[7] 18.08fF
C15073 nmat.col[24] nmat.col[28] 5.00fF
C15074 pmat.en_bit_n[2] _1187_.A2 2.72fF
C15075 a_11067_49871# a_21923_47919# 0.36fF
C15076 a_31214_64162# a_32218_64162# 0.97fF
C15077 a_18546_64204# a_45178_64162# 0.35fF
C15078 a_18546_17522# a_24094_17930# 0.35fF
C15079 a_32405_32463# a_45019_38645# 0.87fF
C15080 ANTENNA__1184__B1.DIODE a_38851_28327# 0.32fF
C15081 a_37238_68178# a_38242_68178# 0.97fF
C15082 VDD a_28078_29967# 0.32fF
C15083 pmat.rowon_n[0] a_5579_12394# 0.33fF
C15084 a_18975_40871# a_14533_39631# 0.50fF
C15085 pmat.rowon_n[11] vcm 0.85fF
C15086 a_13909_39605# a_14107_39958# 0.30fF
C15087 a_33222_8488# m2_32992_7214# 1.00fF
C15088 pmat.rowon_n[5] vcm 0.59fF
C15089 a_26194_13508# a_26194_12504# 1.00fF
C15090 VDD a_9579_26159# 0.38fF
C15091 a_18546_15514# a_24094_15922# 0.35fF
C15092 a_47278_65166# vcm 0.62fF
C15093 a_43262_60146# ctopp 3.58fF
C15094 VDD a_11299_31573# 0.86fF
C15095 VDD a_21087_36649# 0.63fF
C15096 a_27198_70186# vcm 0.62fF
C15097 a_2411_33749# a_5823_34863# 0.31fF
C15098 a_19166_22544# vcm 0.65fF
C15099 VDD a_8831_24501# 1.24fF
C15100 a_2648_29397# a_2564_21959# 0.53fF
C15101 a_21739_29415# a_17139_30503# 0.87fF
C15102 a_48282_14512# ctopn 3.58fF
C15103 pmat.row_n[7] a_3305_15823# 0.38fF
C15104 pmat.sample pmat.row_n[0] 0.40fF
C15105 VDD a_30140_43781# 1.22fF
C15106 a_2149_45717# a_1923_61759# 0.68fF
C15107 m2_17932_8218# m2_17932_7214# 0.99fF
C15108 pmat.col_n[26] m2_45040_54946# 0.42fF
C15109 a_6292_65479# a_5687_71829# 0.57fF
C15110 a_4351_55527# a_3339_70759# 0.93fF
C15111 a_18546_59184# a_40158_59142# 0.35fF
C15112 a_33222_65166# a_33222_64162# 1.00fF
C15113 a_36234_57134# ctopp 3.58fF
C15114 a_5081_53135# pmat.rowon_n[3] 0.81fF
C15115 a_35230_71190# ctopp 3.40fF
C15116 VDD a_45270_57134# 0.52fF
C15117 a_22178_58138# ctopp 3.58fF
C15118 VDD a_44266_71190# 0.55fF
C15119 VDD a_31214_58138# 0.52fF
C15120 a_42258_23548# a_43262_23548# 0.97fF
C15121 a_22178_16520# a_22178_15516# 1.00fF
C15122 _1154_.X clk_ena 0.40fF
C15123 VDD a_11067_30287# 12.02fF
C15124 a_44266_9492# a_45270_9492# 0.97fF
C15125 pmat.row_n[4] a_3746_58487# 0.51fF
C15126 a_9135_60967# a_2046_30184# 0.94fF
C15127 a_40837_46261# nmat.col_n[21] 0.67fF
C15128 VDD a_27887_41271# 0.60fF
C15129 a_18546_24550# a_45178_24958# 0.35fF
C15130 _1192_.B1 a_35244_32411# 0.49fF
C15131 VDD a_26957_39867# 1.35fF
C15132 nmat.col_n[11] m2_29980_24282# 0.37fF
C15133 a_1739_47893# cgen.dlycontrol4_in[0] 8.80fF
C15134 _1179_.X a_1781_9308# 2.44fF
C15135 a_23182_23548# vcm 0.65fF
C15136 nmat.col[19] nmat.col_n[19] 4.10fF
C15137 VDD a_23182_69182# 0.52fF
C15138 a_25190_9492# vcm 0.65fF
C15139 a_47278_61150# vcm 0.62fF
C15140 a_43262_23548# m2_43032_24282# 0.99fF
C15141 m2_51064_18258# a_50290_18528# 0.96fF
C15142 a_18546_22542# a_42166_22950# 0.35fF
C15143 VDD a_4215_15797# 0.42fF
C15144 a_41254_20536# vcm 0.65fF
C15145 a_34226_65166# a_35230_65166# 0.97fF
C15146 a_23182_59142# ctopp 3.58fF
C15147 VDD a_32218_59142# 0.52fF
C15148 a_11149_36924# a_14589_35286# 4.18fF
C15149 pmat.sw vcm 0.51fF
C15150 a_41254_21540# a_42258_21540# 0.97fF
C15151 VDD a_13653_35516# 1.42fF
C15152 VDD pmat.rowon_n[6] 3.58fF
C15153 cgen.dlycontrol4_in[3] a_11317_40188# 0.58fF
C15154 cgen.dlycontrol4_in[4] a_12197_43746# 4.06fF
C15155 a_18546_16518# a_28110_16926# 0.35fF
C15156 a_9643_66389# a_10921_64786# 0.37fF
C15157 a_42258_71190# a_42258_70186# 1.00fF
C15158 a_40105_47375# a_40741_46565# 0.35fF
C15159 VDD a_4421_67477# 0.43fF
C15160 VDD a_5731_58951# 2.15fF
C15161 a_4075_50087# a_2315_44124# 0.53fF
C15162 pmat.col_n[21] vcm 2.80fF
C15163 a_21174_13508# vcm 0.65fF
C15164 VDD a_11021_42619# 1.01fF
C15165 m2_37008_7214# m2_38012_7214# 0.96fF
C15166 a_7717_14735# a_37291_29397# 0.42fF
C15167 a_28704_29568# a_17842_27497# 0.38fF
C15168 pmat.sw _1194_.B1 0.45fF
C15169 a_18162_18528# vcm 6.95fF
C15170 a_24407_31375# a_30571_50959# 2.87fF
C15171 a_18162_56170# ctopp 1.18fF
C15172 VDD a_2051_29973# 0.65fF
C15173 a_1674_68047# a_3136_72515# 0.34fF
C15174 a_3615_71631# a_3936_70197# 0.60fF
C15175 ANTENNA__1195__A1.DIODE a_45277_32687# 0.42fF
C15176 a_40250_13508# a_41254_13508# 0.97fF
C15177 cgen.enable_dlycontrol_in a_12069_36341# 2.08fF
C15178 a_30210_15516# vcm 0.65fF
C15179 a_5687_71829# a_5357_62779# 0.77fF
C15180 VDD a_4505_74005# 0.75fF
C15181 nmat.rowon_n[15] a_18162_8488# 1.33fF
C15182 a_5731_58951# a_4719_30287# 1.86fF
C15183 a_11067_16359# a_12447_16143# 2.51fF
C15184 pmat.col_n[21] _1194_.B1 0.38fF
C15185 pmat.row_n[9] a_18546_65208# 0.35fF
C15186 a_11067_64015# a_4955_40277# 0.43fF
C15187 a_38242_18528# a_39246_18528# 0.97fF
C15188 a_10239_14183# a_2835_13077# 1.58fF
C15189 nmat.col_n[31] nmat.col[18] 1.81fF
C15190 VDD a_2163_71997# 0.51fF
C15191 a_25190_62154# a_25190_61150# 1.00fF
C15192 a_49286_12504# vcm 0.65fF
C15193 a_26194_23548# ctopn 3.40fF
C15194 VDD a_32218_19532# 0.52fF
C15195 a_28202_9492# ctopn 3.57fF
C15196 VDD m2_39016_72014# 1.38fF
C15197 nmat.col[29] nmat.col_n[18] 7.42fF
C15198 nmat.rowon_n[12] nmat.col_n[13] 3.13fF
C15199 a_26194_60146# vcm 0.62fF
C15200 VDD a_31214_10496# 0.52fF
C15201 a_1957_43567# a_2983_48071# 0.68fF
C15202 pmat.rowoff_n[7] a_1823_60949# 0.76fF
C15203 a_44266_20536# ctopn 3.58fF
C15204 VDD a_33395_43455# 0.77fF
C15205 a_10949_42364# a_11921_41814# 4.11fF
C15206 a_25190_15516# a_25190_14512# 1.00fF
C15207 a_49286_15516# a_50290_15516# 0.97fF
C15208 VDD _1192_.A2 20.27fF
C15209 VDD nmat.rowon_n[14] 14.12fF
C15210 pmat.sample_n a_11067_30287# 0.71fF
C15211 a_4383_7093# a_1586_8439# 0.40fF
C15212 a_27198_69182# a_27198_68178# 1.00fF
C15213 a_18546_57176# ctopp 1.58fF
C15214 a_18546_58180# a_38150_58138# 0.35fF
C15215 a_48282_69182# a_49286_69182# 0.97fF
C15216 ANTENNA__1190__B1.DIODE _0467_ 0.53fF
C15217 a_18546_10494# a_38150_10902# 0.35fF
C15218 a_35230_21540# a_35230_20536# 1.00fF
C15219 a_38242_62154# ctopp 3.58fF
C15220 VDD a_47278_62154# 0.52fF
C15221 a_24747_29967# a_28812_29575# 1.59fF
C15222 a_32218_16520# vcm 0.65fF
C15223 a_10873_39605# a_11113_39747# 1.73fF
C15224 VDD a_32871_49007# 0.46fF
C15225 a_11711_60751# a_12155_60751# 0.32fF
C15226 VDD a_9303_22351# 0.57fF
C15227 a_24186_13508# ctopn 3.58fF
C15228 ANTENNA__1183__B1.DIODE nmat.col[24] 0.56fF
C15229 a_22178_18528# ctopn 3.58fF
C15230 VDD a_21981_34191# 3.02fF
C15231 VDD a_4865_12533# 1.11fF
C15232 VDD a_11067_64015# 20.58fF
C15233 a_13091_52047# a_35786_47893# 0.62fF
C15234 a_21371_50087# a_30111_47911# 0.50fF
C15235 pmat.row_n[12] pmat.rowoff_n[11] 1.06fF
C15236 a_20170_10496# a_20170_9492# 1.00fF
C15237 a_37238_70186# ctopp 3.57fF
C15238 a_33222_15516# ctopn 3.58fF
C15239 VDD a_46274_70186# 0.52fF
C15240 a_6283_31591# a_1781_9308# 1.73fF
C15241 a_13643_29415# a_14379_6567# 1.01fF
C15242 a_21739_29415# a_9411_2215# 0.38fF
C15243 VDD a_33222_11500# 0.52fF
C15244 a_43720_32143# a_35244_32411# 0.51fF
C15245 a_46274_23548# a_46274_22544# 1.00fF
C15246 _1154_.X pmat.sw 2.62fF
C15247 a_6927_30503# a_8079_46519# 0.34fF
C15248 a_11041_39860# a_10767_39087# 0.45fF
C15249 a_11435_58791# nmat.rowoff_n[14] 1.11fF
C15250 VDD a_3339_59879# 11.25fF
C15251 a_45270_60146# a_46274_60146# 0.97fF
C15252 pmat.en_bit_n[0] a_22199_30287# 0.52fF
C15253 a_5651_66975# a_9827_53379# 0.61fF
C15254 a_18546_69224# a_33130_69182# 0.35fF
C15255 VDD a_25287_32117# 0.45fF
C15256 nmat.col_n[10] nmat.col_n[7] 0.95fF
C15257 a_12267_36694# a_12069_36341# 0.31fF
C15258 a_29206_11500# a_29206_10496# 1.00fF
C15259 a_48282_56130# vcm 0.62fF
C15260 pmat.sw a_42024_46805# 0.35fF
C15261 VDD a_1591_61519# 1.33fF
C15262 pmat.col[8] m2_26968_54946# 0.40fF
C15263 VDD a_3576_17143# 5.37fF
C15264 m2_48052_24282# m3_48184_24414# 2.79fF
C15265 a_30210_22544# vcm 0.65fF
C15266 a_34226_61150# a_35230_61150# 0.97fF
C15267 a_28202_68178# ctopp 3.58fF
C15268 a_2124_69947# a_2163_69821# 0.58fF
C15269 VDD a_37238_68178# 0.52fF
C15270 _1187_.A2 nmat.col_n[18] 5.44fF
C15271 a_11317_40188# a_11297_36091# 0.76fF
C15272 VDD a_11021_43011# 2.25fF
C15273 a_9963_13967# a_13091_18535# 2.56fF
C15274 a_44266_63158# vcm 0.62fF
C15275 a_28202_20536# a_29206_20536# 0.97fF
C15276 a_18546_20534# a_39154_20942# 0.35fF
C15277 a_35230_16520# ctopn 3.58fF
C15278 a_17154_43671# a_17902_43439# 0.37fF
C15279 VDD a_6292_69831# 2.69fF
C15280 a_18546_62196# a_24094_62154# 0.35fF
C15281 a_41254_67174# a_41254_66170# 1.00fF
C15282 a_27198_9492# a_27198_8488# 1.00fF
C15283 a_18546_21538# vcm 0.40fF
C15284 VDD a_42258_23548# 0.55fF
C15285 VDD a_44266_9492# 0.52fF
C15286 nmat.rowon_n[7] a_11948_49783# 1.10fF
C15287 a_18546_11498# a_42166_11906# 0.35fF
C15288 VDD a_28079_37737# 0.63fF
C15289 m2_40020_7214# m3_40152_7346# 2.79fF
C15290 a_28915_50959# _1183_.A2 0.47fF
C15291 a_15101_29423# a_9785_28879# 0.48fF
C15292 a_47147_44655# a_46968_45743# 0.30fF
C15293 a_40250_17524# a_41254_17524# 0.97fF
C15294 a_38242_57134# a_39246_57134# 0.97fF
C15295 a_11067_16359# a_11435_58791# 2.08fF
C15296 a_43262_20536# a_43262_19532# 1.00fF
C15297 a_37238_71190# a_38242_71190# 0.97fF
C15298 a_49286_67174# vcm 0.62fF
C15299 a_24186_58138# a_25190_58138# 0.97fF
C15300 a_38242_14512# vcm 0.65fF
C15301 _1187_.A2 a_42191_48071# 0.37fF
C15302 inp_analog ANTENNA__1395__A2.DIODE 4.77fF
C15303 a_18546_22542# nmat.rowoff_n[1] 4.09fF
C15304 a_37238_64162# vcm 0.62fF
C15305 VDD m2_43032_24282# 0.62fF
C15306 pmat.row_n[15] a_4979_38127# 3.15fF
C15307 VDD a_30833_46805# 0.61fF
C15308 a_41254_8488# a_42258_8488# 0.97fF
C15309 a_11041_38772# clk_ena 0.57fF
C15310 a_18546_58180# a_20078_58138# 0.35fF
C15311 VDD a_15435_29111# 0.70fF
C15312 a_13459_28111# a_41731_49525# 1.56fF
C15313 pmat.col_n[29] ctopp 2.02fF
C15314 VDD a_2944_56872# 1.10fF
C15315 ANTENNA__1187__B1.DIODE a_18243_28327# 6.80fF
C15316 VDD a_40250_13508# 0.52fF
C15317 a_11435_58791# nmat.rowoff_n[13] 0.36fF
C15318 a_49286_14512# a_49286_13508# 1.00fF
C15319 nmat.col_n[10] nmat.col_n[0] 2.17fF
C15320 a_1923_61759# a_4266_63303# 0.45fF
C15321 nmat.sw a_4703_24527# 0.49fF
C15322 a_33222_22544# ctopn 3.57fF
C15323 ANTENNA__1395__B1.DIODE _1183_.A2 2.80fF
C15324 VDD a_38242_18528# 0.52fF
C15325 m2_24960_24282# vcm 0.42fF
C15326 a_24186_61150# a_24186_60146# 1.00fF
C15327 nmat.col_n[14] vcm 2.80fF
C15328 a_4976_16091# a_7407_17455# 0.35fF
C15329 a_32218_19532# a_32218_18528# 1.00fF
C15330 a_18546_70228# a_22086_70186# 0.35fF
C15331 a_3339_59879# a_12723_64789# 0.58fF
C15332 pmat.rowoff_n[4] a_9528_20407# 1.66fF
C15333 a_13641_23439# nmat.en_C0_n 0.41fF
C15334 VDD a_49286_15516# 0.52fF
C15335 a_33309_41479# a_33765_41317# 0.40fF
C15336 a_18546_14510# a_40158_14918# 0.35fF
C15337 a_21174_62154# vcm 0.62fF
C15338 cgen.dlycontrol3_in[4] a_11497_40719# 1.09fF
C15339 VDD a_4613_19087# 1.28fF
C15340 a_18546_64204# a_38150_64162# 0.35fF
C15341 a_5462_62215# a_10286_60405# 0.34fF
C15342 ANTENNA__1196__A2.DIODE nmat.col_n[13] 0.30fF
C15343 VDD a_24747_29967# 6.43fF
C15344 a_19166_70186# ctopp 3.42fF
C15345 a_25190_59142# a_25190_58138# 1.00fF
C15346 a_18546_72236# a_32126_72194# 0.35fF
C15347 nmat.col_n[3] a_9528_20407# 0.55fF
C15348 VDD a_1757_26159# 0.60fF
C15349 _1224_.X _1179_.X 2.70fF
C15350 a_40250_65166# vcm 0.62fF
C15351 a_11041_38772# a_20534_35431# 1.14fF
C15352 a_47278_21540# vcm 0.65fF
C15353 a_36234_60146# ctopp 3.58fF
C15354 m2_31988_72014# m3_32120_72146# 2.79fF
C15355 VDD a_5963_32117# 0.43fF
C15356 VDD a_45270_60146# 0.52fF
C15357 VDD a_11041_36596# 2.14fF
C15358 a_20170_70186# vcm 0.62fF
C15359 a_11067_64015# pmat.rowoff_n[1] 0.74fF
C15360 a_45019_38645# a_40951_31599# 0.31fF
C15361 a_30210_17524# a_30210_16520# 1.00fF
C15362 a_11067_16359# a_7048_23277# 0.56fF
C15363 _1194_.A2 nmat.col_n[26] 0.93fF
C15364 a_1899_35051# cgen.dlycontrol4_in[0] 1.12fF
C15365 a_2952_25045# a_2683_22089# 1.05fF
C15366 m2_17932_57958# vcm 0.44fF
C15367 a_18546_19530# a_51202_19938# 0.35fF
C15368 a_3866_57399# a_4075_68583# 0.92fF
C15369 a_41254_14512# ctopn 3.58fF
C15370 VDD a_19166_68178# 0.56fF
C15371 a_36234_12504# a_37238_12504# 0.97fF
C15372 a_49286_22544# a_50290_22544# 0.97fF
C15373 a_1781_9308# a_22199_32149# 0.63fF
C15374 a_28131_50069# a_30663_50087# 1.85fF
C15375 pmat.rowon_n[3] a_1781_9308# 0.79fF
C15376 m2_17932_15246# m3_18064_15378# 2.76fF
C15377 pmat.col_n[22] m2_41024_54946# 0.37fF
C15378 a_18546_7482# a_20078_7890# 0.35fF
C15379 VDD a_4123_20693# 0.56fF
C15380 a_18546_59184# a_33130_59142# 0.35fF
C15381 a_25190_59142# a_26194_59142# 0.97fF
C15382 a_29206_57134# ctopp 3.57fF
C15383 a_28202_71190# ctopp 3.40fF
C15384 VDD pmat.col[15] 4.72fF
C15385 VDD a_38242_57134# 0.52fF
C15386 a_18546_20534# a_21082_20942# 0.35fF
C15387 VDD a_37238_71190# 0.55fF
C15388 a_24867_53135# a_17139_30503# 0.79fF
C15389 ANTENNA__1395__A1.DIODE a_28915_50959# 0.97fF
C15390 VDD a_24186_58138# 0.52fF
C15391 ANTENNA__1184__B1.DIODE a_13643_29415# 0.49fF
C15392 a_2263_43719# a_28455_47381# 1.04fF
C15393 pmat.rowon_n[5] pmat.rowoff_n[5] 20.79fF
C15394 VDD a_39111_38825# 0.61fF
C15395 a_10515_61839# a_13643_29415# 0.65fF
C15396 VDD a_45187_38129# 1.53fF
C15397 a_1591_61519# a_1823_60949# 0.42fF
C15398 a_1781_9308# a_2648_29397# 1.07fF
C15399 a_18546_64204# ctopp 1.59fF
C15400 VDD a_3325_40847# 1.13fF
C15401 ANTENNA__1190__B1.DIODE nmat.col[12] 1.61fF
C15402 a_27198_56130# m2_26968_54946# 0.99fF
C15403 a_18546_55168# a_49194_55126# 0.35fF
C15404 a_18546_24550# a_38150_24958# 0.35fF
C15405 a_12228_39605# a_12237_36596# 0.86fF
C15406 a_4399_51157# a_4257_34319# 0.39fF
C15407 a_2046_30184# a_2217_29973# 0.49fF
C15408 a_21174_68178# a_21174_67174# 1.00fF
C15409 a_2879_57487# a_4720_58487# 0.46fF
C15410 VDD a_12789_68021# 0.96fF
C15411 a_40250_61150# vcm 0.62fF
C15412 ANTENNA__1395__A1.DIODE ANTENNA__1395__B1.DIODE 1.85fF
C15413 a_18546_22542# a_35138_22950# 0.35fF
C15414 a_50290_21540# ctopn 3.43fF
C15415 VDD cgen.dlycontrol3_in[0] 9.86fF
C15416 a_20170_14512# vcm 0.65fF
C15417 VDD a_3571_13627# 5.80fF
C15418 a_19166_64162# vcm 0.61fF
C15419 VDD m2_39016_54946# 0.62fF
C15420 VDD a_5221_45199# 0.34fF
C15421 a_34226_20536# vcm 0.65fF
C15422 a_1674_68047# a_2791_57703# 1.84fF
C15423 a_5462_62215# a_6568_59887# 0.36fF
C15424 VDD a_49286_22544# 0.52fF
C15425 a_11113_39747# cgen.dlycontrol2_in[2] 1.55fF
C15426 pmat.rowoff_n[4] a_19541_28879# 1.09fF
C15427 VDD a_18597_31599# 1.49fF
C15428 a_25879_31591# a_31263_28309# 0.85fF
C15429 VDD a_18546_7482# 33.27fF
C15430 VDD a_25190_59142# 0.52fF
C15431 a_7026_24527# _0467_ 0.53fF
C15432 VDD cgen.dlycontrol1_in[1] 7.94fF
C15433 VDD pmat.col_n[22] 5.26fF
C15434 a_45370_48169# a_45450_48695# 0.48fF
C15435 _1194_.B1 a_45450_48695# 0.58fF
C15436 VDD a_22343_50613# 0.37fF
C15437 VDD a_4317_62215# 0.46fF
C15438 a_46274_17524# vcm 0.65fF
C15439 _1194_.A2 a_24407_31375# 0.73fF
C15440 VDD a_20170_18528# 0.52fF
C15441 m2_20944_54946# vcm 0.42fF
C15442 _1183_.A2 a_30111_47911# 0.99fF
C15443 _1192_.A2 a_7840_27247# 0.83fF
C15444 pmat.row_n[14] a_18162_70226# 25.58fF
C15445 a_47278_8488# vcm 0.64fF
C15446 VDD a_19611_27247# 0.60fF
C15447 a_4985_51433# a_4025_54965# 0.50fF
C15448 a_1781_9308# a_30412_31751# 0.42fF
C15449 VDD a_27785_43131# 1.16fF
C15450 nmat.rowoff_n[6] a_13655_26703# 0.46fF
C15451 nmat.col_n[19] nmat.col_n[29] 0.32fF
C15452 a_5363_33551# a_14452_51843# 0.60fF
C15453 m2_17932_12234# m3_18064_12366# 2.76fF
C15454 m2_29980_7214# m2_30984_7214# 0.96fF
C15455 pmat.col_n[27] pmat.col[27] 1.00fF
C15456 nmat.sw cgen.dlycontrol1_in[0] 2.10fF
C15457 a_18546_64204# a_20078_64162# 0.35fF
C15458 pmat.rowoff_n[12] ctopn 1.40fF
C15459 VDD a_8215_69929# 0.42fF
C15460 a_2411_43301# a_7479_53909# 0.56fF
C15461 VDD dummypin[4] 1.14fF
C15462 a_23182_15516# vcm 0.65fF
C15463 VDD a_9155_17455# 0.38fF
C15464 cgen.dlycontrol4_in[2] cgen.dlycontrol2_in[4] 1.30fF
C15465 VDD m2_51064_59966# 1.04fF
C15466 VDD a_2769_22357# 0.65fF
C15467 a_28202_70186# a_28202_69182# 1.00fF
C15468 ANTENNA__1187__B1.DIODE a_30571_50959# 0.55fF
C15469 a_24867_53135# a_26891_28327# 0.95fF
C15470 pmat.en_bit_n[2] nmat.col[30] 3.35fF
C15471 a_42258_12504# vcm 0.65fF
C15472 a_2419_69455# cgen.dlycontrol4_in[0] 0.42fF
C15473 a_47278_64162# ctopp 3.58fF
C15474 a_4865_12533# a_4895_12559# 0.46fF
C15475 a_18162_23548# ctopn 1.18fF
C15476 VDD a_25190_19532# 0.52fF
C15477 a_21174_9492# ctopn 3.57fF
C15478 VDD m2_24960_72014# 0.98fF
C15479 a_21174_57134# a_21174_56130# 1.00fF
C15480 a_4128_64391# a_11067_30287# 3.85fF
C15481 a_25190_19532# a_26194_19532# 0.97fF
C15482 VDD a_24186_10496# 0.52fF
C15483 a_37238_20536# ctopn 3.58fF
C15484 pmat.col[18] ctopp 1.98fF
C15485 a_50290_17524# m2_51064_17254# 0.96fF
C15486 a_18546_58180# a_31122_58138# 0.35fF
C15487 a_24186_10496# a_25190_10496# 0.97fF
C15488 a_18546_10494# a_31122_10902# 0.35fF
C15489 ANTENNA__1395__A2.DIODE ANTENNA__1395__B1.DIODE 1.13fF
C15490 a_49286_17524# ctopn 3.57fF
C15491 VDD a_19166_71190# 0.60fF
C15492 a_31214_62154# ctopp 3.58fF
C15493 a_22199_30287# nmat.col_n[24] 1.45fF
C15494 VDD a_40250_62154# 0.52fF
C15495 a_25190_16520# vcm 0.65fF
C15496 a_21174_62154# pmat.col[2] 0.31fF
C15497 pmat.rowon_n[8] a_3305_17999# 1.30fF
C15498 m2_48052_24282# vcm 0.42fF
C15499 a_50290_8488# ctopn 3.24fF
C15500 a_35230_56130# a_36234_56130# 0.97fF
C15501 VDD a_1591_23445# 0.41fF
C15502 VDD a_12969_40175# 1.15fF
C15503 nmat.col[31] a_42240_29423# 0.67fF
C15504 a_50290_65166# ctopp 3.43fF
C15505 a_2007_25597# a_12437_28585# 0.43fF
C15506 VDD a_10651_42035# 2.04fF
C15507 m2_17932_9222# m3_18064_9354# 2.76fF
C15508 a_18546_55168# a_32126_55126# 0.35fF
C15509 a_28704_29568# a_25575_31055# 0.40fF
C15510 a_1858_25615# a_12079_31061# 0.34fF
C15511 a_15667_27239# nmat.col[29] 1.24fF
C15512 a_30210_70186# ctopp 3.57fF
C15513 nmat.col[5] m2_23956_24282# 0.39fF
C15514 a_18975_40871# a_12345_39100# 0.32fF
C15515 a_26194_15516# ctopn 3.58fF
C15516 VDD a_39246_70186# 0.52fF
C15517 VDD a_26194_11500# 0.52fF
C15518 a_26194_23548# m2_25964_24282# 0.99fF
C15519 a_12585_39355# a_12197_38306# 0.32fF
C15520 a_10515_13967# a_5351_19913# 1.33fF
C15521 a_11948_49783# a_33839_46805# 0.36fF
C15522 a_1674_57711# a_4025_54965# 0.67fF
C15523 a_4128_64391# a_5731_58951# 0.73fF
C15524 a_11021_43011# a_12658_42895# 0.59fF
C15525 a_40250_62154# a_41254_62154# 0.97fF
C15526 a_47278_16520# a_47278_15516# 1.00fF
C15527 a_38242_66170# a_39246_66170# 0.97fF
C15528 a_45270_12504# ctopn 3.58fF
C15529 a_18546_69224# a_26102_69182# 0.35fF
C15530 VDD dummypin[2] 1.05fF
C15531 a_41254_56130# vcm 0.62fF
C15532 a_8491_47911# a_11435_58791# 1.56fF
C15533 a_23021_29199# a_19405_28853# 0.51fF
C15534 nmat.rowon_n[7] cgen.dlycontrol1_in[2] 0.47fF
C15535 a_22186_30485# a_15753_28879# 0.30fF
C15536 a_31214_63158# a_32218_63158# 0.97fF
C15537 a_18546_63200# a_45178_63158# 0.35fF
C15538 a_23182_22544# vcm 0.65fF
C15539 a_5535_57993# a_4843_54826# 0.93fF
C15540 a_21174_68178# ctopp 3.58fF
C15541 a_44266_66170# vcm 0.62fF
C15542 VDD a_30210_68178# 0.52fF
C15543 a_1923_31743# a_1591_26159# 0.34fF
C15544 a_12116_39783# a_11339_39319# 0.50fF
C15545 a_11883_62063# a_12199_62621# 0.37fF
C15546 pmat.col_n[1] vcm 2.79fF
C15547 a_10781_42869# a_11297_36091# 2.09fF
C15548 a_26891_28327# a_38851_28327# 3.26fF
C15549 VDD a_34593_43493# 1.39fF
C15550 VDD a_6853_14967# 1.03fF
C15551 a_12116_40871# a_12116_39783# 0.49fF
C15552 a_5363_33551# a_1781_9308# 1.21fF
C15553 a_37238_63158# vcm 0.62fF
C15554 VDD a_10049_60663# 2.73fF
C15555 ANTENNA__1196__A2.DIODE ANTENNA__1395__B1.DIODE 1.13fF
C15556 a_18546_10494# ctopn 1.59fF
C15557 pmat.rowoff_n[12] pmat.rowon_n[12] 20.66fF
C15558 VDD a_5423_30485# 0.50fF
C15559 _1183_.A2 nmat.col[18] 0.81fF
C15560 a_1769_13103# a_1769_14735# 12.87fF
C15561 a_18546_20534# a_32126_20942# 0.35fF
C15562 a_11317_36924# clk_ena 0.31fF
C15563 a_28202_16520# ctopn 3.58fF
C15564 pmat.row_n[11] cgen.dlycontrol4_in[5] 2.82fF
C15565 a_10515_15055# ANTENNA__1197__A.DIODE 0.48fF
C15566 VDD a_2099_76725# 0.62fF
C15567 pmat.row_n[9] vcm 1.15fF
C15568 m2_51064_21270# vcm 0.51fF
C15569 VDD a_35230_23548# 0.54fF
C15570 a_50290_61150# ctopp 3.43fF
C15571 _1154_.X a_13459_28111# 0.94fF
C15572 a_39246_70186# a_40250_70186# 0.97fF
C15573 VDD a_37238_9492# 0.52fF
C15574 a_18546_11498# a_35138_11906# 0.35fF
C15575 a_26194_11500# a_27198_11500# 0.97fF
C15576 VDD a_12311_19783# 0.41fF
C15577 a_28202_64162# a_28202_63158# 1.00fF
C15578 VDD a_35071_39913# 0.62fF
C15579 a_13459_28111# a_42024_46805# 0.68fF
C15580 a_31214_10496# a_31214_9492# 1.00fF
C15581 a_18546_71232# a_50198_71190# 0.35fF
C15582 a_42258_67174# vcm 0.62fF
C15583 a_28202_58138# a_28202_57134# 1.00fF
C15584 nmat.en_bit_n[1] a_16966_29673# 0.87fF
C15585 _1187_.A2 a_15667_27239# 0.37fF
C15586 VDD config_1_in[1] 1.02fF
C15587 VDD a_19689_44581# 1.17fF
C15588 a_31214_14512# vcm 0.65fF
C15589 a_6927_30503# a_8453_46287# 0.47fF
C15590 VDD a_3367_14906# 0.94fF
C15591 a_30210_64162# vcm 0.62fF
C15592 a_9963_13967# a_7717_14735# 3.07fF
C15593 a_32218_60146# a_32218_59142# 1.00fF
C15594 pmat.row_n[8] a_18162_64202# 25.57fF
C15595 pmat.col[2] m2_20944_54946# 0.39fF
C15596 a_2046_30184# a_5179_31591# 0.34fF
C15597 VDD a_24861_29673# 1.10fF
C15598 a_16800_47213# a_11948_49783# 0.59fF
C15599 a_11067_49871# a_12044_49641# 1.05fF
C15600 pmat.row_n[4] a_2564_21959# 0.92fF
C15601 m2_51064_63982# m2_51064_62978# 0.99fF
C15602 pmat.rowon_n[13] vcm 0.60fF
C15603 a_50290_62154# a_50290_61150# 1.00fF
C15604 VDD a_33222_13508# 0.52fF
C15605 nmat.rowon_n[7] a_2411_43301# 0.99fF
C15606 a_26194_22544# ctopn 3.57fF
C15607 VDD a_31214_18528# 0.52fF
C15608 a_20170_63158# a_20170_62154# 1.00fF
C15609 m2_44036_54946# vcm 0.42fF
C15610 pmat.row_n[10] pmat.rowon_n[10] 20.01fF
C15611 a_36234_67174# a_37238_67174# 0.97fF
C15612 a_11041_38772# a_12513_36924# 0.64fF
C15613 a_33222_66170# a_33222_65166# 1.00fF
C15614 a_26194_22544# a_26194_21540# 1.00fF
C15615 pmat.col_n[24] vcm 2.80fF
C15616 a_1781_9308# nmat.col_n[12] 0.80fF
C15617 VDD a_42258_15516# 0.52fF
C15618 a_1899_35051# a_2419_69455# 1.02fF
C15619 a_50290_15516# a_50290_14512# 1.00fF
C15620 a_25190_14512# a_26194_14512# 0.97fF
C15621 a_18546_14510# a_33130_14918# 0.35fF
C15622 nmat.col_n[10] _0467_ 0.58fF
C15623 a_24186_64162# a_25190_64162# 0.97fF
C15624 a_18546_64204# a_31122_64162# 0.35fF
C15625 a_20572_40517# a_20221_40835# 0.35fF
C15626 _1192_.B1 _1183_.A2 1.39fF
C15627 a_30210_68178# a_31214_68178# 0.97fF
C15628 pmat.row_n[15] pmat.row_n[14] 0.67fF
C15629 a_2419_53351# a_2419_69455# 1.12fF
C15630 VDD a_9777_26935# 0.75fF
C15631 VDD m2_51064_7214# 1.79fF
C15632 a_11067_30287# a_18241_31698# 0.77fF
C15633 a_6283_31591# a_31263_32117# 0.35fF
C15634 VDD a_18162_17524# 2.74fF
C15635 cgen.dlycontrol3_in[0] a_11113_40835# 1.79fF
C15636 VDD a_20411_51157# 0.34fF
C15637 a_33222_65166# vcm 0.62fF
C15638 a_11067_64015# cgen.dlycontrol4_in[4] 0.35fF
C15639 a_40250_21540# vcm 0.65fF
C15640 a_10378_7637# a_10747_6727# 0.33fF
C15641 VDD a_2099_21237# 0.38fF
C15642 a_29206_60146# ctopp 3.58fF
C15643 VDD a_5087_32687# 0.38fF
C15644 VDD a_38242_60146# 0.52fF
C15645 a_2952_25045# a_1586_18231# 0.55fF
C15646 VDD a_26041_36374# 1.12fF
C15647 VDD a_9279_71829# 0.79fF
C15648 a_18546_63200# ctopp 1.59fF
C15649 nmat.col[22] vcm 5.76fF
C15650 a_18546_19530# a_44174_19938# 0.35fF
C15651 m2_30984_54946# m2_31988_54946# 0.96fF
C15652 a_34226_14512# ctopn 3.58fF
C15653 VDD a_13575_68743# 0.34fF
C15654 a_18546_12502# a_48190_12910# 0.35fF
C15655 a_32687_46607# a_17842_27497# 0.47fF
C15656 VDD a_1586_33927# 4.51fF
C15657 VDD a_44266_16520# 0.52fF
C15658 a_19166_63158# vcm 0.61fF
C15659 pmat.col_n[18] m2_37008_54946# 0.38fF
C15660 a_18546_59184# a_26102_59142# 0.35fF
C15661 a_26194_65166# a_26194_64162# 1.00fF
C15662 a_1858_25615# a_4707_32156# 0.44fF
C15663 VDD pmat.en_bit_n[1] 0.78fF
C15664 a_22178_57134# ctopp 3.57fF
C15665 a_2695_76757# a_2861_76757# 0.46fF
C15666 a_21174_71190# ctopp 3.40fF
C15667 VDD a_31214_57134# 0.52fF
C15668 a_6451_67655# a_5595_65301# 0.93fF
C15669 VDD a_6007_33767# 3.58fF
C15670 ANTENNA__1195__A1.DIODE a_45866_38279# 0.87fF
C15671 pmat.sample pmat.row_n[3] 0.53fF
C15672 a_5779_71285# a_5081_53135# 0.67fF
C15673 a_47278_69182# vcm 0.62fF
C15674 a_33957_48437# a_35786_47893# 0.56fF
C15675 VDD a_30210_71190# 0.55fF
C15676 nmat.col_n[30] ctopn 2.03fF
C15677 a_18546_13506# a_20078_13914# 0.35fF
C15678 VDD a_5363_73807# 0.40fF
C15679 a_35230_23548# a_36234_23548# 0.97fF
C15680 a_29206_71190# m2_28976_72014# 1.00fF
C15681 VDD m2_17932_62978# 1.01fF
C15682 a_37238_9492# a_38242_9492# 0.97fF
C15683 a_14641_57167# a_14287_69455# 0.50fF
C15684 a_4719_30287# a_1586_33927# 0.88fF
C15685 a_44266_12504# a_44266_11500# 1.00fF
C15686 a_10873_38517# cgen.dlycontrol1_in[2] 0.38fF
C15687 VDD a_25393_38053# 1.30fF
C15688 VDD a_30523_41245# 1.52fF
C15689 a_1957_43567# a_12263_50959# 0.36fF
C15690 a_34705_51959# a_30663_50087# 1.58fF
C15691 a_18546_55168# a_42166_55126# 0.35fF
C15692 a_18546_24550# a_31122_24958# 0.35fF
C15693 pmat.row_n[5] nmat.col_n[10] 0.46fF
C15694 a_10873_38517# cgen.dlycontrol2_in[1] 1.24fF
C15695 VDD a_2163_55233# 0.47fF
C15696 a_4128_46983# a_4979_38127# 0.32fF
C15697 a_33222_61150# vcm 0.62fF
C15698 a_34226_62154# pmat.col[15] 0.31fF
C15699 a_18546_22542# a_28110_22950# 0.35fF
C15700 a_43262_21540# ctopn 3.58fF
C15701 a_12228_40693# a_23741_42567# 0.50fF
C15702 VDD a_12155_27791# 0.30fF
C15703 VDD a_38557_47381# 0.59fF
C15704 a_25879_31591# nmat.col[31] 0.38fF
C15705 a_27198_20536# vcm 0.65fF
C15706 a_21739_29415# a_25879_31591# 0.33fF
C15707 a_12228_39605# a_12513_39100# 2.05fF
C15708 a_27198_65166# a_28202_65166# 0.97fF
C15709 VDD a_42258_22544# 0.52fF
C15710 VDD a_32771_31599# 0.64fF
C15711 a_34226_21540# a_35230_21540# 0.97fF
C15712 VDD a_6763_13103# 0.40fF
C15713 a_47278_63158# ctopp 3.58fF
C15714 a_14365_22351# a_8443_20719# 2.02fF
C15715 pmat.col_n[1] pmat.col[2] 6.26fF
C15716 ANTENNA__1395__A1.DIODE _1192_.B1 6.35fF
C15717 a_13641_23439# a_20439_27247# 0.61fF
C15718 a_39246_17524# vcm 0.65fF
C15719 m2_18936_23278# m3_19068_23410# 2.76fF
C15720 m2_27972_24282# m2_28976_24282# 0.96fF
C15721 a_35230_71190# a_35230_70186# 1.00fF
C15722 a_40250_8488# vcm 0.64fF
C15723 _1179_.X ANTENNA__1183__B1.DIODE 0.39fF
C15724 a_49286_58138# a_50290_58138# 0.97fF
C15725 a_2564_21959# a_3305_27791# 0.41fF
C15726 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top nmat.col_n[30] 0.50fF
C15727 m2_22952_7214# m2_23956_7214# 0.96fF
C15728 VDD a_3351_27249# 2.65fF
C15729 _1194_.A2 ANTENNA__1187__B1.DIODE 2.03fF
C15730 m2_51064_70006# vcm 0.50fF
C15731 _1224_.X pmat.en_bit_n[2] 0.38fF
C15732 a_37820_30485# a_43720_32143# 0.63fF
C15733 VDD a_14287_70543# 8.23fF
C15734 a_33222_13508# a_34226_13508# 0.97fF
C15735 a_18546_13506# a_49194_13914# 0.35fF
C15736 VDD a_16311_28327# 8.32fF
C15737 VDD a_2149_45717# 16.12fF
C15738 a_48282_71190# m2_48052_72014# 1.00fF
C15739 VDD a_45502_48463# 0.32fF
C15740 a_49286_61150# a_49286_60146# 1.00fF
C15741 pmat.col_n[11] ANTENNA__1184__B1.DIODE 0.36fF
C15742 a_31214_18528# a_32218_18528# 0.97fF
C15743 a_18546_18526# a_45178_18934# 0.35fF
C15744 pmat.rowon_n[11] pmat.row_n[5] 6.09fF
C15745 pmat.row_n[5] pmat.rowon_n[5] 20.07fF
C15746 a_35230_12504# vcm 0.65fF
C15747 a_40250_64162# ctopp 3.58fF
C15748 a_6664_26159# a_4339_27804# 1.29fF
C15749 VDD a_50290_14512# 0.54fF
C15750 m2_45040_7214# m3_45172_7346# 2.79fF
C15751 m2_51064_9222# vcm 0.50fF
C15752 VDD a_49286_64162# 0.52fF
C15753 a_1781_9308# a_2021_9563# 0.72fF
C15754 a_12228_39605# a_17996_36391# 0.46fF
C15755 a_10055_31591# a_4075_31591# 0.55fF
C15756 a_1899_35051# cgen.dlycontrol4_in[3] 0.76fF
C15757 m2_22952_54946# m3_23084_55078# 2.79fF
C15758 a_50290_59142# a_50290_58138# 1.00fF
C15759 a_17842_27497# a_16965_27247# 0.32fF
C15760 pmat.sample pmat.row_n[1] 0.44fF
C15761 a_13091_28327# nmat.en_bit_n[0] 3.42fF
C15762 a_30210_20536# ctopn 3.58fF
C15763 VDD a_32219_44535# 0.60fF
C15764 a_10781_42364# a_14497_42658# 1.23fF
C15765 a_42258_15516# a_43262_15516# 0.97fF
C15766 VDD m2_51064_24282# 1.13fF
C15767 a_18546_58180# a_24094_58138# 0.35fF
C15768 a_20170_69182# a_20170_68178# 1.00fF
C15769 a_41254_69182# a_42258_69182# 0.97fF
C15770 a_18546_10494# a_24094_10902# 0.35fF
C15771 a_28202_21540# a_28202_20536# 1.00fF
C15772 VDD a_45107_34863# 0.50fF
C15773 a_42258_17524# ctopn 3.58fF
C15774 _1154_.A a_11067_30287# 0.48fF
C15775 a_24186_62154# ctopp 3.58fF
C15776 VDD a_33222_62154# 0.52fF
C15777 pmat.sw a_41443_28879# 0.34fF
C15778 a_43262_8488# ctopn 3.40fF
C15779 a_18546_56172# a_46182_56130# 0.35fF
C15780 VDD a_45178_24958# 0.44fF
C15781 pmat.row_n[2] a_18162_10496# 25.57fF
C15782 a_6664_26159# a_10223_26703# 0.30fF
C15783 a_13459_28111# nmat.col_n[0] 0.33fF
C15784 a_43262_65166# ctopp 3.58fF
C15785 VDD a_27913_42333# 1.10fF
C15786 a_18546_55168# a_25098_55126# 0.35fF
C15787 a_36234_24552# vcm 0.62fF
C15788 a_23182_70186# ctopp 3.57fF
C15789 VDD a_4123_52789# 0.35fF
C15790 a_18162_15516# ctopn 1.49fF
C15791 VDD a_32218_70186# 0.52fF
C15792 VDD a_18162_11500# 2.76fF
C15793 ANTENNA__1395__B1.DIODE a_2007_25597# 0.31fF
C15794 a_18546_72236# a_35138_72194# 0.35fF
C15795 a_10814_29111# a_11897_21263# 0.40fF
C15796 VDD m3_51196_69134# 0.34fF
C15797 a_39246_23548# a_39246_22544# 1.00fF
C15798 pmat.row_n[11] a_12263_50959# 0.62fF
C15799 _1187_.A2 a_11067_27239# 0.66fF
C15800 pmat.rowon_n[8] a_9963_13967# 0.36fF
C15801 a_38242_60146# a_39246_60146# 0.97fF
C15802 pmat.rowon_n[9] a_18162_65206# 1.19fF
C15803 a_18546_65208# a_19074_65166# 0.35fF
C15804 a_35244_32411# a_7717_14735# 0.71fF
C15805 m2_37008_72014# m3_37140_72146# 2.79fF
C15806 a_4075_31591# a_13688_47893# 0.35fF
C15807 a_38242_12504# ctopn 3.58fF
C15808 a_22178_11500# a_22178_10496# 1.00fF
C15809 a_34226_56130# vcm 0.62fF
C15810 VDD a_13779_36595# 1.43fF
C15811 VDD a_21082_72194# 0.32fF
C15812 a_6292_65479# a_6970_67191# 0.39fF
C15813 a_10515_13967# a_4383_7093# 1.33fF
C15814 a_38851_28327# nmat.col[24] 0.53fF
C15815 a_18546_63200# a_38150_63158# 0.35fF
C15816 a_30663_50087# a_37820_30485# 1.34fF
C15817 a_46274_68178# a_46274_67174# 1.00fF
C15818 a_18546_67216# a_19074_67174# 0.35fF
C15819 a_27198_61150# a_28202_61150# 0.97fF
C15820 pmat.rowoff_n[12] ctopp 0.60fF
C15821 nmat.rowon_n[12] a_5991_23983# 1.86fF
C15822 ANTENNA__1395__B1.DIODE a_19405_28853# 0.42fF
C15823 a_2791_57703# a_1823_68565# 0.47fF
C15824 a_37238_66170# vcm 0.62fF
C15825 VDD a_23182_68178# 0.52fF
C15826 ANTENNA__1395__A1.DIODE a_43720_32143# 2.54fF
C15827 a_13327_70741# a_14641_57167# 1.13fF
C15828 a_4075_50087# a_2419_69455# 0.41fF
C15829 m2_47048_72014# m2_48052_72014# 0.96fF
C15830 VDD a_20848_41605# 1.38fF
C15831 cgen.enable_dlycontrol_in clk_ena 0.55fF
C15832 a_30210_63158# vcm 0.62fF
C15833 VDD a_3751_64757# 0.74fF
C15834 pmat.sample ANTENNA__1195__A1.DIODE 1.30fF
C15835 VDD a_25315_28335# 1.67fF
C15836 a_1923_69823# a_7663_71317# 0.35fF
C15837 cgen.dlycontrol1_in[3] a_2953_33237# 0.59fF
C15838 VDD a_44174_55126# 0.42fF
C15839 a_18546_20534# a_25098_20942# 0.35fF
C15840 a_21174_20536# a_22178_20536# 0.97fF
C15841 a_21174_16520# ctopn 3.58fF
C15842 VDD a_3136_72515# 0.50fF
C15843 a_1591_43029# a_1757_43029# 0.72fF
C15844 a_44266_16520# a_45270_16520# 0.97fF
C15845 VDD cgen.dlycontrol3_in[3] 4.83fF
C15846 a_34226_67174# a_34226_66170# 1.00fF
C15847 VDD a_28202_23548# 0.55fF
C15848 VDD a_7521_47081# 2.85fF
C15849 a_43262_61150# ctopp 3.58fF
C15850 _1192_.B1 ANTENNA__1196__A2.DIODE 0.78fF
C15851 VDD a_30210_9492# 0.52fF
C15852 a_13357_37429# a_12237_36596# 4.51fF
C15853 a_18546_11498# a_28110_11906# 0.35fF
C15854 VDD a_4031_37191# 0.40fF
C15855 VDD a_19689_41317# 1.19fF
C15856 a_12447_16143# a_8305_20871# 0.46fF
C15857 pmat.row_n[0] nmat.rowon_n[12] 2.79fF
C15858 a_5351_19913# a_8861_24527# 0.37fF
C15859 a_12228_39605# a_14773_37218# 0.44fF
C15860 VDD a_46274_20536# 0.52fF
C15861 VDD a_18975_40871# 2.64fF
C15862 a_33222_17524# a_34226_17524# 0.97fF
C15863 VDD a_21124_39655# 1.13fF
C15864 a_31214_57134# a_32218_57134# 0.97fF
C15865 pmat.row_n[14] pmat.rowoff_n[2] 1.49fF
C15866 pmat.rowon_n[3] a_18546_11498# 4.09fF
C15867 a_13091_28327# pmat.col[20] 0.50fF
C15868 a_36234_20536# a_36234_19532# 1.00fF
C15869 a_2411_16101# a_6375_15279# 0.54fF
C15870 a_30210_71190# a_31214_71190# 0.97fF
C15871 a_18546_71232# a_43170_71190# 0.35fF
C15872 a_2727_58470# a_3838_70455# 0.50fF
C15873 a_35230_67174# vcm 0.62fF
C15874 _1192_.A2 nmat.col[15] 1.22fF
C15875 a_19541_28879# a_11823_46973# 0.63fF
C15876 VDD pmat.col[26] 4.52fF
C15877 ANTENNA__1190__B1.DIODE ANTENNA__1395__B1.DIODE 2.06fF
C15878 ANTENNA__1190__A1.DIODE a_13459_28111# 1.63fF
C15879 a_24591_28327# a_21739_29415# 0.60fF
C15880 VDD m3_51196_16382# 0.35fF
C15881 a_32687_46607# a_26479_32117# 0.49fF
C15882 cgen.enable_dlycontrol_in a_20534_35431# 1.61fF
C15883 a_24186_14512# vcm 0.65fF
C15884 a_4719_30287# cgen.dlycontrol3_in[3] 0.46fF
C15885 VDD a_14195_7351# 1.35fF
C15886 VDD nmat.en_bit_n[2] 0.58fF
C15887 a_23182_64162# vcm 0.62fF
C15888 a_18162_58178# pmat.row_n[2] 25.58fF
C15889 a_18546_8486# a_51202_8894# 0.35fF
C15890 a_34226_8488# a_35230_8488# 0.97fF
C15891 a_18546_65208# a_48190_65166# 0.35fF
C15892 VDD a_10747_6727# 0.39fF
C15893 a_22541_36603# a_22085_36374# 0.30fF
C15894 a_13091_18535# a_4533_38279# 0.95fF
C15895 VDD pmat.col_n[25] 5.08fF
C15896 VDD a_26194_13508# 0.52fF
C15897 pmat.col[29] ctopp 1.97fF
C15898 a_42258_14512# a_42258_13508# 1.00fF
C15899 VDD a_11711_62313# 0.42fF
C15900 a_2263_43719# a_33423_47695# 1.32fF
C15901 VDD a_24186_18528# 0.52fF
C15902 a_18546_67216# a_48190_67174# 0.35fF
C15903 a_46274_57134# a_46274_56130# 1.00fF
C15904 _1194_.B1 a_32405_32463# 2.12fF
C15905 a_25190_19532# a_25190_18528# 1.00fF
C15906 a_11391_69831# a_11487_69653# 0.36fF
C15907 nmat.col_n[26] m2_45040_24282# 0.44fF
C15908 a_5651_66975# a_6175_60039# 0.33fF
C15909 VDD a_39193_43131# 1.19fF
C15910 VDD a_35230_15516# 0.52fF
C15911 a_18546_14510# a_26102_14918# 0.35fF
C15912 a_29937_31055# a_46522_34293# 0.52fF
C15913 a_18546_7482# a_48190_7890# 0.35fF
C15914 a_18546_64204# a_24094_64162# 0.35fF
C15915 VDD a_45915_29941# 1.32fF
C15916 a_49286_10496# a_50290_10496# 0.97fF
C15917 a_33467_46261# a_45112_47607# 0.37fF
C15918 VDD a_3408_11849# 0.31fF
C15919 VDD m2_37008_7214# 0.91fF
C15920 pmat.col[12] ctopp 1.97fF
C15921 a_13503_43421# a_11021_43011# 1.19fF
C15922 VDD a_2747_74549# 0.42fF
C15923 a_26194_65166# vcm 0.62fF
C15924 VDD a_31152_48071# 1.62fF
C15925 a_33222_21540# vcm 0.65fF
C15926 pmat.rowon_n[10] ctopp 1.57fF
C15927 VDD a_10071_17999# 0.75fF
C15928 a_22178_60146# ctopp 3.58fF
C15929 a_20170_12504# ctopn 3.57fF
C15930 a_14287_70543# a_13718_68591# 0.53fF
C15931 VDD a_31214_60146# 0.52fF
C15932 a_21739_29415# a_43659_28853# 0.30fF
C15933 a_18243_28327# nmat.col_n[1] 0.47fF
C15934 a_48282_58138# vcm 0.62fF
C15935 a_49286_56130# m2_49056_54946# 0.99fF
C15936 nmat.col[11] vcm 5.76fF
C15937 nmat.col_n[12] comp_latch 2.07fF
C15938 pmat.sample pmat.row_n[7] 1.31fF
C15939 a_18546_63200# a_20078_63158# 0.35fF
C15940 a_23182_17524# a_23182_16520# 1.00fF
C15941 pmat.rowon_n[11] pmat.row_n[11] 20.55fF
C15942 _1179_.X nmat.col[31] 0.37fF
C15943 ANTENNA__1395__B1.DIODE a_7109_29423# 0.62fF
C15944 _1179_.X a_21739_29415# 5.70fF
C15945 pmat.rowon_n[5] a_18162_61190# 1.19fF
C15946 a_18546_61192# a_19074_61150# 0.35fF
C15947 a_18546_19530# a_37146_19938# 0.35fF
C15948 m2_23956_54946# m2_24960_54946# 0.96fF
C15949 a_19166_66170# vcm 0.61fF
C15950 a_27198_14512# ctopn 3.58fF
C15951 a_3339_70759# a_2411_43301# 1.96fF
C15952 a_6559_33767# a_4075_31591# 1.69fF
C15953 a_4025_54965# a_4243_54991# 0.40fF
C15954 a_18546_12502# a_41162_12910# 0.35fF
C15955 a_29206_12504# a_30210_12504# 0.97fF
C15956 a_42258_22544# a_43262_22544# 0.97fF
C15957 VDD a_27509_44219# 1.31fF
C15958 VDD a_37238_16520# 0.52fF
C15959 pmat.col[27] ctopp 1.97fF
C15960 a_30278_30511# a_32957_30287# 0.41fF
C15961 VDD a_1987_45370# 0.76fF
C15962 pmat.row_n[14] nmat.rowoff_n[0] 0.43fF
C15963 VDD a_27106_55126# 0.43fF
C15964 _1179_.X a_21215_48071# 0.34fF
C15965 VDD a_47186_7890# 0.34fF
C15966 pmat.col_n[1] ANTENNA__1190__A1.DIODE 0.31fF
C15967 VDD a_24186_57134# 0.52fF
C15968 _1196_.B1 _1187_.A2 0.49fF
C15969 pmat.row_n[15] pmat.rowon_n[15] 20.19fF
C15970 a_40250_69182# vcm 0.62fF
C15971 a_9411_2215# a_13643_29415# 1.64fF
C15972 VDD a_23182_71190# 0.55fF
C15973 a_19166_10496# vcm 0.65fF
C15974 VDD a_10443_12879# 0.36fF
C15975 pmat.col[8] vcm 5.88fF
C15976 _1154_.X pmat.en_bit_n[0] 0.41fF
C15977 pmat.sw nmat.col[12] 3.39fF
C15978 a_18546_23546# a_46182_23954# 0.35fF
C15979 a_11149_40188# cgen.dlycontrol4_in[0] 3.55fF
C15980 VDD a_6467_29415# 11.05fF
C15981 a_13091_7655# cgen.start_conv_in 0.41fF
C15982 a_18546_9490# a_50198_9898# 0.35fF
C15983 VDD a_5271_23447# 0.30fF
C15984 a_18162_55166# vcm 7.69fF
C15985 a_49286_59142# vcm 0.62fF
C15986 nmat.col[18] nmat.col_n[17] 6.77fF
C15987 VDD a_23884_40517# 1.22fF
C15988 pmat.rowoff_n[4] ctopn 1.40fF
C15989 a_18546_18526# ctopn 1.59fF
C15990 VDD a_17959_42089# 0.58fF
C15991 a_1957_43567# a_2389_45859# 0.45fF
C15992 pmat.row_n[2] a_12263_50959# 1.21fF
C15993 m2_17932_12234# vcm 0.44fF
C15994 VDD a_4266_63303# 0.58fF
C15995 VDD start_conversion_in 0.69fF
C15996 a_18546_24550# a_24094_24958# 0.35fF
C15997 nmat.col[24] nmat.col_n[19] 0.65fF
C15998 a_4399_51157# a_4313_44111# 0.33fF
C15999 a_44266_56130# ctopp 3.40fF
C16000 VDD a_13091_52047# 13.33fF
C16001 a_38242_8488# m2_38012_7214# 1.00fF
C16002 a_33423_47695# a_40105_47375# 0.33fF
C16003 a_26194_61150# vcm 0.62fF
C16004 a_2879_57487# a_2727_58470# 0.32fF
C16005 nmat.col_n[3] ctopn 2.02fF
C16006 a_36234_21540# ctopn 3.58fF
C16007 VDD a_47147_44655# 0.63fF
C16008 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top inn_analog 1.72fF
C16009 a_47278_66170# ctopp 3.58fF
C16010 VDD a_35230_22544# 0.52fF
C16011 VDD a_1643_58773# 0.38fF
C16012 VDD a_34924_36165# 1.28fF
C16013 a_40250_63158# ctopp 3.58fF
C16014 VDD a_49286_63158# 0.52fF
C16015 a_11041_38772# a_11113_38659# 0.62fF
C16016 a_32218_17524# vcm 0.65fF
C16017 a_2263_43719# a_6283_31591# 1.85fF
C16018 a_1586_8439# config_1_in[2] 0.51fF
C16019 a_25695_28111# a_29937_31055# 2.54fF
C16020 pmat.rowoff_n[8] _1194_.B1 0.71fF
C16021 a_18546_61192# a_48190_61150# 0.35fF
C16022 a_24867_53135# a_25879_31591# 0.63fF
C16023 ANTENNA__1395__A2.DIODE a_30663_50087# 0.36fF
C16024 VDD result_out[0] 0.71fF
C16025 m2_20944_24282# m2_21948_24282# 0.96fF
C16026 a_33222_8488# vcm 0.64fF
C16027 a_29937_31055# a_1781_9308# 0.84fF
C16028 pmat.rowon_n[8] a_4516_21531# 0.92fF
C16029 a_49286_19532# vcm 0.65fF
C16030 a_10515_15055# a_10515_61839# 1.87fF
C16031 a_45270_18528# a_45270_17524# 1.00fF
C16032 a_48282_10496# vcm 0.65fF
C16033 VDD result_out[9] 0.60fF
C16034 a_18546_13506# a_42166_13914# 0.35fF
C16035 pmat.row_n[4] a_4979_38127# 2.22fF
C16036 a_45270_63158# a_45270_62154# 1.00fF
C16037 pmat.rowon_n[3] a_2411_16101# 1.87fF
C16038 pmat.rowon_n[2] ctopp 1.57fF
C16039 a_45270_67174# ctopp 3.58fF
C16040 a_18546_18526# a_38150_18934# 0.35fF
C16041 a_21174_70186# a_21174_69182# 1.00fF
C16042 nmat.col_n[18] comp_latch 0.59fF
C16043 VDD a_22059_37683# 1.32fF
C16044 m2_17932_66994# m2_17932_65990# 0.99fF
C16045 a_2835_13077# a_4383_7093# 0.62fF
C16046 a_10190_60663# a_10195_59861# 0.35fF
C16047 a_10239_14183# a_11067_16359# 2.53fF
C16048 a_28202_12504# vcm 0.65fF
C16049 a_33222_64162# ctopp 3.58fF
C16050 VDD a_43262_14512# 0.52fF
C16051 pmat.row_n[10] a_18546_18526# 0.35fF
C16052 pmat.row_n[7] a_1923_31743# 0.58fF
C16053 VDD a_42258_64162# 0.52fF
C16054 a_2411_43301# a_6651_51733# 0.69fF
C16055 a_15667_27239# a_25695_28111# 0.79fF
C16056 a_24160_30199# a_22628_30485# 0.71fF
C16057 a_49286_64162# a_50290_64162# 0.97fF
C16058 nmat.col_n[19] m2_38012_24282# 0.40fF
C16059 _1196_.B1 pmat.col[1] 0.37fF
C16060 a_1674_57711# a_2124_56891# 0.46fF
C16061 a_13529_34951# clk_ena 0.78fF
C16062 nmat.rowon_n[10] ctopn 1.40fF
C16063 VDD a_18487_50069# 0.48fF
C16064 a_20170_12504# a_21174_12504# 0.97fF
C16065 a_44266_13508# a_44266_12504# 1.00fF
C16066 a_48282_23548# m2_48052_24282# 0.99fF
C16067 a_23182_20536# ctopn 3.58fF
C16068 VDD a_29404_44869# 1.31fF
C16069 m2_50060_54946# ctopp 0.69fF
C16070 a_19605_32149# a_18241_31698# 0.59fF
C16071 VDD a_18869_46831# 0.31fF
C16072 a_10239_14183# nmat.rowoff_n[13] 0.30fF
C16073 VDD nmat.col_n[26] 9.71fF
C16074 nmat.col[1] ctopn 1.92fF
C16075 a_20475_49783# a_19283_49783# 0.51fF
C16076 a_35230_17524# ctopn 3.58fF
C16077 a_50290_11500# vcm 0.65fF
C16078 nmat.en_bit_n[1] a_11067_30287# 0.41fF
C16079 a_11067_16359# a_9457_51163# 0.38fF
C16080 VDD a_26194_62154# 0.52fF
C16081 VDD m2_51064_14242# 1.01fF
C16082 cgen.dlycontrol4_in[4] a_1586_33927# 2.53fF
C16083 ANTENNA__1196__A2.DIODE a_30663_50087# 1.12fF
C16084 m2_17932_24282# vcm 0.42fF
C16085 a_36234_8488# ctopn 3.40fF
C16086 a_13432_62581# pmat.rowon_n[8] 2.11fF
C16087 a_28202_56130# a_29206_56130# 0.97fF
C16088 a_18546_56172# a_39154_56130# 0.35fF
C16089 VDD a_38150_24958# 0.44fF
C16090 pmat.rowon_n[0] a_2315_44124# 1.67fF
C16091 nmat.sw cgen.start_conv_in 0.37fF
C16092 VDD a_9135_60967# 7.29fF
C16093 a_1586_8439# a_3413_6037# 0.61fF
C16094 pmat.rowon_n[7] nmat.sw 0.82fF
C16095 a_6664_26159# a_11927_27399# 0.42fF
C16096 pmat.sample_n a_13091_52047# 1.59fF
C16097 pmat.col_n[27] vcm 2.80fF
C16098 a_36234_65166# ctopp 3.58fF
C16099 VDD a_13227_42333# 1.04fF
C16100 _1194_.A2 a_18243_28327# 1.04fF
C16101 VDD a_45270_65166# 0.52fF
C16102 a_50290_58138# m2_51064_57958# 0.96fF
C16103 a_11113_40835# a_18975_40871# 1.17fF
C16104 a_18546_68220# a_47186_68178# 0.35fF
C16105 VDD a_17702_29967# 1.01fF
C16106 VDD a_25190_70186# 0.52fF
C16107 _1183_.A2 a_10883_3303# 0.90fF
C16108 nmat.rowoff_n[14] ctopn 0.60fF
C16109 ANTENNA__1184__B1.DIODE nmat.col[19] 0.32fF
C16110 a_33222_62154# a_34226_62154# 0.97fF
C16111 a_40250_16520# a_40250_15516# 1.00fF
C16112 a_31214_66170# a_32218_66170# 0.97fF
C16113 a_36234_63158# pmat.col[17] 0.31fF
C16114 pmat.row_n[11] a_12447_16143# 3.04fF
C16115 a_11435_58791# a_1957_43567# 0.50fF
C16116 a_31214_12504# ctopn 3.58fF
C16117 VDD a_47499_32687# 0.41fF
C16118 a_27198_56130# vcm 0.62fF
C16119 VDD a_44757_37289# 1.09fF
C16120 VDD a_2791_57703# 9.48fF
C16121 a_15101_29423# nmat.col_n[3] 0.87fF
C16122 VDD a_7479_53909# 0.51fF
C16123 nmat.col_n[24] vcm 6.13fF
C16124 a_43720_32143# a_44966_43255# 0.43fF
C16125 pmat.row_n[13] a_18546_21538# 0.35fF
C16126 a_24186_63158# a_25190_63158# 0.97fF
C16127 a_18546_63200# a_31122_63158# 0.35fF
C16128 inp_analog clk_ena 16.85fF
C16129 a_50290_69182# ctopp 3.43fF
C16130 pmat.row_n[7] a_2935_38279# 0.64fF
C16131 a_30210_66170# vcm 0.62fF
C16132 VDD a_12597_68279# 0.62fF
C16133 a_13139_54599# a_12895_53359# 0.32fF
C16134 ANTENNA__1395__B1.DIODE nmat.col_n[21] 1.32fF
C16135 _1184_.A2 a_6664_26159# 2.48fF
C16136 m2_40020_72014# m2_41024_72014# 0.96fF
C16137 pmat.rowon_n[10] pmat.rowon_n[7] 0.32fF
C16138 a_9411_2215# a_20439_27247# 1.63fF
C16139 a_2407_49289# a_5081_53135# 0.61fF
C16140 a_23182_63158# vcm 0.62fF
C16141 a_10515_75895# a_5687_71829# 0.40fF
C16142 VDD a_24407_31375# 14.23fF
C16143 VDD a_37146_55126# 0.42fF
C16144 a_39246_63158# pmat.col[20] 0.31fF
C16145 pmat.sw _1519_.A 0.91fF
C16146 a_11927_27399# a_12061_26703# 0.71fF
C16147 pmat.rowoff_n[12] a_9427_50095# 0.34fF
C16148 VDD a_21174_23548# 0.55fF
C16149 VDD a_30913_38779# 1.25fF
C16150 a_36234_61150# ctopp 3.58fF
C16151 a_32218_70186# a_33222_70186# 0.97fF
C16152 VDD a_23182_9492# 0.52fF
C16153 VDD a_45270_61150# 0.52fF
C16154 a_11921_37462# a_11317_36924# 2.39fF
C16155 VDD a_34277_37462# 1.04fF
C16156 pmat.rowon_n[7] a_1858_25615# 1.00fF
C16157 ANTENNA__1197__A.DIODE a_17139_30503# 0.77fF
C16158 VDD a_39246_20536# 0.52fF
C16159 VDD a_5989_40303# 0.50fF
C16160 a_21174_64162# a_21174_63158# 1.00fF
C16161 a_24186_10496# a_24186_9492# 1.00fF
C16162 a_28202_67174# vcm 0.62fF
C16163 a_18546_71232# a_36142_71190# 0.35fF
C16164 a_21174_58138# a_21174_57134# 1.00fF
C16165 nmat.en_bit_n[1] _1192_.A2 1.06fF
C16166 a_9411_2215# a_6664_26159# 1.62fF
C16167 VDD m2_30984_54946# 0.62fF
C16168 a_40837_46261# a_32405_32463# 0.78fF
C16169 a_2983_48071# cgen.dlycontrol3_in[4] 0.41fF
C16170 a_18546_8486# a_44174_8894# 0.35fF
C16171 a_25190_60146# a_25190_59142# 1.00fF
C16172 a_18546_65208# a_41162_65166# 0.35fF
C16173 VDD a_32319_32143# 0.35fF
C16174 VDD a_20848_36165# 1.19fF
C16175 nmat.rowoff_n[13] ctopn 0.60fF
C16176 a_43262_62154# a_43262_61150# 1.00fF
C16177 VDD a_18162_13508# 2.74fF
C16178 cgen.dlycontrol3_in[4] a_12237_36596# 0.74fF
C16179 a_11435_58791# cgen.enable_dlycontrol_in 0.39fF
C16180 a_1717_13647# a_1761_11471# 0.38fF
C16181 ANTENNA__1190__B1.DIODE _1192_.B1 7.73fF
C16182 ANTENNA__1187__B1.DIODE ANTENNA__1197__B.DIODE 3.77fF
C16183 a_27001_30511# a_23021_29199# 0.52fF
C16184 _1194_.A2 a_18547_51565# 0.49fF
C16185 a_29206_67174# a_30210_67174# 0.97fF
C16186 a_18546_67216# a_41162_67174# 0.35fF
C16187 nmat.col_n[30] m2_49056_24282# 0.45fF
C16188 a_10055_31591# a_6283_31591# 0.56fF
C16189 a_34226_55126# m3_34128_55078# 2.08fF
C16190 a_3351_27249# a_3305_15823# 0.35fF
C16191 VDD a_7163_53333# 1.22fF
C16192 a_26194_66170# a_26194_65166# 1.00fF
C16193 a_18546_65208# ctopp 1.59fF
C16194 VDD a_28202_15516# 0.52fF
C16195 a_43262_15516# a_43262_14512# 1.00fF
C16196 nmat.rowoff_n[9] a_18546_14510# 4.09fF
C16197 VDD a_10814_29111# 1.13fF
C16198 a_18546_7482# a_41162_7890# 0.35fF
C16199 ANTENNA__1190__B1.DIODE a_23395_53135# 2.63fF
C16200 a_23182_68178# a_24186_68178# 0.97fF
C16201 a_45270_69182# a_45270_68178# 1.00fF
C16202 vcm ctopn 33.24fF
C16203 _1184_.A2 a_8197_20871# 0.34fF
C16204 VDD a_47278_12504# 0.52fF
C16205 ANTENNA__1187__B1.DIODE a_31675_47695# 0.66fF
C16206 a_9528_20407# a_8305_20871# 0.71fF
C16207 VDD m2_22952_7214# 1.26fF
C16208 a_30819_40191# cgen.dlycontrol2_in[4] 1.83fF
C16209 a_4523_21276# a_10071_17999# 0.73fF
C16210 cgen.dlycontrol3_in[1] a_12116_40871# 0.34fF
C16211 a_26194_21540# vcm 0.65fF
C16212 a_4991_69831# a_11435_58791# 0.44fF
C16213 VDD a_24186_60146# 0.52fF
C16214 a_3305_17999# a_3576_17143# 1.23fF
C16215 VDD dummypin[12] 0.99fF
C16216 a_41254_58138# vcm 0.62fF
C16217 m2_50060_7214# m3_50192_7346# 2.79fF
C16218 VDD nmat.col[6] 4.32fF
C16219 a_23821_35279# a_11041_36596# 0.51fF
C16220 m2_27972_54946# m3_28104_55078# 2.79fF
C16221 _1194_.A2 a_2046_30184# 1.66fF
C16222 a_18546_19530# a_30118_19938# 0.35fF
C16223 a_7521_47081# a_4128_64391# 1.68fF
C16224 a_18546_12502# a_34134_12910# 0.35fF
C16225 ANTENNA__1197__A.DIODE a_26891_28327# 0.44fF
C16226 VDD a_3983_43567# 0.40fF
C16227 VDD a_30210_16520# 0.52fF
C16228 a_26479_32117# a_24374_29941# 0.39fF
C16229 VDD a_17424_27497# 0.41fF
C16230 VDD pmat.en_C0_n 0.59fF
C16231 VDD a_17842_27497# 4.60fF
C16232 VDD a_40158_7890# 0.33fF
C16233 a_47278_11500# a_47278_10496# 1.00fF
C16234 m3_20072_24702# ctopn 0.35fF
C16235 _1179_.X a_24867_53135# 0.46fF
C16236 a_33222_69182# vcm 0.62fF
C16237 VDD a_12809_69679# 1.12fF
C16238 a_2215_47375# a_6559_57167# 0.58fF
C16239 a_2419_69455# a_5065_63669# 0.39fF
C16240 a_18546_23546# a_39154_23954# 0.35fF
C16241 a_28202_23548# a_29206_23548# 0.97fF
C16242 a_6448_5755# a_6487_5629# 0.76fF
C16243 pmat.sw inp_analog 3.37fF
C16244 a_1781_9308# cgen.dlycontrol4_in[1] 0.90fF
C16245 a_30210_9492# a_31214_9492# 0.97fF
C16246 a_18546_9490# a_43170_9898# 0.35fF
C16247 a_18546_61192# ctopp 1.59fF
C16248 a_4991_69831# a_10991_68591# 0.47fF
C16249 VDD a_18546_67216# 32.63fF
C16250 a_42258_59142# vcm 0.62fF
C16251 a_37238_12504# a_37238_11500# 1.00fF
C16252 pmat.row_n[6] pmat.rowoff_n[11] 0.69fF
C16253 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top vcm 138.49fF
C16254 VDD pmat.col[16] 4.59fF
C16255 VDD a_36801_42405# 1.25fF
C16256 VDD nmat.rowon_n[7] 19.41fF
C16257 a_1923_69823# a_1674_57711# 0.60fF
C16258 pmat.row_n[9] pmat.row_n[5] 1.40fF
C16259 a_37238_56130# ctopp 3.40fF
C16260 VDD a_46274_56130# 0.55fF
C16261 a_46274_20536# a_47278_20536# 0.97fF
C16262 a_18975_40871# a_20179_41046# 0.31fF
C16263 pmat.row_n[10] vcm 1.29fF
C16264 VDD a_14653_53458# 4.42fF
C16265 a_33957_48437# a_35540_46983# 0.36fF
C16266 a_18546_72236# a_38150_72194# 0.35fF
C16267 a_29206_21540# ctopn 3.58fF
C16268 a_45270_9492# a_45270_8488# 1.00fF
C16269 a_20170_65166# a_21174_65166# 0.97fF
C16270 VDD a_28202_22544# 0.52fF
C16271 a_40250_66170# ctopp 3.58fF
C16272 m2_42028_72014# m3_42160_72146# 2.79fF
C16273 VDD a_49286_66170# 0.52fF
C16274 VDD a_2655_59317# 0.40fF
C16275 a_14600_37607# a_26552_36165# 0.31fF
C16276 a_27198_21540# a_28202_21540# 0.97fF
C16277 VDD a_23700_36391# 1.16fF
C16278 VDD a_24094_72194# 0.32fF
C16279 pmat.rowoff_n[4] pmat.rowon_n[4] 20.95fF
C16280 nmat.rowon_n[7] a_4719_30287# 1.33fF
C16281 a_33222_63158# ctopp 3.58fF
C16282 a_5081_53135# a_6568_59887# 0.55fF
C16283 VDD a_42258_63158# 0.52fF
C16284 a_25190_17524# vcm 0.65fF
C16285 a_5558_9527# a_5654_9527# 0.79fF
C16286 a_18546_61192# a_41162_61150# 0.35fF
C16287 a_20170_55126# m3_20072_55078# 2.44fF
C16288 m2_47048_54946# m2_48052_54946# 0.96fF
C16289 a_28202_71190# a_28202_70186# 1.00fF
C16290 a_26194_8488# vcm 0.64fF
C16291 a_31105_46805# a_30833_46805# 0.48fF
C16292 a_42258_58138# a_43262_58138# 0.97fF
C16293 VDD nmat.rowoff_n[11] 2.38fF
C16294 pmat.col_n[0] pmat.row_n[8] 0.31fF
C16295 VDD a_10569_64489# 0.63fF
C16296 _1187_.A2 nmat.sw 0.30fF
C16297 a_42258_19532# vcm 0.65fF
C16298 _1192_.A2 a_19584_52423# 0.46fF
C16299 a_1674_57711# a_1586_63927# 0.94fF
C16300 pmat.rowon_n[12] vcm 0.61fF
C16301 a_50290_9492# m2_51064_9222# 0.96fF
C16302 a_41254_10496# vcm 0.65fF
C16303 a_18546_13506# a_35138_13914# 0.35fF
C16304 a_26194_13508# a_27198_13508# 0.97fF
C16305 a_5687_71829# a_3866_57399# 1.68fF
C16306 a_12197_43746# a_11497_40719# 0.71fF
C16307 a_42258_61150# a_42258_60146# 1.00fF
C16308 a_38242_67174# ctopp 3.58fF
C16309 a_18546_18526# a_31122_18934# 0.35fF
C16310 a_24186_18528# a_25190_18528# 0.97fF
C16311 a_50290_19532# a_50290_18528# 1.00fF
C16312 a_7109_29423# a_46027_44905# 0.43fF
C16313 VDD a_47278_67174# 0.52fF
C16314 VDD a_8841_60405# 0.60fF
C16315 ANTENNA__1183__B1.DIODE nmat.col_n[18] 2.09fF
C16316 pmat.en_bit_n[2] nmat.col[31] 0.39fF
C16317 a_21174_12504# vcm 0.65fF
C16318 pmat.en_bit_n[2] a_21739_29415# 1.23fF
C16319 a_26194_64162# ctopp 3.58fF
C16320 VDD a_36234_14512# 0.52fF
C16321 a_32218_56130# m2_31988_54946# 0.99fF
C16322 ANTENNA__1196__A2.DIODE a_10883_3303# 2.22fF
C16323 VDD a_35230_64162# 0.52fF
C16324 pmat.en_bit_n[2] a_20310_28029# 0.33fF
C16325 VDD a_21621_40955# 1.38fF
C16326 pmat.rowoff_n[15] a_12263_50959# 0.50fF
C16327 a_18546_57176# a_49194_57134# 0.35fF
C16328 a_43262_59142# a_43262_58138# 1.00fF
C16329 a_3688_17179# a_3576_17143# 0.56fF
C16330 ANTENNA__1190__A1.DIODE nmat.col[11] 0.30fF
C16331 a_33839_46805# a_35540_46983# 0.41fF
C16332 a_15667_27239# nmat.col_n[15] 0.38fF
C16333 VDD a_2847_50069# 0.47fF
C16334 a_35230_15516# a_36234_15516# 0.97fF
C16335 VDD m2_20944_24282# 0.61fF
C16336 a_34226_69182# a_35230_69182# 0.97fF
C16337 cgen.dlycontrol2_in[0] cgen.dlycontrol1_in[2] 1.25fF
C16338 a_1586_18231# a_1757_20181# 0.61fF
C16339 a_21174_21540# a_21174_20536# 1.00fF
C16340 VDD a_11921_35286# 2.16fF
C16341 a_28202_17524# ctopn 3.58fF
C16342 VDD pmat.col_n[28] 5.26fF
C16343 a_43262_11500# vcm 0.65fF
C16344 pmat.rowoff_n[4] ctopp 0.60fF
C16345 a_10873_40693# clk_ena 0.38fF
C16346 a_6787_47607# a_11435_58791# 0.61fF
C16347 a_18546_23546# a_21082_23954# 0.35fF
C16348 cgen.dlycontrol4_in[3] a_11149_40188# 0.39fF
C16349 a_48282_17524# a_48282_16520# 1.00fF
C16350 a_12309_38659# a_38711_37683# 0.31fF
C16351 a_29206_8488# ctopn 3.40fF
C16352 a_10883_3303# a_11337_25071# 1.04fF
C16353 cgen.dlycontrol2_in[1] cgen.dlycontrol2_in[0] 1.33fF
C16354 a_7109_29423# a_43720_32143# 1.12fF
C16355 a_18546_56172# a_32126_56130# 0.35fF
C16356 VDD a_31122_24958# 0.44fF
C16357 m2_44036_24282# m2_45040_24282# 0.96fF
C16358 VDD a_5307_67655# 2.04fF
C16359 VDD a_6583_61519# 0.49fF
C16360 a_31675_47695# a_25575_31055# 0.56fF
C16361 a_45270_19532# ctopn 3.58fF
C16362 a_29206_65166# ctopp 3.58fF
C16363 nmat.col[27] nmat.col_n[27] 0.86fF
C16364 a_17842_27497# nmat.col[20] 0.63fF
C16365 VDD a_38242_65166# 0.52fF
C16366 a_19166_18528# vcm 0.65fF
C16367 VDD a_45270_21540# 0.52fF
C16368 pmat.row_n[14] a_18546_22542# 0.35fF
C16369 a_43262_59142# a_44266_59142# 0.97fF
C16370 nmat.sample a_2007_25597# 0.42fF
C16371 a_44266_10496# ctopn 3.58fF
C16372 a_18546_68220# a_40158_68178# 0.35fF
C16373 a_2411_16101# a_1586_8439# 0.51fF
C16374 a_47278_68178# vcm 0.62fF
C16375 pmat.row_n[12] pmat.row_n[6] 0.74fF
C16376 a_32218_23548# a_32218_22544# 1.00fF
C16377 a_6283_31591# a_25688_32117# 0.42fF
C16378 a_31095_42367# a_24833_40719# 0.77fF
C16379 a_17902_43439# a_10949_43124# 0.41fF
C16380 cgen.dlycontrol3_in[1] a_28116_39655# 0.32fF
C16381 VDD a_1769_13103# 4.98fF
C16382 VDD a_4351_55527# 7.82fF
C16383 pmat.row_n[7] a_18546_15514# 0.35fF
C16384 a_9135_60967# a_8583_29199# 0.62fF
C16385 a_31214_60146# a_32218_60146# 0.97fF
C16386 a_18546_60188# a_45178_60146# 0.35fF
C16387 pmat.row_n[9] a_18162_65206# 25.57fF
C16388 a_24186_12504# ctopn 3.58fF
C16389 a_20170_56130# vcm 0.62fF
C16390 pmat.rowoff_n[12] a_2564_21959# 0.63fF
C16391 a_18546_21538# a_18162_21540# 2.61fF
C16392 cgen.dlycontrol3_in[2] config_2_in[12] 0.45fF
C16393 pmat.row_n[13] pmat.row_n[9] 1.96fF
C16394 a_15101_29423# a_22186_30485# 0.55fF
C16395 a_22628_30485# a_15753_28879# 0.69fF
C16396 a_18546_63200# a_24094_63158# 0.35fF
C16397 VDD m2_40020_72014# 1.11fF
C16398 a_39246_68178# a_39246_67174# 1.00fF
C16399 a_20170_61150# a_21174_61150# 0.97fF
C16400 a_43262_69182# ctopp 3.58fF
C16401 a_23182_66170# vcm 0.62fF
C16402 a_12263_50959# a_15899_47939# 0.42fF
C16403 ANTENNA__1395__A2.DIODE a_10589_22351# 0.39fF
C16404 m2_32992_72014# m2_33996_72014# 0.96fF
C16405 pmat.rowoff_n[15] clk_ena 0.66fF
C16406 VDD a_10873_38517# 8.03fF
C16407 VDD a_44733_44431# 0.57fF
C16408 m2_51064_17254# m3_51196_17386# 2.76fF
C16409 VDD a_14825_50095# 0.89fF
C16410 a_46274_11500# ctopn 3.58fF
C16411 a_18162_57174# ctopp 1.47fF
C16412 VDD a_13335_31359# 0.43fF
C16413 VDD a_10090_58093# 1.00fF
C16414 a_50290_20536# m2_51064_20266# 0.96fF
C16415 VDD a_13801_34427# 1.20fF
C16416 _1192_.B1 nmat.col_n[21] 0.44fF
C16417 cgen.enable_dlycontrol_in a_11921_37462# 0.38fF
C16418 a_37238_16520# a_38242_16520# 0.97fF
C16419 a_2215_47375# a_5784_52423# 1.22fF
C16420 VDD a_33957_48437# 1.83fF
C16421 a_27198_67174# a_27198_66170# 1.00fF
C16422 VDD a_7693_22365# 3.24fF
C16423 VDD ANTENNA__1187__B1.DIODE 22.52fF
C16424 a_29206_61150# ctopp 3.58fF
C16425 pmat.row_n[13] pmat.rowon_n[13] 20.11fF
C16426 VDD a_38242_61150# 0.52fF
C16427 VDD a_29163_38545# 1.00fF
C16428 a_13357_37429# a_24015_36911# 0.78fF
C16429 VDD a_14773_38306# 2.69fF
C16430 a_18546_71232# vcm 0.39fF
C16431 a_50290_13508# vcm 0.65fF
C16432 a_15435_29111# a_14691_29575# 0.35fF
C16433 VDD nmat.rowoff_n[9] 2.58fF
C16434 VDD a_12199_62621# 0.66fF
C16435 a_48282_18528# vcm 0.65fF
C16436 VDD a_32218_20536# 0.52fF
C16437 a_26194_17524# a_27198_17524# 0.97fF
C16438 pmat.row_n[1] pmat.rowon_n[1] 20.07fF
C16439 a_24186_57134# a_25190_57134# 0.97fF
C16440 pmat.col[30] m2_49056_54946# 0.39fF
C16441 a_29206_20536# a_29206_19532# 1.00fF
C16442 a_21174_67174# vcm 0.62fF
C16443 a_18546_71232# a_29114_71190# 0.35fF
C16444 a_23182_71190# a_24186_71190# 0.97fF
C16445 a_1674_68047# a_3267_74817# 0.48fF
C16446 a_31214_23548# m2_30984_24282# 0.99fF
C16447 a_11711_12565# a_11877_12565# 0.61fF
C16448 pmat.row_n[11] pmat.row_n[9] 4.91fF
C16449 nmat.col_n[7] ctopn 2.02fF
C16450 a_4128_64391# a_9135_60967# 3.22fF
C16451 VDD a_46797_45993# 0.54fF
C16452 pmat.row_n[3] nmat.rowon_n[12] 20.17fF
C16453 VDD a_44266_17524# 0.52fF
C16454 a_27198_8488# a_28202_8488# 0.97fF
C16455 a_18546_8486# a_37146_8894# 0.35fF
C16456 VDD a_10811_77437# 0.45fF
C16457 a_18546_65208# a_34134_65166# 0.35fF
C16458 VDD a_26479_32117# 1.28fF
C16459 a_46274_70186# a_46274_69182# 1.00fF
C16460 VDD a_45270_8488# 0.55fF
C16461 a_10873_36341# a_12069_36341# 0.40fF
C16462 a_18546_21538# a_48190_21946# 0.35fF
C16463 a_3615_71631# a_12003_52815# 0.40fF
C16464 a_35230_14512# a_35230_13508# 1.00fF
C16465 VDD a_3345_62839# 3.08fF
C16466 a_18546_67216# a_34134_67174# 0.35fF
C16467 a_39246_57134# a_39246_56130# 1.00fF
C16468 a_4075_68583# a_5341_59317# 0.37fF
C16469 VDD a_12147_24233# 0.35fF
C16470 ANTENNA__1196__A2.DIODE a_10589_22351# 0.88fF
C16471 a_43262_19532# a_44266_19532# 0.97fF
C16472 a_17842_27497# a_7840_27247# 0.31fF
C16473 nmat.col_n[9] m2_27972_24282# 0.37fF
C16474 a_11149_40188# a_11297_36091# 0.54fF
C16475 a_9963_13967# nmat.rowon_n[14] 3.02fF
C16476 VDD a_21174_15516# 0.52fF
C16477 m2_51064_14242# m3_51196_14374# 2.76fF
C16478 pmat.col_n[20] pmat.col[20] 0.79fF
C16479 a_18546_7482# a_34134_7890# 0.35fF
C16480 a_12069_36341# cgen.dlycontrol1_in[3] 0.54fF
C16481 a_42258_10496# a_43262_10496# 0.97fF
C16482 VDD a_9103_56383# 0.47fF
C16483 VDD a_3936_70197# 0.63fF
C16484 VDD a_40250_12504# 0.52fF
C16485 a_1899_35051# a_4843_54826# 0.31fF
C16486 VDD a_82815_54965# 0.48fF
C16487 VDD a_10245_51335# 0.41fF
C16488 VDD a_33839_46805# 1.22fF
C16489 _1224_.X a_11067_27239# 1.23fF
C16490 VDD pmat.rowoff_n[11] 2.81fF
C16491 a_48282_57134# vcm 0.62fF
C16492 VDD a_30765_37692# 1.21fF
C16493 a_47278_71190# vcm 0.60fF
C16494 a_11067_64015# a_9963_13967# 0.43fF
C16495 a_10055_31591# a_5363_33551# 2.21fF
C16496 a_34226_58138# vcm 0.62fF
C16497 a_50290_56130# m2_51064_55950# 0.96fF
C16498 a_12463_22351# a_11159_23145# 0.53fF
C16499 nmat.col[22] m2_41024_24282# 0.39fF
C16500 nmat.col_n[25] nmat.col[25] 0.83fF
C16501 a_18546_19530# a_23090_19938# 0.35fF
C16502 pmat.rowon_n[4] vcm 0.58fF
C16503 a_17139_30503# nmat.col[19] 1.35fF
C16504 VDD a_46211_50095# 0.48fF
C16505 a_22178_12504# a_23182_12504# 0.97fF
C16506 a_18546_12502# a_27106_12910# 0.35fF
C16507 a_35230_22544# a_36234_22544# 0.97fF
C16508 a_4259_73807# a_5211_57172# 0.34fF
C16509 VDD a_23182_16520# 0.52fF
C16510 VDD m2_44036_24282# 0.62fF
C16511 nmat.col_n[0] ctopn 1.81fF
C16512 VDD nmat.rowon_n[5] 8.34fF
C16513 VDD a_33130_7890# 0.33fF
C16514 ANTENNA__1197__B.DIODE a_18243_28327# 0.48fF
C16515 ANTENNA__1184__B1.DIODE a_13091_28327# 1.29fF
C16516 a_26194_69182# vcm 0.62fF
C16517 a_11067_16359# a_7779_22583# 1.17fF
C16518 a_18546_23546# a_32126_23954# 0.35fF
C16519 a_49286_63158# a_50290_63158# 0.97fF
C16520 m2_25964_24282# vcm 0.42fF
C16521 a_18546_9490# a_36142_9898# 0.35fF
C16522 nmat.col[14] vcm 5.76fF
C16523 a_10055_31591# a_4128_46983# 1.27fF
C16524 a_35230_59142# vcm 0.62fF
C16525 a_13641_23439# a_10223_26703# 0.46fF
C16526 a_13459_28111# nmat.col_n[4] 0.33fF
C16527 a_2411_16101# a_2879_19093# 0.38fF
C16528 pmat.col_n[30] vcm 2.81fF
C16529 a_50290_11500# m2_51064_11230# 0.96fF
C16530 m2_51064_11230# m3_51196_11362# 2.76fF
C16531 pmat.rowon_n[7] pmat.rowoff_n[4] 5.28fF
C16532 a_1586_33927# config_2_in[6] 0.36fF
C16533 a_30210_56130# ctopp 3.40fF
C16534 VDD a_28715_28879# 0.50fF
C16535 a_7658_71543# a_4075_50087# 0.65fF
C16536 pmat.rowoff_n[7] nmat.rowon_n[4] 1.10fF
C16537 VDD a_39246_56130# 0.55fF
C16538 VDD pmat.col[3] 5.93fF
C16539 a_1781_9308# a_2835_13077# 1.03fF
C16540 VDD m3_44168_72146# 0.33fF
C16541 a_22178_21540# ctopn 3.58fF
C16542 a_18546_66212# a_49194_66170# 0.35fF
C16543 cgen.dlycontrol3_in[1] a_1757_40853# 0.53fF
C16544 VDD a_21174_22544# 0.52fF
C16545 a_33222_66170# ctopp 3.58fF
C16546 _1192_.B1 a_44635_46025# 0.35fF
C16547 VDD a_5179_31591# 2.07fF
C16548 VDD a_42258_66170# 0.52fF
C16549 a_12237_36596# a_10873_36341# 0.50fF
C16550 a_44266_11500# a_45270_11500# 0.97fF
C16551 VDD a_3615_71631# 9.80fF
C16552 a_26194_63158# ctopp 3.58fF
C16553 a_15753_28879# a_8443_20719# 0.54fF
C16554 VDD a_16800_47213# 7.11fF
C16555 a_5363_70543# a_10049_60663# 0.86fF
C16556 VDD a_35230_63158# 0.52fF
C16557 a_46274_64162# a_46274_63158# 1.00fF
C16558 m2_23956_24282# m3_24088_24414# 2.79fF
C16559 a_49286_10496# a_49286_9492# 1.00fF
C16560 a_18546_61192# a_34134_61150# 0.35fF
C16561 m2_40020_54946# m2_41024_54946# 0.96fF
C16562 a_18162_8488# vcm 6.95fF
C16563 a_46274_58138# a_46274_57134# 1.00fF
C16564 vcm ctopp 33.24fF
C16565 a_19166_22544# m2_17932_22274# 0.96fF
C16566 VDD a_2952_25045# 5.32fF
C16567 a_35230_19532# vcm 0.65fF
C16568 a_50290_60146# a_50290_59142# 1.00fF
C16569 a_38242_18528# a_38242_17524# 1.00fF
C16570 VDD a_25575_31055# 2.56fF
C16571 a_19166_20536# a_20170_20536# 0.97fF
C16572 m2_51064_61974# m2_51064_60970# 0.99fF
C16573 _1192_.B1 nmat.col_n[10] 3.36fF
C16574 ANTENNA__1184__B1.DIODE a_17139_30503# 0.63fF
C16575 a_34226_10496# vcm 0.65fF
C16576 a_18546_13506# a_28110_13914# 0.35fF
C16577 a_11067_16359# a_5351_19913# 0.77fF
C16578 VDD a_3339_70759# 9.03fF
C16579 a_2263_43719# a_28621_47381# 0.52fF
C16580 cgen.dlycontrol4_in[1] cgen.dlycontrol4_in[2] 1.31fF
C16581 a_38242_63158# a_38242_62154# 1.00fF
C16582 a_34226_71190# m2_33996_72014# 1.00fF
C16583 _1192_.B1 clk_ena 0.66fF
C16584 VDD a_36936_49257# 0.41fF
C16585 pmat.rowon_n[4] a_18162_60186# 1.19fF
C16586 a_31214_67174# ctopp 3.58fF
C16587 a_18546_18526# a_24094_18934# 0.35fF
C16588 a_18546_70228# a_51202_70186# 0.35fF
C16589 VDD a_40250_67174# 0.52fF
C16590 _1192_.A2 a_18823_50247# 0.45fF
C16591 a_44266_22544# a_44266_21540# 1.00fF
C16592 VDD a_29206_14512# 0.52fF
C16593 a_43262_14512# a_44266_14512# 0.97fF
C16594 a_50290_62154# vcm 0.62fF
C16595 VDD a_28202_64162# 0.52fF
C16596 m2_51064_8218# m3_51196_8350# 2.76fF
C16597 a_9307_31068# nmat.col[10] 0.45fF
C16598 a_11067_49871# a_29076_48695# 0.32fF
C16599 VDD a_13653_40956# 1.35fF
C16600 a_42258_64162# a_43262_64162# 0.97fF
C16601 a_18546_17522# a_46182_17930# 0.35fF
C16602 a_48282_68178# a_49286_68178# 0.97fF
C16603 a_18546_57176# a_42166_57134# 0.35fF
C16604 a_23395_53135# clk_ena 1.32fF
C16605 a_4399_51157# a_4979_38127# 0.45fF
C16606 VDD pmat.row_n[12] 18.15fF
C16607 a_37238_13508# a_37238_12504# 1.00fF
C16608 VDD a_11785_16367# 0.66fF
C16609 pmat.en_bit_n[2] a_24867_53135# 0.67fF
C16610 VDD a_20583_28529# 0.37fF
C16611 a_18546_15514# a_46182_15922# 0.35fF
C16612 VDD m2_40020_54946# 0.62fF
C16613 a_11067_64015# a_18823_50247# 0.50fF
C16614 VDD a_42791_32375# 0.57fF
C16615 a_30663_50087# nmat.col_n[21] 1.19fF
C16616 VDD a_19074_7890# 0.34fF
C16617 a_11803_49551# a_11067_49871# 0.35fF
C16618 a_49286_70186# vcm 0.62fF
C16619 a_21174_17524# ctopn 3.58fF
C16620 a_36234_11500# vcm 0.65fF
C16621 pmat.col[10] ctopp 1.97fF
C16622 _1224_.X _1196_.B1 5.07fF
C16623 VDD pmat.col[5] 4.62fF
C16624 VDD a_4520_60975# 0.44fF
C16625 a_22178_8488# ctopn 3.40fF
C16626 m2_21948_54946# vcm 0.42fF
C16627 a_13091_18535# cgen.dlycontrol4_in[5] 1.88fF
C16628 a_21174_56130# a_22178_56130# 0.97fF
C16629 a_18546_56172# a_25098_56130# 0.35fF
C16630 VDD a_24094_24958# 0.44fF
C16631 m2_37008_24282# m2_38012_24282# 0.96fF
C16632 pmat.rowoff_n[14] a_18546_70228# 4.09fF
C16633 a_9135_69679# a_9301_69679# 0.39fF
C16634 a_29159_37607# a_11681_35823# 0.56fF
C16635 a_17139_30503# a_19439_30511# 0.63fF
C16636 pmat.row_n[9] nmat.rowoff_n[6] 1.43fF
C16637 a_38242_19532# ctopn 3.58fF
C16638 a_1899_35051# pmat.rowon_n[0] 1.00fF
C16639 a_22178_65166# ctopp 3.58fF
C16640 VDD a_28907_43177# 0.64fF
C16641 VDD a_31214_65166# 0.52fF
C16642 VDD a_38242_21540# 0.52fF
C16643 a_44266_65166# a_44266_64162# 1.00fF
C16644 a_10781_42869# ndecision_finish 0.64fF
C16645 a_37238_10496# ctopn 3.58fF
C16646 a_18546_68220# a_33130_68178# 0.35fF
C16647 a_2149_45717# a_6292_65479# 0.91fF
C16648 pmat.row_n[12] nmat.rowoff_n[2] 0.54fF
C16649 ANTENNA__1190__A1.DIODE vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top 0.40fF
C16650 a_44266_58138# ctopp 3.58fF
C16651 a_40250_68178# vcm 0.62fF
C16652 VDD a_9135_69679# 0.40fF
C16653 VDD a_2683_22089# 4.50fF
C16654 VDD a_14287_17455# 0.38fF
C16655 a_33222_16520# a_33222_15516# 1.00fF
C16656 a_26194_62154# a_27198_62154# 0.97fF
C16657 VDD m2_17932_58962# 1.12fF
C16658 a_24186_66170# a_25190_66170# 0.97fF
C16659 a_18546_60188# a_38150_60146# 0.35fF
C16660 a_18162_60186# ctopp 1.49fF
C16661 ANTENNA__1184__B1.DIODE a_26891_28327# 1.74fF
C16662 ANTENNA__1197__B.DIODE a_30571_50959# 0.39fF
C16663 a_32687_46607# a_44444_32233# 1.20fF
C16664 pmat.rowoff_n[8] pmat.row_n[5] 0.53fF
C16665 a_3325_20175# a_7048_23277# 0.49fF
C16666 a_28704_29568# a_28812_29575# 0.91fF
C16667 m2_32992_54946# m3_33124_55078# 2.79fF
C16668 VDD m2_25964_72014# 1.00fF
C16669 a_45270_23548# vcm 0.65fF
C16670 a_36234_69182# ctopp 3.58fF
C16671 a_47278_9492# vcm 0.65fF
C16672 a_33986_47375# a_35186_47375# 0.53fF
C16673 VDD a_45270_69182# 0.52fF
C16674 a_3351_27249# a_3305_17999# 1.52fF
C16675 m2_25964_72014# m2_26968_72014# 0.96fF
C16676 a_33423_47695# nmat.en_bit_n[0] 0.34fF
C16677 _1192_.A2 a_35244_32411# 0.65fF
C16678 VDD a_6651_51733# 0.49fF
C16679 a_26194_62154# pmat.col[7] 0.31fF
C16680 a_45270_65166# a_46274_65166# 0.97fF
C16681 a_45270_59142# ctopp 3.58fF
C16682 a_4383_7093# a_7436_16519# 0.30fF
C16683 a_39246_11500# ctopn 3.58fF
C16684 VDD a_2957_58255# 0.88fF
C16685 a_11317_36924# cgen.dlycontrol1_in[0] 2.55fF
C16686 m3_35132_24990# ctopn 0.31fF
C16687 VDD a_15107_34743# 0.62fF
C16688 ANTENNA__1395__A2.DIODE ANTENNA__1195__A1.DIODE 0.41fF
C16689 ANTENNA__1184__B1.DIODE _1184_.A2 17.56fF
C16690 a_4075_50087# a_4843_54826# 1.10fF
C16691 a_2419_53351# a_2727_58470# 1.05fF
C16692 a_18546_16518# a_50198_16926# 0.35fF
C16693 m2_49056_24282# vcm 0.41fF
C16694 a_22178_61150# ctopp 3.58fF
C16695 a_18546_55168# vcm 0.37fF
C16696 nmat.rowoff_n[8] ctopn 0.60fF
C16697 a_25190_70186# a_26194_70186# 0.97fF
C16698 VDD a_31214_61150# 0.52fF
C16699 VDD a_13985_40229# 1.40fF
C16700 pmat.rowon_n[8] a_18162_64202# 1.19fF
C16701 a_43262_13508# vcm 0.65fF
C16702 VDD a_10591_42089# 0.57fF
C16703 VDD a_2439_13889# 0.56fF
C16704 nmat.rowoff_n[10] a_18546_13506# 4.09fF
C16705 nmat.rowoff_n[14] nmat.rowoff_n[1] 0.46fF
C16706 a_41254_18528# vcm 0.65fF
C16707 a_22499_49783# a_33957_48437# 0.67fF
C16708 VDD a_25190_20536# 0.52fF
C16709 cgen.start_conv_in clk_dig 2.74fF
C16710 m2_51064_65990# vcm 0.50fF
C16711 VDD a_83196_3561# 0.66fF
C16712 VDD dummypin[8] 0.99fF
C16713 a_10239_14183# a_8305_20871# 0.32fF
C16714 a_12513_39100# a_11497_38543# 3.32fF
C16715 a_18546_71232# a_22086_71190# 0.35fF
C16716 a_6200_70919# a_5497_73719# 0.36fF
C16717 VDD a_5123_52423# 0.60fF
C16718 a_18546_72236# a_41162_72194# 0.35fF
C16719 a_1823_68565# a_1823_64213# 0.55fF
C16720 VDD a_37238_17524# 0.52fF
C16721 pmat.sw _1192_.B1 0.91fF
C16722 a_1739_47893# a_1775_35113# 0.37fF
C16723 VDD a_23823_47679# 0.51fF
C16724 a_18546_8486# a_30118_8894# 0.35fF
C16725 a_18546_65208# a_27106_65166# 0.35fF
C16726 m2_47048_72014# m3_47180_72146# 2.79fF
C16727 a_49286_18528# a_50290_18528# 0.97fF
C16728 VDD a_38242_8488# 0.55fF
C16729 a_18546_21538# a_41162_21946# 0.35fF
C16730 VDD a_28247_34191# 0.72fF
C16731 pmat.rowoff_n[12] a_1895_26372# 0.34fF
C16732 VDD a_27106_72194# 0.33fF
C16733 a_36234_62154# a_36234_61150# 1.00fF
C16734 pmat.col[2] ctopp 1.98fF
C16735 ANTENNA__1184__B1.DIODE a_9411_2215# 7.50fF
C16736 a_48282_23548# ctopn 3.40fF
C16737 VDD a_6343_18517# 0.36fF
C16738 a_50290_9492# ctopn 3.42fF
C16739 a_22178_67174# a_23182_67174# 0.97fF
C16740 a_18546_67216# a_27106_67174# 0.35fF
C16741 a_6787_47607# a_11203_62037# 0.89fF
C16742 a_4351_55527# a_4128_64391# 0.32fF
C16743 a_2419_69455# pmat.rowon_n[0] 3.02fF
C16744 a_48282_60146# vcm 0.62fF
C16745 nmat.col[13] nmat.col[19] 0.51fF
C16746 VDD a_82971_11989# 0.35fF
C16747 a_12116_39783# a_12585_40443# 0.73fF
C16748 a_10767_39087# a_11339_39319# 1.24fF
C16749 nmat.sw a_1781_9308# 0.59fF
C16750 a_20170_19532# ctopn 3.57fF
C16751 VDD a_7085_15055# 0.37fF
C16752 a_10873_40693# a_29217_41570# 0.54fF
C16753 a_36234_15516# a_36234_14512# 1.00fF
C16754 VDD a_11521_64239# 0.54fF
C16755 VDD a_26355_29673# 0.41fF
C16756 a_18546_7482# a_27106_7890# 0.35fF
C16757 VDD a_20170_21540# 0.52fF
C16758 ANTENNA__1196__A2.DIODE ANTENNA__1195__A1.DIODE 8.99fF
C16759 a_13459_28111# ANTENNA__1395__B1.DIODE 0.85fF
C16760 a_38242_69182# a_38242_68178# 1.00fF
C16761 a_41731_49525# nmat.col[29] 1.97fF
C16762 a_46274_21540# a_46274_20536# 1.00fF
C16763 ANTENNA__1197__A.DIODE a_25879_31591# 6.02fF
C16764 VDD a_33222_12504# 0.52fF
C16765 a_19166_13508# m2_17932_13238# 0.96fF
C16766 nmat.col_n[2] m2_20944_24282# 0.37fF
C16767 VDD a_18243_28327# 9.11fF
C16768 cgen.dlycontrol4_in[2] a_17902_43439# 1.21fF
C16769 VDD a_2999_76922# 0.85fF
C16770 pmat.row_n[5] a_10239_14183# 0.38fF
C16771 pmat.rowon_n[7] vcm 0.62fF
C16772 m2_17932_20266# vcm 0.44fF
C16773 a_18546_60188# a_20078_60146# 0.35fF
C16774 a_46274_13508# ctopn 3.58fF
C16775 nmat.col_n[7] m2_25964_24282# 0.37fF
C16776 a_14719_37737# a_13503_36893# 0.45fF
C16777 a_41254_57134# vcm 0.62fF
C16778 a_40250_71190# vcm 0.60fF
C16779 a_44266_18528# ctopn 3.58fF
C16780 a_27198_58138# vcm 0.62fF
C16781 VDD a_5087_19319# 0.32fF
C16782 VDD a_13909_39605# 4.26fF
C16783 VDD a_38972_39655# 1.14fF
C16784 a_10515_15055# nmat.rowon_n[13] 0.91fF
C16785 nmat.col_n[16] nmat.col[17] 6.87fF
C16786 a_18546_69224# ctopp 1.59fF
C16787 a_2411_16101# a_3063_14741# 0.34fF
C16788 a_2879_57487# a_3770_57399# 0.61fF
C16789 a_2727_58470# a_2419_69455# 0.94fF
C16790 a_18546_12502# a_19074_12910# 0.35fF
C16791 VDD m3_31116_7346# 0.37fF
C16792 VDD config_1_in[9] 1.00fF
C16793 VDD a_17867_44535# 0.64fF
C16794 a_7717_14735# a_2007_25597# 0.94fF
C16795 nmat.col[1] a_4383_7093# 0.34fF
C16796 a_1591_58799# a_1823_58237# 0.44fF
C16797 a_20170_18528# a_20170_17524# 1.00fF
C16798 pmat.row_n[12] a_13718_68591# 0.39fF
C16799 VDD a_28704_29568# 5.00fF
C16800 a_5081_53135# a_1586_63927# 0.51fF
C16801 VDD a_26102_7890# 0.33fF
C16802 a_40250_11500# a_40250_10496# 1.00fF
C16803 VDD pmat.col_n[31] 5.42fF
C16804 a_14365_22351# a_10589_22351# 0.48fF
C16805 a_1923_61759# a_1591_63701# 0.37fF
C16806 a_18546_23546# a_25098_23954# 0.35fF
C16807 a_21174_23548# a_22178_23548# 0.97fF
C16808 m2_45040_54946# vcm 0.42fF
C16809 a_23182_9492# a_24186_9492# 0.97fF
C16810 a_18546_9490# a_29114_9898# 0.35fF
C16811 a_45270_61150# a_46274_61150# 0.97fF
C16812 a_50290_68178# ctopp 3.43fF
C16813 VDD a_34226_24552# 0.59fF
C16814 _1192_.A2 nmat.col_n[31] 1.71fF
C16815 a_6830_22895# a_12175_27221# 0.43fF
C16816 nmat.rowoff_n[1] vcm 0.30fF
C16817 a_28202_59142# vcm 0.62fF
C16818 a_50290_22544# m2_51064_22274# 0.96fF
C16819 a_30210_12504# a_30210_11500# 1.00fF
C16820 a_12345_39100# cgen.dlycontrol2_in[1] 2.94fF
C16821 pmat.row_n[2] a_12079_9615# 1.43fF
C16822 a_6829_26703# a_8568_26703# 1.81fF
C16823 a_23182_56130# ctopp 3.40fF
C16824 pmat.rowoff_n[7] a_3045_19093# 0.60fF
C16825 a_12341_57141# a_12613_57141# 0.50fF
C16826 a_1923_61759# a_3175_59585# 0.34fF
C16827 VDD a_32218_56130# 0.55fF
C16828 a_39246_20536# a_40250_20536# 0.97fF
C16829 a_8491_47911# a_3746_58487# 0.35fF
C16830 a_24186_8488# m2_23956_7214# 1.00fF
C16831 a_10239_14183# a_1957_43567# 0.47fF
C16832 VDD m2_17246_6268# 0.59fF
C16833 VDD a_19166_17524# 0.56fF
C16834 a_18546_62196# a_46182_62154# 0.35fF
C16835 a_18546_66212# a_42166_66170# 0.35fF
C16836 a_38242_9492# a_38242_8488# 1.00fF
C16837 a_26194_66170# ctopp 3.58fF
C16838 VDD a_5253_32687# 0.59fF
C16839 VDD a_35230_66170# 0.52fF
C16840 VDD a_20170_8488# 0.56fF
C16841 VDD a_27605_37127# 1.06fF
C16842 VDD a_11019_71543# 1.38fF
C16843 nmat.col_n[23] vcm 2.80fF
C16844 VDD a_28202_63158# 0.52fF
C16845 pmat.en_bit_n[0] a_23021_29199# 0.92fF
C16846 a_2564_21959# a_4308_21495# 0.30fF
C16847 a_11927_27399# a_10223_26703# 1.00fF
C16848 pmat.row_n[11] pmat.rowoff_n[8] 1.40fF
C16849 a_49286_57134# a_50290_57134# 0.97fF
C16850 a_18546_61192# a_27106_61150# 0.35fF
C16851 a_21739_29415# a_15667_27239# 0.48fF
C16852 nmat.en_bit_n[0] nmat.col[17] 0.32fF
C16853 a_21174_71190# a_21174_70186# 1.00fF
C16854 a_48282_71190# a_49286_71190# 0.97fF
C16855 nmat.col[24] nmat.col[19] 12.89fF
C16856 a_10883_3303# a_7026_24527# 1.74fF
C16857 ANTENNA__1196__A2.DIODE a_7415_29397# 0.31fF
C16858 a_35230_58138# a_36234_58138# 0.97fF
C16859 a_10055_31591# pmat.row_n[4] 3.04fF
C16860 a_33423_47695# a_6664_26159# 0.66fF
C16861 VDD a_1895_43194# 0.55fF
C16862 a_2835_13077# comp_latch 0.55fF
C16863 VDD m2_51064_22274# 1.00fF
C16864 VDD a_40645_46519# 0.32fF
C16865 VDD a_18547_51565# 3.89fF
C16866 a_28202_19532# vcm 0.65fF
C16867 VDD a_12851_28853# 2.22fF
C16868 VDD a_4503_6335# 0.40fF
C16869 a_27198_10496# vcm 0.65fF
C16870 VDD a_7847_73493# 0.58fF
C16871 a_7693_22365# a_3305_15823# 1.13fF
C16872 a_10873_39605# cgen.dlycontrol4_in[2] 0.96fF
C16873 a_14691_27399# nmat.col_n[1] 0.38fF
C16874 a_2935_38279# a_3325_40847# 0.34fF
C16875 a_35230_61150# a_35230_60146# 1.00fF
C16876 a_24186_67174# ctopp 3.58fF
C16877 VDD a_14833_23089# 0.38fF
C16878 VDD a_22541_38779# 1.30fF
C16879 nmat.col[30] nmat.col_n[30] 1.33fF
C16880 cgen.enable_dlycontrol_in a_20221_40835# 3.21fF
C16881 a_43262_19532# a_43262_18528# 1.00fF
C16882 a_18546_70228# a_44174_70186# 0.35fF
C16883 VDD a_33222_67174# 0.52fF
C16884 pmat.row_n[5] ctopn 1.65fF
C16885 VDD a_23847_38007# 0.64fF
C16886 VDD a_34611_42089# 0.64fF
C16887 VDD a_22178_14512# 0.52fF
C16888 a_43262_62154# vcm 0.62fF
C16889 VDD a_21174_64162# 0.52fF
C16890 a_7840_27247# a_2683_22089# 0.59fF
C16891 VDD a_3199_40455# 0.51fF
C16892 a_18546_17522# a_39154_17930# 0.35fF
C16893 a_18546_57176# a_35138_57134# 0.35fF
C16894 cgen.dlycontrol4_in[1] a_2411_16101# 0.47fF
C16895 a_36234_59142# a_36234_58138# 1.00fF
C16896 a_4128_46983# a_5173_45993# 0.34fF
C16897 a_11067_30287# a_26155_46831# 0.63fF
C16898 a_43262_8488# m2_43032_7214# 1.00fF
C16899 pmat.col_n[3] pmat.col[3] 0.76fF
C16900 pmat.col_n[29] pmat.col[30] 5.95fF
C16901 a_18546_15514# a_39154_15922# 0.35fF
C16902 a_28202_15516# a_29206_15516# 0.97fF
C16903 a_10239_14183# cgen.enable_dlycontrol_in 0.86fF
C16904 a_1923_31743# a_1591_23445# 0.33fF
C16905 pmat.rowoff_n[5] ctopp 0.60fF
C16906 VDD a_11948_49783# 10.74fF
C16907 VDD a_29163_29423# 1.05fF
C16908 a_27198_69182# a_28202_69182# 0.97fF
C16909 VDD a_18546_59184# 32.64fF
C16910 VDD a_2046_30184# 10.95fF
C16911 a_42258_70186# vcm 0.62fF
C16912 a_29206_11500# vcm 0.65fF
C16913 VDD a_10383_13077# 0.55fF
C16914 a_1769_13103# config_2_in[11] 0.67fF
C16915 _1192_.B1 nmat.col_n[14] 0.46fF
C16916 VDD a_30571_50959# 11.34fF
C16917 VDD a_9301_62613# 0.65fF
C16918 a_35230_24552# a_35230_23548# 1.00fF
C16919 a_31263_28309# a_30699_29397# 0.48fF
C16920 nmat.col[29] vcm 6.39fF
C16921 VDD a_12171_18005# 0.44fF
C16922 a_41254_17524# a_41254_16520# 1.00fF
C16923 a_41731_49525# a_46753_41935# 0.59fF
C16924 a_47278_12504# a_48282_12504# 0.97fF
C16925 nmat.col_n[14] m2_32992_24282# 0.37fF
C16926 nmat.col[19] m2_38012_24282# 0.39fF
C16927 a_4128_64391# a_5179_31591# 0.74fF
C16928 a_31214_19532# ctopn 3.58fF
C16929 a_20572_40517# a_10767_39087# 0.93fF
C16930 VDD a_24186_65166# 0.52fF
C16931 VDD a_1586_18231# 13.87fF
C16932 VDD a_31214_21540# 0.52fF
C16933 _1194_.A2 ANTENNA__1197__B.DIODE 0.55fF
C16934 a_36234_59142# a_37238_59142# 0.97fF
C16935 m2_17932_69002# vcm 0.44fF
C16936 a_13091_28327# a_17139_30503# 1.12fF
C16937 a_30210_10496# ctopn 3.58fF
C16938 a_18546_68220# a_26102_68178# 0.35fF
C16939 a_50290_71190# ctopp 3.24fF
C16940 VDD a_11444_55535# 0.42fF
C16941 a_2683_22089# a_4523_21276# 0.54fF
C16942 a_37238_58138# ctopp 3.58fF
C16943 a_33222_68178# vcm 0.62fF
C16944 VDD a_46274_58138# 0.52fF
C16945 VDD ANTENNA__1190__A2.DIODE 11.84fF
C16946 a_25190_23548# a_25190_22544# 1.00fF
C16947 a_22085_42902# a_15049_42902# 0.36fF
C16948 pmat.rowoff_n[12] nmat.rowon_n[2] 0.39fF
C16949 a_24186_60146# a_25190_60146# 0.97fF
C16950 a_18546_60188# a_31122_60146# 0.35fF
C16951 pmat.row_n[9] pmat.row_n[8] 1.42fF
C16952 a_2021_9563# a_2972_9991# 0.83fF
C16953 a_24747_29967# nmat.col_n[31] 1.95fF
C16954 VDD a_44811_36469# 1.04fF
C16955 pmat.row_n[11] a_10239_14183# 3.60fF
C16956 m2_17932_8218# vcm 0.42fF
C16957 VDD a_18546_19530# 32.63fF
C16958 a_8491_47911# pmat.rowon_n[7] 0.72fF
C16959 a_12447_16143# pmat.row_n[0] 0.31fF
C16960 a_32218_68178# a_32218_67174# 1.00fF
C16961 a_10515_61839# nmat.rowon_n[13] 0.35fF
C16962 a_38242_23548# vcm 0.65fF
C16963 a_29206_69182# ctopp 3.58fF
C16964 a_40250_9492# vcm 0.65fF
C16965 VDD a_38242_69182# 0.52fF
C16966 m2_18936_72014# m2_19940_72014# 0.96fF
C16967 VDD a_46947_39215# 0.84fF
C16968 cgen.enable_dlycontrol_in cgen.dlycontrol1_in[0] 1.05fF
C16969 VDD m2_17932_23278# 1.02fF
C16970 a_2007_25597# a_9963_28111# 1.07fF
C16971 a_38242_59142# ctopp 3.58fF
C16972 a_20438_35431# a_12228_39605# 0.34fF
C16973 a_4075_31591# a_14379_6567# 0.50fF
C16974 a_32218_11500# ctopn 3.58fF
C16975 VDD a_47278_59142# 0.52fF
C16976 VDD a_11409_34789# 1.26fF
C16977 a_30210_16520# a_31214_16520# 0.97fF
C16978 a_18546_16518# a_43170_16926# 0.35fF
C16979 a_20170_67174# a_20170_66170# 1.00fF
C16980 VDD a_11883_62063# 1.22fF
C16981 VDD a_24186_61150# 0.52fF
C16982 a_11067_16359# a_4259_31375# 0.38fF
C16983 a_36234_13508# vcm 0.65fF
C16984 _1179_.X ANTENNA__1197__A.DIODE 2.77fF
C16985 VDD a_1823_64213# 1.11fF
C16986 a_2315_44124# a_4128_46983# 0.43fF
C16987 a_34226_18528# vcm 0.65fF
C16988 a_18546_17522# a_21082_17930# 0.35fF
C16989 pmat.sample_n a_11948_49783# 0.61fF
C16990 _1196_.B1 ANTENNA__1183__B1.DIODE 0.74fF
C16991 a_22178_20536# a_22178_19532# 1.00fF
C16992 a_19166_15516# ctopn 3.43fF
C16993 pmat.col_n[13] clk_ena 0.51fF
C16994 VDD a_19166_11500# 0.58fF
C16995 VDD a_3325_26159# 1.05fF
C16996 nmat.col[12] ctopn 1.97fF
C16997 a_45270_15516# vcm 0.65fF
C16998 VDD a_30210_17524# 0.52fF
C16999 a_18546_15514# a_21082_15922# 0.35fF
C17000 _1187_.A2 _1194_.B1 0.45fF
C17001 a_18546_8486# a_23090_8894# 0.35fF
C17002 pmat.row_n[13] ctopn 1.65fF
C17003 a_18546_69224# a_19074_69182# 0.35fF
C17004 pmat.rowon_n[13] a_18162_69222# 1.19fF
C17005 a_39246_70186# a_39246_69182# 1.00fF
C17006 VDD a_31214_8488# 0.55fF
C17007 a_14773_37218# a_10873_36341# 0.50fF
C17008 a_11149_36924# a_28431_34735# 0.33fF
C17009 cgen.dlycontrol3_in[1] a_14589_40726# 3.03fF
C17010 a_18546_21538# a_34134_21946# 0.35fF
C17011 VDD a_13719_36649# 0.57fF
C17012 m2_17932_64986# m2_17932_63982# 0.99fF
C17013 a_35312_31599# a_38913_31055# 0.38fF
C17014 a_28202_14512# a_28202_13508# 1.00fF
C17015 a_41254_23548# ctopn 3.40fF
C17016 a_2659_35015# a_3325_43023# 0.34fF
C17017 VDD a_47278_19532# 0.52fF
C17018 a_43262_9492# ctopn 3.57fF
C17019 m2_28976_24282# m3_29108_24414# 2.79fF
C17020 VDD m2_51064_71010# 1.05fF
C17021 a_32218_57134# a_32218_56130# 1.00fF
C17022 nmat.col_n[28] m2_47048_24282# 0.47fF
C17023 VDD nmat.col_n[1] 13.02fF
C17024 a_36234_19532# a_37238_19532# 0.97fF
C17025 a_41254_60146# vcm 0.62fF
C17026 pmat.col_n[7] pmat.col[8] 5.97fF
C17027 VDD a_46274_10496# 0.52fF
C17028 a_6467_29415# a_3688_17179# 0.56fF
C17029 VDD a_22361_41479# 1.82fF
C17030 VDD a_9485_15279# 0.35fF
C17031 VDD a_4259_65103# 0.74fF
C17032 VDD a_15667_28111# 4.10fF
C17033 pmat.row_n[7] a_18162_63198# 25.57fF
C17034 a_13091_28327# _1184_.A2 0.95fF
C17035 a_1858_25615# a_19439_32149# 0.96fF
C17036 a_35230_10496# a_36234_10496# 0.97fF
C17037 pmat.rowoff_n[12] cgen.dlycontrol4_in[2] 0.41fF
C17038 VDD a_26194_12504# 0.52fF
C17039 VDD m2_51064_10226# 1.03fF
C17040 a_47278_16520# vcm 0.65fF
C17041 a_10883_3303# nmat.col_n[10] 1.66fF
C17042 VDD a_1769_14735# 6.34fF
C17043 a_45019_38645# nmat.col[28] 0.39fF
C17044 a_20170_9492# a_20170_8488# 1.00fF
C17045 a_46274_56130# a_47278_56130# 0.97fF
C17046 a_39246_13508# ctopn 3.58fF
C17047 _1192_.B1 a_13459_28111# 0.88fF
C17048 VDD a_5351_60663# 0.53fF
C17049 a_10883_3303# clk_ena 0.30fF
C17050 a_34226_57134# vcm 0.62fF
C17051 VDD cgen.dlycontrol2_in[0] 5.22fF
C17052 a_33222_71190# vcm 0.60fF
C17053 a_37238_18528# ctopn 3.58fF
C17054 a_20170_58138# vcm 0.62fF
C17055 nmat.sw comp_latch 0.39fF
C17056 m2_21948_7214# m3_22080_7346# 2.79fF
C17057 pmat.en_bit_n[2] nmat.en_bit_n[0] 1.05fF
C17058 nmat.col_n[18] nmat.col_n[19] 0.95fF
C17059 VDD a_14533_39631# 1.75fF
C17060 pmat.row_n[11] ctopn 1.65fF
C17061 a_20170_23548# vcm 0.65fF
C17062 a_13091_28327# pmat.col[22] 0.35fF
C17063 a_32687_46607# a_31675_47695# 0.31fF
C17064 a_48282_15516# ctopn 3.58fF
C17065 VDD a_48282_11500# 0.52fF
C17066 a_18243_28327# a_8583_29199# 0.40fF
C17067 ANTENNA__1190__B1.DIODE ANTENNA__1195__A1.DIODE 0.34fF
C17068 a_11067_27239# a_21739_29415# 2.00fF
C17069 a_12069_38517# a_12197_38306# 1.28fF
C17070 a_28202_22544# a_29206_22544# 0.97fF
C17071 VDD a_11133_44581# 1.14fF
C17072 a_7847_73493# a_8013_73493# 0.69fF
C17073 a_12069_38517# a_12116_39783# 1.73fF
C17074 a_49286_66170# a_50290_66170# 0.97fF
C17075 a_17139_30503# a_26891_28327# 2.97fF
C17076 VDD dummypin[10] 0.90fF
C17077 a_43533_30761# a_28704_29568# 0.32fF
C17078 pmat.col[6] ctopp 1.97fF
C17079 pmat.col[1] vcm 5.88fF
C17080 a_18546_69224# a_48190_69182# 0.35fF
C17081 pmat.row_n[13] pmat.row_n[10] 7.48fF
C17082 VDD a_6337_6825# 0.33fF
C17083 nmat.col_n[5] m2_23956_24282# 0.37fF
C17084 a_13091_28327# a_9411_2215# 2.01fF
C17085 a_19166_21540# a_19166_20536# 1.00fF
C17086 a_2411_33749# cgen.dlycontrol1_in[0] 0.45fF
C17087 cgen.dlycontrol3_in[4] a_22537_36911# 2.39fF
C17088 _1154_.X _1187_.A2 0.61fF
C17089 nmat.rowon_n[1] ctopn 1.39fF
C17090 a_42258_63158# a_43262_63158# 0.97fF
C17091 a_18546_9490# a_22086_9898# 0.35fF
C17092 a_11797_60431# a_12237_60431# 0.36fF
C17093 a_45270_22544# vcm 0.65fF
C17094 a_2263_43719# a_10515_13967# 0.60fF
C17095 a_43262_68178# ctopp 3.58fF
C17096 nmat.sw cgen.dlycontrol4_in[2] 2.49fF
C17097 VDD a_1643_67477# 0.35fF
C17098 a_21174_59142# vcm 0.62fF
C17099 a_7109_29423# a_9963_28111# 3.74fF
C17100 pmat.col_n[16] a_35230_55126# 0.31fF
C17101 a_14825_50095# a_11711_50959# 0.34fF
C17102 a_6883_51335# a_6979_51157# 0.37fF
C17103 VDD a_25190_56130# 0.55fF
C17104 a_10873_36341# clk_ena 2.83fF
C17105 a_19541_28879# a_15899_47939# 0.60fF
C17106 a_50290_16520# ctopn 3.43fF
C17107 a_19166_8488# m2_18936_7214# 1.00fF
C17108 a_10239_14183# pmat.row_n[2] 0.47fF
C17109 VDD a_5746_11703# 0.98fF
C17110 pmat.col[4] vcm 5.88fF
C17111 VDD m2_38012_7214# 0.93fF
C17112 pmat.rowon_n[3] a_1739_47893# 0.31fF
C17113 VDD a_2467_16341# 0.86fF
C17114 VDD a_12559_51325# 0.51fF
C17115 VDD a_3267_74817# 0.54fF
C17116 a_18546_62196# a_39154_62154# 0.35fF
C17117 a_1586_8439# a_2199_13887# 0.79fF
C17118 VDD a_35786_47893# 1.03fF
C17119 a_18546_66212# a_35138_66170# 0.35fF
C17120 VDD a_28202_66170# 0.52fF
C17121 a_34924_37253# a_11297_36091# 0.49fF
C17122 a_37238_11500# a_38242_11500# 0.97fF
C17123 a_15101_29423# nmat.col[12] 0.71fF
C17124 nmat.col_n[11] vcm 2.80fF
C17125 VDD a_21174_63158# 0.52fF
C17126 pmat.sample a_20848_41605# 0.49fF
C17127 a_39246_64162# a_39246_63158# 1.00fF
C17128 m2_39016_54946# m3_39148_55078# 2.79fF
C17129 a_5651_66975# a_5267_65479# 0.38fF
C17130 pmat.row_n[11] pmat.row_n[10] 0.49fF
C17131 a_42258_10496# a_42258_9492# 1.00fF
C17132 a_39246_58138# a_39246_57134# 1.00fF
C17133 pmat.en_bit_n[0] ANTENNA__1395__B1.DIODE 2.25fF
C17134 a_4025_54965# a_4587_53505# 0.34fF
C17135 VDD a_26276_39429# 1.05fF
C17136 VDD a_26552_43781# 0.96fF
C17137 _1224_.X nmat.col_n[30] 0.90fF
C17138 a_10239_14183# nmat.col_n[13] 0.49fF
C17139 a_21174_19532# vcm 0.65fF
C17140 a_18546_59184# a_19074_59142# 0.35fF
C17141 a_43262_60146# a_43262_59142# 1.00fF
C17142 a_31214_18528# a_31214_17524# 1.00fF
C17143 a_32218_63158# pmat.col[13] 0.31fF
C17144 a_12513_36924# nmat.sample 0.38fF
C17145 m3_50192_24414# ctopn 0.35fF
C17146 VDD cgen.dlycontrol1_in[2] 5.23fF
C17147 a_24867_53135# a_15667_27239# 0.54fF
C17148 VDD a_10845_12559# 0.39fF
C17149 pmat.col_n[18] pmat.col[19] 6.74fF
C17150 a_48282_22544# ctopn 3.57fF
C17151 a_11041_39860# cgen.dlycontrol4_in[0] 0.32fF
C17152 VDD dummypin[11] 0.87fF
C17153 a_16083_50069# a_19283_49783# 0.43fF
C17154 pmat.row_n[10] nmat.rowon_n[1] 0.34fF
C17155 a_31214_63158# a_31214_62154# 1.00fF
C17156 VDD a_17191_48981# 0.31fF
C17157 a_47278_67174# a_48282_67174# 0.97fF
C17158 VDD cgen.dlycontrol2_in[1] 6.00fF
C17159 a_14287_69455# pmat.rowon_n[0] 0.88fF
C17160 a_12171_18005# a_12337_18005# 0.63fF
C17161 a_18546_70228# a_37146_70186# 0.35fF
C17162 VDD a_26194_67174# 0.52fF
C17163 VDD a_6559_8527# 0.44fF
C17164 a_9335_51727# a_9463_50877# 0.32fF
C17165 a_9675_10396# a_11501_10927# 0.44fF
C17166 a_44266_66170# a_44266_65166# 1.00fF
C17167 a_37238_22544# a_37238_21540# 1.00fF
C17168 VDD a_20645_42044# 1.38fF
C17169 a_2411_43301# a_4955_40277# 0.50fF
C17170 a_36234_14512# a_37238_14512# 0.97fF
C17171 a_36234_62154# vcm 0.62fF
C17172 a_15435_29111# nmat.col[10] 0.37fF
C17173 a_8583_29199# a_12851_28853# 0.46fF
C17174 a_18546_17522# a_32126_17930# 0.35fF
C17175 a_35230_64162# a_36234_64162# 0.97fF
C17176 a_11067_16359# a_6173_22895# 0.71fF
C17177 a_1858_25615# a_15660_31029# 0.37fF
C17178 a_41254_68178# a_42258_68178# 0.97fF
C17179 a_18546_57176# a_28110_57134# 0.35fF
C17180 a_14773_39394# cgen.dlycontrol2_in[1] 4.02fF
C17181 VDD _1194_.A2 33.01fF
C17182 a_33423_47695# a_45112_47607# 1.27fF
C17183 a_11067_30287# nmat.rowon_n[12] 0.32fF
C17184 a_30210_13508# a_30210_12504# 1.00fF
C17185 a_8695_12801# a_8656_12675# 0.75fF
C17186 a_18546_72236# a_44174_72194# 0.35fF
C17187 VDD a_46968_45743# 0.38fF
C17188 a_31095_42367# a_10781_42364# 0.76fF
C17189 a_18546_15514# a_32126_15922# 0.35fF
C17190 a_40837_46261# a_45325_38127# 0.72fF
C17191 config_1_in[6] VSS 1.17fF
C17192 config_1_in[7] VSS 1.21fF
C17193 config_1_in[8] VSS 1.11fF
C17194 config_1_in[9] VSS 1.17fF
C17195 config_1_in[0] VSS 1.08fF
C17196 config_1_in[1] VSS 1.04fF
C17197 config_1_in[2] VSS 1.27fF
C17198 config_1_in[3] VSS 1.38fF
C17199 config_1_in[4] VSS 0.85fF
C17200 config_1_in[5] VSS 1.07fF
C17201 config_1_in[10] VSS 1.11fF
C17202 config_1_in[11] VSS 0.88fF
C17203 config_1_in[12] VSS 1.06fF
C17204 config_1_in[13] VSS 1.67fF
C17205 config_1_in[14] VSS 0.87fF
C17206 config_1_in[15] VSS 1.49fF
C17207 rst_n VSS 1.33fF
C17208 start_conversion_in VSS 0.94fF
C17209 config_2_in[0] VSS 0.96fF
C17210 config_2_in[1] VSS 1.00fF
C17211 config_2_in[2] VSS 1.03fF
C17212 config_2_in[3] VSS 0.87fF
C17213 clk_dig VSS 4.34fF
C17214 config_2_in[4] VSS 1.02fF
C17215 config_2_in[5] VSS 1.04fF
C17216 config_2_in[6] VSS 0.91fF
C17217 ndecision_finish VSS 6.09fF
C17218 clk_comp VSS 3.51fF
C17219 comp_latch VSS 24.38fF
C17220 ctopn VSS -372.32fF
C17221 config_2_in[7] VSS 1.02fF
C17222 config_2_in[8] VSS 0.99fF
C17223 config_2_in[9] VSS 0.92fF
C17224 config_2_in[10] VSS 1.12fF
C17225 config_2_in[12] VSS 1.19fF
C17226 config_2_in[11] VSS 1.31fF
C17227 config_2_in[13] VSS 0.85fF
C17228 config_2_in[14] VSS 1.18fF
C17229 config_2_in[15] VSS 1.32fF
C17230 result_out[0] VSS 0.60fF
C17231 result_out[1] VSS 0.69fF
C17232 ctopp VSS -372.75fF
C17233 clk_ena VSS 39.10fF
C17234 result_out[2] VSS 0.83fF
C17235 result_out[3] VSS 0.58fF
C17236 result_out[4] VSS 0.84fF
C17237 result_out[5] VSS 0.85fF
C17238 result_out[6] VSS 0.61fF
C17239 result_out[7] VSS 0.88fF
C17240 result_out[8] VSS 0.76fF
C17241 result_out[9] VSS 0.66fF
C17242 result_out[10] VSS 0.78fF
C17243 result_out[11] VSS 0.77fF
C17244 result_out[12] VSS 0.77fF
C17245 result_out[13] VSS 0.79fF
C17246 vcm VSS 23346.50fF
C17247 result_out[14] VSS 0.72fF
C17248 result_out[15] VSS 0.88fF
C17249 conversion_finished_out VSS 0.75fF
C17550 dummypin[15] VSS 0.95fF
C17551 adc_top_96.HI VSS 0.32fF
C17552 a_82735_2223# VSS 0.38fF
C17553 a_84090_3087# VSS 0.39fF
C17554 a_83630_3311# VSS 0.38fF
C17555 a_83238_4175# VSS 0.49fF
C17556 a_82778_4399# VSS 0.49fF
C17557 a_83170_5263# VSS 0.39fF
C17558 a_2219_4943# VSS 0.43fF
C17559 a_1775_5059# VSS 0.30fF
C17560 a_1761_2767# VSS 0.65fF
C17561 a_6487_5629# VSS 0.55fF
C17562 a_5967_5461# VSS 0.37fF
C17563 dummypin[14] VSS 0.84fF
C17564 adc_top_95.HI VSS 0.34fF
C17565 a_84028_9615# VSS 0.32fF
C17566 a_9655_6335# VSS 0.40fF
C17567 a_8703_6202# VSS 0.34fF
C17568 a_8399_6037# VSS 0.49fF
C17569 a_6559_6031# VSS 0.32fF
C17570 a_4503_6335# VSS 0.41fF
C17571 a_3247_6037# VSS 0.48fF
C17572 a_1761_6031# VSS 0.35fF
C17573 a_51202_7890# VSS 0.49fF
C17574 a_50198_7890# VSS 0.40fF
C17575 a_49194_7890# VSS 0.39fF
C17576 a_48190_7890# VSS 0.38fF
C17577 a_47186_7890# VSS 0.38fF
C17578 a_46182_7890# VSS 0.39fF
C17579 a_45178_7890# VSS 0.39fF
C17580 a_44174_7890# VSS 0.38fF
C17581 a_43170_7890# VSS 0.38fF
C17582 a_42166_7890# VSS 0.39fF
C17583 a_41162_7890# VSS 0.39fF
C17584 a_40158_7890# VSS 0.38fF
C17585 a_39154_7890# VSS 0.38fF
C17586 a_38150_7890# VSS 0.39fF
C17587 a_37146_7890# VSS 0.40fF
C17588 a_36142_7890# VSS 0.38fF
C17589 a_35138_7890# VSS 0.38fF
C17590 a_34134_7890# VSS 0.39fF
C17591 a_33130_7890# VSS 0.40fF
C17592 a_32126_7890# VSS 0.38fF
C17593 a_31122_7890# VSS 0.38fF
C17594 a_30118_7890# VSS 0.39fF
C17595 a_29114_7890# VSS 0.40fF
C17596 a_28110_7890# VSS 0.38fF
C17597 a_27106_7890# VSS 0.38fF
C17598 a_26102_7890# VSS 0.40fF
C17599 a_25098_7890# VSS 0.39fF
C17600 a_24094_7890# VSS 0.38fF
C17601 a_23090_7890# VSS 0.38fF
C17602 a_22086_7890# VSS 0.40fF
C17603 a_21082_7890# VSS 0.40fF
C17604 a_9459_5461# VSS 0.69fF
C17605 a_6337_6825# VSS 0.39fF
C17606 nmat.rowoff_n[1] VSS 1.83fF
C17607 a_20078_7890# VSS 0.38fF
C17608 a_19074_7890# VSS 0.39fF
C17609 a_18162_7484# VSS 5.71fF
C17610 a_18546_7482# VSS 8.97fF
C17611 a_9195_7423# VSS 0.41fF
C17612 a_8105_7125# VSS 0.33fF
C17613 a_7939_7125# VSS 0.54fF
C17614 a_3551_6202# VSS 0.96fF
C17615 a_1761_7119# VSS 0.58fF
C17616 a_18162_8488# VSS 4.97fF
C17617 a_18546_8486# VSS 3.53fF
C17618 a_4254_7351# VSS 0.60fF
C17619 a_8243_7290# VSS 0.58fF
C17620 a_14071_8511# VSS 0.42fF
C17621 a_12257_8527# VSS 0.39fF
C17622 a_12815_8213# VSS 0.47fF
C17623 a_2847_8511# VSS 0.53fF
C17624 a_1591_8213# VSS 0.56fF
C17625 nmat.rowon_n[15] VSS 4.29fF
C17626 a_18162_9492# VSS 4.95fF
C17627 a_18546_9490# VSS 3.50fF
C17628 nmat.rowoff_n[3] VSS 1.82fF
C17629 a_12133_9001# VSS 0.43fF
C17630 a_10378_7637# VSS 1.10fF
C17631 a_10047_8751# VSS 0.57fF
C17632 a_1895_8378# VSS 0.53fF
C17633 a_6559_8527# VSS 0.96fF
C17634 a_7040_8725# VSS 0.36fF
C17635 a_6872_8725# VSS 0.49fF
C17636 a_6412_8725# VSS 0.36fF
C17637 nmat.rowoff_n[2] VSS 1.55fF
C17638 a_5654_9527# VSS 1.41fF
C17639 a_5558_9527# VSS 0.93fF
C17640 a_4865_8181# VSS 0.97fF
C17641 a_5325_9269# VSS 0.31fF
C17642 dummypin[13] VSS 0.83fF
C17643 adc_top_94.HI VSS 0.31fF
C17644 a_82971_11989# VSS 0.33fF
C17645 a_82787_13077# VSS 0.31fF
C17646 a_18162_10496# VSS 4.95fF
C17647 a_18546_10494# VSS 3.50fF
C17648 a_9583_10121# VSS 2.94fF
C17649 a_4611_9839# VSS 0.79fF
C17650 a_3415_9839# VSS 0.43fF
C17651 a_3663_9269# VSS 1.18fF
C17652 a_4338_9839# VSS 0.30fF
C17653 a_3609_9295# VSS 0.80fF
C17654 a_4167_9615# VSS 0.52fF
C17655 a_2972_9991# VSS 1.84fF
C17656 a_11051_8903# VSS 0.44fF
C17657 a_13795_10687# VSS 0.40fF
C17658 a_11987_10089# VSS 0.35fF
C17659 a_12539_10389# VSS 0.56fF
C17660 a_9668_10651# VSS 1.74fF
C17661 a_8481_10396# VSS 1.06fF
C17662 a_6607_10615# VSS 0.33fF
C17663 a_18162_11500# VSS 4.95fF
C17664 a_18546_11498# VSS 3.50fF
C17665 a_11501_10927# VSS 0.33fF
C17666 a_8111_11209# VSS 0.45fF
C17667 a_1959_10615# VSS 0.38fF
C17668 a_1761_9839# VSS 0.39fF
C17669 a_11167_11177# VSS 0.33fF
C17670 a_9675_10396# VSS 0.95fF
C17671 a_11207_11079# VSS 0.34fF
C17672 a_5012_10927# VSS 0.87fF
C17673 a_4989_11079# VSS 0.58fF
C17674 nmat.rowoff_n[5] VSS 1.68fF
C17675 a_5223_11079# VSS 0.31fF
C17676 a_8693_11769# VSS 0.30fF
C17677 a_8479_11484# VSS 0.60fF
C17678 a_8472_11739# VSS 0.36fF
C17679 a_2021_11043# VSS 2.87fF
C17680 a_7283_11484# VSS 0.77fF
C17681 a_2021_9563# VSS 3.20fF
C17682 a_5768_9527# VSS 0.57fF
C17683 a_5746_11703# VSS 0.37fF
C17684 a_3583_11775# VSS 0.55fF
C17685 a_2129_10383# VSS 0.68fF
C17686 a_2327_11477# VSS 0.40fF
C17687 a_18162_12504# VSS 4.95fF
C17688 a_18546_12502# VSS 3.51fF
C17689 a_5363_12015# VSS 0.55fF
C17690 a_1761_11471# VSS 0.60fF
C17691 a_10839_11989# VSS 1.34fF
C17692 a_12967_12863# VSS 0.41fF
C17693 a_10845_12559# VSS 0.70fF
C17694 a_11711_12565# VSS 0.54fF
C17695 a_10471_12791# VSS 0.37fF
C17696 a_8695_12801# VSS 0.60fF
C17697 a_8175_12533# VSS 0.42fF
C17698 a_18162_13508# VSS 4.96fF
C17699 a_18546_13506# VSS 3.50fF
C17700 nmat.rowoff_n[8] VSS 1.17fF
C17701 a_8031_13353# VSS 1.38fF
C17702 a_4895_12559# VSS 0.79fF
C17703 a_10383_13077# VSS 0.58fF
C17704 a_5579_12394# VSS 2.34fF
C17705 a_5173_9839# VSS 1.31fF
C17706 a_5227_13077# VSS 0.31fF
C17707 a_2499_13077# VSS 0.42fF
C17708 dummypin[12] VSS 0.68fF
C17709 adc_top_93.HI VSS 0.34fF
C17710 a_82787_14709# VSS 0.31fF
C17711 a_18162_14512# VSS 4.95fF
C17712 a_18546_14510# VSS 3.50fF
C17713 a_13686_13967# VSS 0.49fF
C17714 nmat.rowoff_n[9] VSS 1.25fF
C17715 a_4865_12533# VSS 0.81fF
C17716 a_1717_13647# VSS 5.39fF
C17717 a_5331_13951# VSS 0.37fF
C17718 a_4075_13653# VSS 0.56fF
C17719 a_2129_12559# VSS 0.42fF
C17720 a_2439_13889# VSS 0.41fF
C17721 a_2199_13887# VSS 9.32fF
C17722 a_1687_13621# VSS 0.60fF
C17723 nmat.rowon_n[10] VSS 4.00fF
C17724 nmat.rowon_n[9] VSS 4.03fF
C17725 a_13446_14191# VSS 0.30fF
C17726 a_12047_14165# VSS 0.66fF
C17727 a_10791_14191# VSS 0.41fF
C17728 a_7419_14379# VSS 0.52fF
C17729 a_18162_15516# VSS 4.95fF
C17730 a_18546_15514# VSS 3.50fF
C17731 nmat.rowoff_n[10] VSS 1.02fF
C17732 a_7085_15055# VSS 0.62fF
C17733 a_7295_14441# VSS 0.39fF
C17734 a_6853_14967# VSS 0.58fF
C17735 a_5547_14735# VSS 0.46fF
C17736 a_4319_15039# VSS 0.48fF
C17737 a_3063_14741# VSS 0.59fF
C17738 nmat.rowoff_n[11] VSS 1.25fF
C17739 a_10575_15253# VSS 0.48fF
C17740 a_9319_15279# VSS 0.40fF
C17741 a_7631_15253# VSS 0.70fF
C17742 a_6375_15279# VSS 0.39fF
C17743 a_18162_16520# VSS 4.95fF
C17744 a_18546_16518# VSS 3.50fF
C17745 a_14457_15823# VSS 0.62fF
C17746 a_8937_15823# VSS 0.36fF
C17747 a_3367_14906# VSS 0.41fF
C17748 a_8767_16055# VSS 0.50fF
C17749 a_4215_15797# VSS 0.49fF
C17750 a_2847_16127# VSS 0.66fF
C17751 a_1591_15829# VSS 0.53fF
C17752 a_1586_8439# VSS 4.71fF
C17753 a_14195_7351# VSS 0.67fF
C17754 a_12875_16341# VSS 0.63fF
C17755 a_11619_16367# VSS 0.42fF
C17756 a_3571_13627# VSS 2.71fF
C17757 a_7387_16367# VSS 0.37fF
C17758 a_1895_15994# VSS 0.71fF
C17759 nmat.rowon_n[6] VSS 4.55fF
C17760 a_18162_17524# VSS 4.97fF
C17761 a_18546_17522# VSS 3.50fF
C17762 nmat.rowoff_n[13] VSS 1.15fF
C17763 a_6621_16885# VSS 0.38fF
C17764 a_5266_17143# VSS 1.05fF
C17765 a_2467_16341# VSS 0.50fF
C17766 a_3909_17209# VSS 0.32fF
C17767 a_11421_17455# VSS 0.55fF
C17768 a_14287_17455# VSS 0.48fF
C17769 a_5715_16911# VSS 0.41fF
C17770 a_4871_17429# VSS 0.56fF
C17771 dummypin[11] VSS 0.80fF
C17772 adc_top_92.HI VSS 0.34fF
C17773 a_18162_18528# VSS 4.95fF
C17774 a_18546_18526# VSS 3.50fF
C17775 a_13427_18303# VSS 0.70fF
C17776 a_11145_17999# VSS 0.79fF
C17777 a_12171_18005# VSS 0.52fF
C17778 a_9557_17705# VSS 0.30fF
C17779 a_8399_18115# VSS 0.34fF
C17780 a_7809_17705# VSS 0.37fF
C17781 a_6795_18319# VSS 0.50fF
C17782 a_3576_17143# VSS 3.14fF
C17783 a_2847_18303# VSS 0.69fF
C17784 a_1591_18005# VSS 0.52fF
C17785 nmat.rowon_n[13] VSS 4.53fF
C17786 a_4383_7093# VSS 10.45fF
C17787 a_10975_18231# VSS 0.39fF
C17788 a_6343_18517# VSS 0.42fF
C17789 a_5087_18543# VSS 0.40fF
C17790 a_1895_18170# VSS 0.68fF
C17791 a_2467_18517# VSS 0.68fF
C17792 nmat.rowon_n[4] VSS 4.27fF
C17793 a_18162_19532# VSS 4.95fF
C17794 a_18546_19530# VSS 3.50fF
C17795 a_14011_19087# VSS 0.41fF
C17796 a_9749_19061# VSS 0.39fF
C17797 a_5257_19087# VSS 0.32fF
C17798 a_4135_19391# VSS 0.43fF
C17799 a_2879_19093# VSS 0.57fF
C17800 a_5087_19319# VSS 0.30fF
C17801 a_7521_19631# VSS 0.65fF
C17802 a_18162_20536# VSS 4.95fF
C17803 a_18546_20534# VSS 3.50fF
C17804 a_10239_20291# VSS 0.30fF
C17805 a_3688_17179# VSS 2.50fF
C17806 a_4976_16091# VSS 3.75fF
C17807 a_9227_20291# VSS 0.38fF
C17808 a_6821_18543# VSS 0.65fF
C17809 a_5179_20175# VSS 0.41fF
C17810 a_4613_19087# VSS 0.99fF
C17811 a_2847_20479# VSS 0.41fF
C17812 a_1591_20181# VSS 0.53fF
C17813 nmat.rowon_n[2] VSS 5.25fF
C17814 a_18162_21540# VSS 4.96fF
C17815 a_18546_21538# VSS 3.50fF
C17816 nmat.rowoff_n[14] VSS 2.04fF
C17817 a_7847_20719# VSS 0.33fF
C17818 a_7644_16341# VSS 2.24fF
C17819 a_3183_19258# VSS 0.88fF
C17820 a_8305_20871# VSS 2.31fF
C17821 a_7533_19087# VSS 0.45fF
C17822 a_13467_21263# VSS 0.34fF
C17823 a_6981_21263# VSS 0.35fF
C17824 a_4123_20693# VSS 0.41fF
C17825 a_12155_20719# VSS 0.31fF
C17826 a_10498_19631# VSS 0.41fF
C17827 a_1895_20346# VSS 0.36fF
C17828 dummypin[10] VSS 0.87fF
C17829 adc_top_91.HI VSS 0.34fF
C17830 nmat.rowon_n[1] VSS 4.77fF
C17831 a_18162_22544# VSS 4.95fF
C17832 a_18546_22542# VSS 3.50fF
C17833 a_8507_20175# VSS 0.79fF
C17834 a_2099_21237# VSS 0.48fF
C17835 a_11897_21813# VSS 0.31fF
C17836 a_10932_21959# VSS 0.34fF
C17837 a_9135_22057# VSS 0.41fF
C17838 a_6469_21813# VSS 0.32fF
C17839 a_5455_22057# VSS 0.41fF
C17840 a_3305_15823# VSS 4.34fF
C17841 a_8197_20871# VSS 0.89fF
C17842 a_10071_17999# VSS 0.74fF
C17843 a_8859_22467# VSS 0.34fF
C17844 a_7479_22467# VSS 0.32fF
C17845 a_4811_22351# VSS 0.35fF
C17846 a_3859_22655# VSS 0.47fF
C17847 a_2603_22357# VSS 0.44fF
C17848 a_18162_23548# VSS 5.01fF
C17849 a_18546_23546# VSS 3.60fF
C17850 nmat.rowoff_n[0] VSS 1.32fF
C17851 a_11159_23145# VSS 1.95fF
C17852 a_7048_23277# VSS 0.97fF
C17853 a_3305_17999# VSS 2.11fF
C17854 a_2907_22522# VSS 0.59fF
C17855 a_12247_20175# VSS 0.88fF
C17856 a_5899_21807# VSS 3.04fF
C17857 a_7693_22365# VSS 2.24fF
C17858 a_10097_22895# VSS 0.67fF
C17859 a_9303_22351# VSS 0.53fF
C17860 a_6800_22869# VSS 0.36fF
C17861 a_5825_22901# VSS 0.32fF
C17862 a_4043_22869# VSS 0.58fF
C17863 a_8356_23671# VSS 0.31fF
C17864 a_6639_23413# VSS 0.41fF
C17865 a_5271_23447# VSS 0.31fF
C17866 a_2411_16101# VSS 8.27fF
C17867 a_2835_13077# VSS 10.93fF
C17868 a_3859_23699# VSS 0.53fF
C17869 a_2847_23743# VSS 0.38fF
C17870 a_1591_23445# VSS 0.48fF
C17871 a_51202_24958# VSS 0.36fF
C17872 a_36234_24552# VSS 0.53fF
C17873 a_35230_24552# VSS 0.39fF
C17874 a_34226_24552# VSS 0.39fF
C17875 a_20170_24552# VSS 0.40fF
C17876 a_10513_24135# VSS 0.55fF
C17877 a_3325_20175# VSS 4.56fF
C17878 a_3387_22869# VSS 0.53fF
C17879 a_14475_24233# VSS 0.32fF
C17880 a_13768_22325# VSS 0.63fF
C17881 a_13151_23957# VSS 0.46fF
C17882 a_12245_21807# VSS 0.37fF
C17883 a_7847_24233# VSS 0.30fF
C17884 a_5547_24233# VSS 0.38fF
C17885 a_18162_24552# VSS 6.82fF
C17886 a_18546_24550# VSS 4.46fF
C17887 a_13563_24527# VSS 0.31fF
C17888 a_12463_22351# VSS 1.04fF
C17889 a_11892_21959# VSS 0.73fF
C17890 a_10959_23983# VSS 0.46fF
C17891 a_11897_21263# VSS 0.44fF
C17892 a_8333_24847# VSS 0.75fF
C17893 a_8831_24501# VSS 1.49fF
C17894 a_6173_22895# VSS 1.01fF
C17895 a_8307_23439# VSS 0.42fF
C17896 a_4703_24527# VSS 0.79fF
C17897 a_6564_24527# VSS 0.54fF
C17898 a_4259_24643# VSS 0.31fF
C17899 a_4337_22351# VSS 1.11fF
C17900 a_3325_23439# VSS 0.85fF
C17901 a_3399_24787# VSS 0.48fF
C17902 a_1895_23610# VSS 0.32fF
C17903 nmat.col_n[1] VSS 9.82fF
C17904 a_14371_25071# VSS 0.84fF
C17905 a_9528_20407# VSS 4.59fF
C17906 a_2191_24501# VSS 0.60fF
C17907 a_9441_20189# VSS 2.61fF
C17908 nmat.col[3] VSS 9.78fF
C17909 a_4523_21276# VSS 3.84fF
C17910 a_7665_25731# VSS 0.32fF
C17911 a_6747_25731# VSS 0.31fF
C17912 a_3891_25623# VSS 0.30fF
C17913 a_2511_25615# VSS 0.42fF
C17914 dummypin[9] VSS 0.79fF
C17915 adc_top_90.HI VSS 0.35fF
C17916 nmat.col[1] VSS 9.31fF
C17917 a_6406_26159# VSS 0.37fF
C17918 a_9579_26159# VSS 0.55fF
C17919 a_2191_25045# VSS 0.47fF
C17920 a_3325_26159# VSS 0.70fF
C17921 a_8013_25615# VSS 3.61fF
C17922 a_9135_26409# VSS 0.32fF
C17923 a_7186_25615# VSS 0.52fF
C17924 a_7072_26311# VSS 0.53fF
C17925 a_2847_26133# VSS 0.36fF
C17926 a_1591_26159# VSS 0.50fF
C17927 a_8861_24527# VSS 0.50fF
C17928 a_12449_22895# VSS 0.58fF
C17929 a_13145_26935# VSS 0.45fF
C17930 a_9779_26819# VSS 0.40fF
C17931 a_9777_26935# VSS 1.01fF
C17932 a_8031_26703# VSS 0.47fF
C17933 a_7779_22583# VSS 1.48fF
C17934 a_5320_27023# VSS 0.95fF
C17935 a_4712_27023# VSS 0.49fF
C17936 a_2879_26703# VSS 0.43fF
C17937 nmat.col_n[24] VSS 23.91fF
C17938 nmat.col[26] VSS 19.69fF
C17939 nmat.col_n[27] VSS 8.69fF
C17940 nmat.col[27] VSS 6.33fF
C17941 nmat.col[25] VSS 6.18fF
C17942 nmat.col_n[23] VSS 8.71fF
C17943 nmat.col[22] VSS 6.31fF
C17944 nmat.col_n[17] VSS 8.11fF
C17945 nmat.col[17] VSS 6.06fF
C17946 nmat.col_n[29] VSS 20.12fF
C17947 nmat.col_n[19] VSS 20.63fF
C17948 nmat.col[16] VSS 6.42fF
C17949 a_16965_27247# VSS 1.26fF
C17950 nmat.col_n[11] VSS 8.47fF
C17951 nmat.col[11] VSS 6.49fF
C17952 nmat.col_n[8] VSS 8.82fF
C17953 nmat.col[8] VSS 6.20fF
C17954 nmat.col[6] VSS 6.39fF
C17955 nmat.col_n[5] VSS 8.59fF
C17956 nmat.col[5] VSS 6.25fF
C17957 nmat.col[2] VSS 6.34fF
C17958 a_9485_27247# VSS 0.51fF
C17959 a_37525_27221# VSS 0.33fF
C17960 a_8568_26703# VSS 0.81fF
C17961 a_6829_26703# VSS 1.90fF
C17962 a_14471_27247# VSS 0.49fF
C17963 a_11337_25071# VSS 1.50fF
C17964 a_11091_26311# VSS 0.61fF
C17965 a_6634_26133# VSS 0.80fF
C17966 a_4443_27247# VSS 0.42fF
C17967 nmat.col_n[25] VSS 8.64fF
C17968 nmat.col_n[22] VSS 8.59fF
C17969 nmat.col[23] VSS 6.25fF
C17970 nmat.col_n[26] VSS 19.58fF
C17971 nmat.col_n[20] VSS 8.47fF
C17972 nmat.col[20] VSS 6.25fF
C17973 nmat.col_n[16] VSS 8.11fF
C17974 nmat.col_n[15] VSS 8.08fF
C17975 nmat.col[14] VSS 7.39fF
C17976 nmat.col_n[14] VSS 8.35fF
C17977 nmat.col_n[9] VSS 8.55fF
C17978 nmat.col[19] VSS 18.09fF
C17979 nmat.col[9] VSS 6.41fF
C17980 nmat.col[18] VSS 24.61fF
C17981 nmat.col_n[0] VSS 8.84fF
C17982 nmat.col_n[6] VSS 8.41fF
C17983 nmat.col_n[4] VSS 8.40fF
C17984 nmat.col[4] VSS 6.46fF
C17985 nmat.col_n[2] VSS 8.42fF
C17986 a_12061_26703# VSS 1.22fF
C17987 a_19746_28111# VSS 0.49fF
C17988 a_17323_28111# VSS 0.59fF
C17989 a_20164_27791# VSS 0.41fF
C17990 a_12987_26159# VSS 1.14fF
C17991 a_17845_27791# VSS 0.47fF
C17992 _0467_ VSS 1.62fF
C17993 a_7026_24527# VSS 3.03fF
C17994 nmat.col[7] VSS 8.23fF
C17995 a_8951_27907# VSS 0.32fF
C17996 a_2683_22089# VSS 2.87fF
C17997 a_7023_27907# VSS 0.32fF
C17998 a_7140_27805# VSS 0.51fF
C17999 a_2283_27221# VSS 0.53fF
C18000 a_3305_27791# VSS 2.37fF
C18001 a_2564_21959# VSS 2.88fF
C18002 a_2847_28095# VSS 0.59fF
C18003 a_1895_27962# VSS 0.34fF
C18004 a_1591_27797# VSS 0.47fF
C18005 ANTENNA__1190__A2.DIODE VSS 16.37fF
C18006 nmat.col[28] VSS 13.72fF
C18007 nmat.col[21] VSS 15.08fF
C18008 inn_analog VSS 13.67fF
C18009 nmat.col_n[30] VSS 27.08fF
C18010 nmat.col_n[31] VSS 32.39fF
C18011 nmat.col_n[18] VSS 20.65fF
C18012 nmat.col[13] VSS 8.35fF
C18013 a_27763_27221# VSS 1.94fF
C18014 nmat.en_bit_n[2] VSS 1.29fF
C18015 a_12053_27497# VSS 5.45fF
C18016 a_46863_28585# VSS 0.43fF
C18017 a_10223_26703# VSS 3.73fF
C18018 nmat.en_C0_n VSS 1.42fF
C18019 a_9075_28023# VSS 0.96fF
C18020 a_5991_23983# VSS 2.78fF
C18021 a_7840_27247# VSS 2.59fF
C18022 a_11927_27399# VSS 2.75fF
C18023 a_12175_27221# VSS 0.57fF
C18024 a_12155_27791# VSS 0.32fF
C18025 a_5351_19913# VSS 9.14fF
C18026 a_5331_28309# VSS 0.46fF
C18027 a_4075_28335# VSS 0.58fF
C18028 a_46395_29199# VSS 0.48fF
C18029 a_44463_29199# VSS 0.48fF
C18030 nmat.col[24] VSS 13.72fF
C18031 nmat.col_n[28] VSS 21.94fF
C18032 nmat.col[29] VSS 21.32fF
C18033 a_27355_28995# VSS 0.32fF
C18034 nmat.col_n[13] VSS 9.77fF
C18035 a_22015_28995# VSS 0.30fF
C18036 nmat.col[0] VSS 6.70fF
C18037 a_19083_28879# VSS 0.47fF
C18038 nmat.col_n[7] VSS 11.64fF
C18039 a_10589_22351# VSS 0.52fF
C18040 a_12437_28585# VSS 0.67fF
C18041 nmat.col_n[3] VSS 10.58fF
C18042 a_10957_28879# VSS 1.10fF
C18043 a_10609_28995# VSS 0.31fF
C18044 a_10814_29111# VSS 1.16fF
C18045 a_9741_28585# VSS 1.04fF
C18046 a_9395_27791# VSS 0.96fF
C18047 a_9323_28879# VSS 0.49fF
C18048 a_4516_21531# VSS 3.35fF
C18049 a_4068_25615# VSS 5.79fF
C18050 a_1586_18231# VSS 5.81fF
C18051 a_3351_27249# VSS 1.89fF
C18052 a_4679_28853# VSS 0.31fF
C18053 a_3944_28853# VSS 0.32fF
C18054 a_2743_28853# VSS 0.38fF
C18055 a_47043_29423# VSS 0.32fF
C18056 a_43659_28853# VSS 0.97fF
C18057 a_37237_29423# VSS 0.32fF
C18058 nmat.col[30] VSS 14.42fF
C18059 nmat.col[12] VSS 8.31fF
C18060 nmat.col_n[10] VSS 10.54fF
C18061 a_17830_29423# VSS 0.73fF
C18062 a_16966_29423# VSS 0.49fF
C18063 a_21365_27247# VSS 1.44fF
C18064 a_19405_28853# VSS 0.72fF
C18065 a_8443_20719# VSS 2.53fF
C18066 a_14943_26703# VSS 0.77fF
C18067 a_47212_29673# VSS 0.43fF
C18068 a_41703_29423# VSS 0.45fF
C18069 a_41443_28879# VSS 0.68fF
C18070 a_41237_28585# VSS 0.34fF
C18071 a_36453_29199# VSS 0.49fF
C18072 a_31217_29429# VSS 0.31fF
C18073 a_28626_29423# VSS 0.34fF
C18074 a_27794_28879# VSS 0.79fF
C18075 a_15667_28111# VSS 0.65fF
C18076 a_16478_29423# VSS 0.39fF
C18077 a_22307_27791# VSS 1.84fF
C18078 a_16966_29673# VSS 0.42fF
C18079 a_17306_28879# VSS 0.79fF
C18080 a_12437_28879# VSS 0.78fF
C18081 a_13655_26703# VSS 0.63fF
C18082 a_14466_28879# VSS 0.37fF
C18083 a_14691_29575# VSS 0.98fF
C18084 a_6830_22895# VSS 3.70fF
C18085 a_4339_27804# VSS 2.44fF
C18086 a_2952_25045# VSS 4.43fF
C18087 a_6981_28879# VSS 0.52fF
C18088 dummypin[8] VSS 0.92fF
C18089 adc_top_89.HI VSS 0.34fF
C18090 a_35559_30209# VSS 0.43fF
C18091 a_35039_29941# VSS 0.38fF
C18092 a_20439_27247# VSS 2.12fF
C18093 a_33011_29941# VSS 0.59fF
C18094 a_27995_30287# VSS 1.23fF
C18095 a_30699_29397# VSS 0.57fF
C18096 a_30603_29575# VSS 0.86fF
C18097 a_28812_29575# VSS 0.87fF
C18098 a_25681_28879# VSS 1.95fF
C18099 a_28715_28879# VSS 0.49fF
C18100 a_25325_29125# VSS 0.46fF
C18101 a_24747_29967# VSS 1.51fF
C18102 a_24214_29967# VSS 0.30fF
C18103 a_23043_28335# VSS 0.34fF
C18104 a_22871_29967# VSS 0.54fF
C18105 a_18566_30287# VSS 0.75fF
C18106 a_17702_30287# VSS 0.49fF
C18107 a_17702_29967# VSS 0.44fF
C18108 a_12461_29673# VSS 1.22fF
C18109 a_10441_21263# VSS 1.47fF
C18110 a_14365_22351# VSS 0.54fF
C18111 a_7939_29967# VSS 0.41fF
C18112 a_3622_29967# VSS 0.55fF
C18113 a_3052_29967# VSS 0.35fF
C18114 a_2500_30345# VSS 0.35fF
C18115 a_2217_29973# VSS 0.39fF
C18116 a_2051_29973# VSS 0.41fF
C18117 a_43869_30511# VSS 0.36fF
C18118 a_45915_29941# VSS 1.08fF
C18119 ANTENNA__1183__B1.DIODE VSS 15.19fF
C18120 a_22576_30511# VSS 0.47fF
C18121 a_37827_30793# VSS 0.94fF
C18122 a_23021_29199# VSS 1.61fF
C18123 a_27001_30511# VSS 0.73fF
C18124 a_47685_30517# VSS 0.31fF
C18125 a_45405_30511# VSS 0.56fF
C18126 a_41227_29423# VSS 0.78fF
C18127 a_28336_29967# VSS 0.96fF
C18128 a_40969_30287# VSS 0.36fF
C18129 a_31399_30511# VSS 0.43fF
C18130 a_31323_29967# VSS 0.33fF
C18131 a_15753_28879# VSS 5.19fF
C18132 a_22186_30485# VSS 0.87fF
C18133 a_20695_30485# VSS 0.39fF
C18134 a_19439_30511# VSS 0.37fF
C18135 a_10147_29415# VSS 4.76fF
C18136 a_10287_29941# VSS 0.81fF
C18137 a_10851_30485# VSS 0.63fF
C18138 a_9899_30724# VSS 0.53fF
C18139 a_9595_30511# VSS 0.39fF
C18140 a_2648_29397# VSS 7.42fF
C18141 a_5423_30485# VSS 0.61fF
C18142 a_4167_30511# VSS 0.61fF
C18143 a_34204_27765# VSS 2.28fF
C18144 a_37291_29397# VSS 0.72fF
C18145 a_47011_31029# VSS 0.38fF
C18146 a_46339_31029# VSS 0.85fF
C18147 a_40125_31029# VSS 0.31fF
C18148 nmat.col_n[21] VSS 25.74fF
C18149 a_6664_26159# VSS 13.03fF
C18150 a_31263_28309# VSS 1.28fF
C18151 a_7415_29397# VSS 8.80fF
C18152 a_29493_31375# VSS 0.43fF
C18153 a_29455_31293# VSS 0.59fF
C18154 a_9785_28879# VSS 8.24fF
C18155 a_22459_28879# VSS 0.93fF
C18156 a_13641_23439# VSS 6.22fF
C18157 a_25575_31055# VSS 4.28fF
C18158 a_25042_31055# VSS 0.31fF
C18159 a_15101_29423# VSS 2.80fF
C18160 a_22628_30485# VSS 2.57fF
C18161 a_24160_30199# VSS 0.51fF
C18162 a_18563_27791# VSS 5.61fF
C18163 nmat.col[10] VSS 8.56fF
C18164 a_20310_28029# VSS 0.89fF
C18165 a_12851_28853# VSS 3.13fF
C18166 nmat.en_bit_n[0] VSS 6.14fF
C18167 a_15660_31029# VSS 0.49fF
C18168 a_13479_26935# VSS 1.66fF
C18169 a_13335_31359# VSS 0.51fF
C18170 a_5535_29980# VSS 1.73fF
C18171 a_12079_31061# VSS 0.42fF
C18172 a_7619_30485# VSS 0.41fF
C18173 a_9307_31068# VSS 0.68fF
C18174 a_7999_31359# VSS 0.48fF
C18175 a_6743_31061# VSS 0.42fF
C18176 a_4951_31029# VSS 0.50fF
C18177 a_17842_27497# VSS 7.11fF
C18178 a_30121_31599# VSS 0.32fF
C18179 nmat.col_n[12] VSS 13.12fF
C18180 a_8583_29199# VSS 5.63fF
C18181 a_25084_31287# VSS 0.31fF
C18182 a_14917_23983# VSS 0.85fF
C18183 a_14691_27399# VSS 0.45fF
C18184 nmat.rowon_n[5] VSS 4.45fF
C18185 a_15435_29111# VSS 1.03fF
C18186 a_47039_31599# VSS 0.95fF
C18187 a_45589_31599# VSS 0.52fF
C18188 a_41949_30761# VSS 0.73fF
C18189 a_42240_29423# VSS 0.74fF
C18190 a_42307_31756# VSS 0.82fF
C18191 a_38913_31055# VSS 0.58fF
C18192 a_39939_29967# VSS 0.65fF
C18193 a_37143_31573# VSS 0.36fF
C18194 a_33869_31599# VSS 0.35fF
C18195 a_31339_31787# VSS 1.56fF
C18196 a_31210_31751# VSS 0.40fF
C18197 a_30527_31573# VSS 0.31fF
C18198 a_30219_29967# VSS 0.39fF
C18199 a_28704_29568# VSS 1.49fF
C18200 a_20616_27791# VSS 2.46fF
C18201 a_24861_29673# VSS 1.27fF
C18202 a_21279_31599# VSS 0.50fF
C18203 a_16635_31573# VSS 0.84fF
C18204 a_15543_31573# VSS 0.41fF
C18205 a_14287_31599# VSS 0.58fF
C18206 a_2422_29575# VSS 0.55fF
C18207 a_2163_31741# VSS 0.43fF
C18208 a_1643_31573# VSS 0.40fF
C18209 a_38905_28853# VSS 2.17fF
C18210 a_45282_32143# VSS 1.63fF
C18211 a_44571_32143# VSS 0.70fF
C18212 a_42791_32375# VSS 0.44fF
C18213 a_43543_32151# VSS 0.33fF
C18214 a_18597_31599# VSS 2.30fF
C18215 a_41427_32143# VSS 0.50fF
C18216 a_40903_32375# VSS 0.39fF
C18217 a_40567_32403# VSS 0.52fF
C18218 a_38727_32447# VSS 0.54fF
C18219 a_37637_32149# VSS 0.32fF
C18220 a_37471_32149# VSS 0.51fF
C18221 a_33684_32143# VSS 0.48fF
C18222 a_34243_32143# VSS 0.49fF
C18223 a_33205_32143# VSS 0.33fF
C18224 a_32957_30287# VSS 0.76fF
C18225 a_29163_29423# VSS 0.65fF
C18226 a_30278_30511# VSS 0.47fF
C18227 a_32771_31599# VSS 0.44fF
C18228 a_31263_32117# VSS 1.88fF
C18229 a_9963_28111# VSS 6.42fF
C18230 a_27976_32463# VSS 0.32fF
C18231 a_27443_32143# VSS 0.30fF
C18232 a_24374_29941# VSS 1.35fF
C18233 a_27498_32117# VSS 0.76fF
C18234 a_26479_32117# VSS 3.66fF
C18235 a_25688_32117# VSS 0.33fF
C18236 a_23933_32143# VSS 1.08fF
C18237 a_18241_31698# VSS 2.01fF
C18238 a_23455_32447# VSS 0.54fF
C18239 a_2007_25597# VSS 10.14fF
C18240 a_22365_32149# VSS 0.32fF
C18241 a_22199_32149# VSS 0.49fF
C18242 a_20695_32447# VSS 0.52fF
C18243 a_19605_32149# VSS 0.30fF
C18244 a_19439_32149# VSS 0.48fF
C18245 a_7717_14735# VSS 7.56fF
C18246 nmat.rowoff_n[6] VSS 1.93fF
C18247 a_14839_20871# VSS 0.85fF
C18248 a_7939_31591# VSS 2.73fF
C18249 a_9983_32385# VSS 0.45fF
C18250 a_9231_32117# VSS 0.75fF
C18251 a_5179_31591# VSS 3.11fF
C18252 a_5963_32117# VSS 0.53fF
C18253 a_4707_32156# VSS 0.90fF
C18254 a_45277_32687# VSS 1.06fF
C18255 a_45119_32661# VSS 0.51fF
C18256 a_47499_32687# VSS 0.42fF
C18257 a_6343_32661# VSS 0.63fF
C18258 a_5391_32900# VSS 0.66fF
C18259 a_5087_32687# VSS 0.53fF
C18260 a_4123_32661# VSS 0.47fF
C18261 a_46386_33231# VSS 1.63fF
C18262 a_44888_33205# VSS 0.51fF
C18263 a_7387_33231# VSS 0.43fF
C18264 a_4043_33535# VSS 0.73fF
C18265 a_2787_33237# VSS 0.42fF
C18266 a_45908_33749# VSS 0.51fF
C18267 a_44533_33749# VSS 1.54fF
C18268 a_46994_34639# VSS 0.76fF
C18269 a_46130_34639# VSS 0.50fF
C18270 a_46130_34319# VSS 0.48fF
C18271 nmat.sample_n VSS 15.46fF
C18272 a_17808_34215# VSS 0.48fF
C18273 nmat.sample VSS 14.94fF
C18274 a_17867_34473# VSS 0.34fF
C18275 a_14864_34215# VSS 0.48fF
C18276 a_37823_34191# VSS 0.56fF
C18277 a_36946_34191# VSS 0.55fF
C18278 a_35382_34191# VSS 0.55fF
C18279 a_34002_34191# VSS 0.49fF
C18280 a_32162_34191# VSS 0.63fF
C18281 cgen.dlycontrol1_in[3] VSS 3.48fF
C18282 a_24667_34191# VSS 0.46fF
C18283 a_21815_34191# VSS 0.45fF
C18284 a_20711_34191# VSS 0.46fF
C18285 a_19834_34191# VSS 0.31fF
C18286 a_16745_34427# VSS 3.03fF
C18287 a_14923_34473# VSS 0.32fF
C18288 a_12196_34215# VSS 0.48fF
C18289 a_12255_34473# VSS 0.33fF
C18290 a_1923_31743# VSS 11.80fF
C18291 a_6007_33767# VSS 3.43fF
C18292 a_2847_33749# VSS 0.37fF
C18293 a_1591_33775# VSS 0.50fF
C18294 a_13801_34427# VSS 3.04fF
C18295 a_11133_34427# VSS 2.99fF
C18296 a_46522_34293# VSS 1.00fF
C18297 cgen.dlycontrol1_in[0] VSS 3.46fF
C18298 a_27687_34967# VSS 0.31fF
C18299 a_26767_34967# VSS 0.95fF
C18300 a_25628_35077# VSS 0.47fF
C18301 cgen.dlycontrol1_in[2] VSS 2.69fF
C18302 a_24565_34789# VSS 2.86fF
C18303 a_20752_35077# VSS 0.46fF
C18304 a_19689_34789# VSS 2.93fF
C18305 a_18176_35077# VSS 0.44fF
C18306 a_17113_34789# VSS 2.87fF
C18307 a_15048_35077# VSS 0.43fF
C18308 a_15144_35077# VSS 1.71fF
C18309 a_13985_34789# VSS 2.93fF
C18310 a_13529_34951# VSS 2.30fF
C18311 a_12472_35077# VSS 0.43fF
C18312 a_4831_34561# VSS 0.37fF
C18313 a_4227_34293# VSS 0.47fF
C18314 a_2511_34319# VSS 0.40fF
C18315 a_1858_25615# VSS 8.19fF
C18316 a_12568_35077# VSS 1.72fF
C18317 a_11409_34789# VSS 2.78fF
C18318 a_10953_34951# VSS 1.65fF
C18319 a_45107_34863# VSS 0.45fF
C18320 a_47591_35407# VSS 0.46fF
C18321 a_45829_35407# VSS 0.75fF
C18322 a_28112_35303# VSS 0.49fF
C18323 a_28171_35561# VSS 0.32fF
C18324 a_27049_35515# VSS 3.14fF
C18325 a_22684_35303# VSS 0.47fF
C18326 a_22743_35561# VSS 0.30fF
C18327 a_17900_35303# VSS 0.44fF
C18328 a_25667_35253# VSS 0.41fF
C18329 a_23655_35279# VSS 0.41fF
C18330 a_21621_35515# VSS 2.81fF
C18331 a_20534_35431# VSS 3.43fF
C18332 a_19086_34343# VSS 0.43fF
C18333 a_17959_35561# VSS 0.32fF
C18334 a_16381_35286# VSS 2.33fF
C18335 a_17996_35303# VSS 1.49fF
C18336 a_16837_35515# VSS 2.96fF
C18337 a_13345_35303# VSS 0.47fF
C18338 a_14589_35286# VSS 1.75fF
C18339 a_13259_35561# VSS 0.30fF
C18340 a_10677_35303# VSS 0.47fF
C18341 a_7079_34837# VSS 0.64fF
C18342 a_6127_35076# VSS 0.83fF
C18343 a_5823_34863# VSS 0.50fF
C18344 a_1775_35113# VSS 0.41fF
C18345 a_11921_35286# VSS 2.49fF
C18346 a_10591_35561# VSS 0.32fF
C18347 a_13653_35516# VSS 2.92fF
C18348 a_10985_35516# VSS 2.89fF
C18349 a_10651_35507# VSS 1.59fF
C18350 a_44763_34293# VSS 0.70fF
C18351 a_47592_35643# VSS 0.41fF
C18352 a_35799_35831# VSS 0.32fF
C18353 a_35885_36165# VSS 0.45fF
C18354 a_36193_35805# VSS 3.26fF
C18355 a_34828_36165# VSS 0.43fF
C18356 a_33765_35877# VSS 2.96fF
C18357 a_25755_34343# VSS 3.42fF
C18358 a_26583_34343# VSS 0.95fF
C18359 a_29308_36165# VSS 0.44fF
C18360 a_26515_35831# VSS 0.33fF
C18361 cgen.dlycontrol1_in[1] VSS 2.37fF
C18362 a_28245_35877# VSS 3.10fF
C18363 a_27789_36039# VSS 1.50fF
C18364 a_26456_36165# VSS 0.48fF
C18365 a_26552_36165# VSS 1.30fF
C18366 a_25393_35877# VSS 2.96fF
C18367 a_24937_36039# VSS 1.38fF
C18368 a_23420_36165# VSS 0.47fF
C18369 a_22357_35877# VSS 2.88fF
C18370 a_20752_36165# VSS 0.47fF
C18371 a_18235_35831# VSS 0.32fF
C18372 a_20848_36165# VSS 1.14fF
C18373 a_19689_35877# VSS 3.00fF
C18374 a_18272_35077# VSS 1.66fF
C18375 a_18176_36165# VSS 0.48fF
C18376 a_17113_35877# VSS 2.90fF
C18377 a_15048_36165# VSS 0.44fF
C18378 a_15144_36165# VSS 1.61fF
C18379 a_13985_35877# VSS 2.90fF
C18380 a_13319_35507# VSS 1.21fF
C18381 a_11681_35823# VSS 0.81fF
C18382 a_2046_30184# VSS 11.31fF
C18383 a_5271_35407# VSS 0.38fF
C18384 a_4601_35727# VSS 0.36fF
C18385 a_4267_35407# VSS 0.35fF
C18386 a_4307_35639# VSS 0.33fF
C18387 a_11297_36091# VSS 2.60fF
C18388 a_11057_35836# VSS 2.84fF
C18389 a_40951_31599# VSS 1.67fF
C18390 a_37680_36391# VSS 0.50fF
C18391 a_37739_36649# VSS 0.39fF
C18392 a_34552_36391# VSS 0.49fF
C18393 a_34924_36165# VSS 1.91fF
C18394 a_44423_36815# VSS 0.51fF
C18395 a_37129_36130# VSS 1.74fF
C18396 a_36617_36603# VSS 3.23fF
C18397 a_34611_36649# VSS 0.33fF
C18398 a_31976_36391# VSS 0.47fF
C18399 a_33309_36039# VSS 1.72fF
C18400 a_33489_36603# VSS 3.10fF
C18401 a_32035_36649# VSS 0.33fF
C18402 a_29404_36165# VSS 1.83fF
C18403 a_30913_36603# VSS 2.99fF
C18404 a_28247_34191# VSS 0.93fF
C18405 a_24833_34191# VSS 1.78fF
C18406 a_27560_36391# VSS 0.50fF
C18407 a_28431_34735# VSS 0.62fF
C18408 a_27619_36649# VSS 0.35fF
C18409 a_26497_36603# VSS 3.20fF
C18410 a_23604_36391# VSS 0.48fF
C18411 a_23663_36649# VSS 0.32fF
C18412 a_21028_36391# VSS 0.44fF
C18413 a_22085_36374# VSS 1.52fF
C18414 a_23700_36391# VSS 1.30fF
C18415 a_22541_36603# VSS 2.91fF
C18416 a_21087_36649# VSS 0.31fF
C18417 a_17900_36391# VSS 0.45fF
C18418 a_21124_36391# VSS 1.59fF
C18419 a_19965_36603# VSS 2.97fF
C18420 a_17959_36649# VSS 0.33fF
C18421 a_17996_36391# VSS 1.44fF
C18422 a_16837_36603# VSS 3.05fF
C18423 a_13805_36391# VSS 0.48fF
C18424 a_15049_36374# VSS 1.53fF
C18425 a_13719_36649# VSS 0.31fF
C18426 a_14113_36604# VSS 2.97fF
C18427 a_13779_36595# VSS 1.37fF
C18428 a_12309_36483# VSS 0.83fF
C18429 a_12069_36341# VSS 2.26fF
C18430 a_11225_35836# VSS 1.79fF
C18431 cgen.dlycontrol1_in[4] VSS 1.98fF
C18432 a_11113_36483# VSS 1.27fF
C18433 a_11041_36596# VSS 1.46fF
C18434 a_10873_36341# VSS 3.35fF
C18435 a_47207_35951# VSS 0.73fF
C18436 a_46636_36469# VSS 0.58fF
C18437 a_45625_36495# VSS 0.33fF
C18438 a_34887_36919# VSS 0.31fF
C18439 a_40399_36911# VSS 0.48fF
C18440 a_34828_37253# VSS 0.44fF
C18441 a_33765_36965# VSS 3.02fF
C18442 a_31425_37218# VSS 1.47fF
C18443 a_30095_36919# VSS 0.33fF
C18444 a_29183_36919# VSS 0.30fF
C18445 a_30181_37253# VSS 0.48fF
C18446 a_30489_36893# VSS 2.99fF
C18447 a_30155_36893# VSS 1.39fF
C18448 a_29124_37253# VSS 0.44fF
C18449 a_26331_36919# VSS 0.32fF
C18450 a_28061_36965# VSS 3.17fF
C18451 a_27605_37127# VSS 1.50fF
C18452 a_26272_37253# VSS 0.49fF
C18453 a_26041_36374# VSS 1.34fF
C18454 a_25209_36965# VSS 3.15fF
C18455 a_22537_36911# VSS 1.24fF
C18456 a_19891_36919# VSS 0.31fF
C18457 a_19832_37253# VSS 0.44fF
C18458 a_18769_36965# VSS 3.07fF
C18459 a_16890_36911# VSS 0.68fF
C18460 a_14773_37218# VSS 2.04fF
C18461 a_13443_36919# VSS 0.31fF
C18462 a_13529_37253# VSS 0.47fF
C18463 a_17675_37001# VSS 0.80fF
C18464 a_12934_35823# VSS 0.38fF
C18465 a_13837_36893# VSS 2.91fF
C18466 a_13503_36893# VSS 1.37fF
C18467 a_12237_36596# VSS 0.94fF
C18468 a_2847_36799# VSS 0.41fF
C18469 a_1895_36666# VSS 0.38fF
C18470 a_1591_36501# VSS 0.54fF
C18471 a_12585_37179# VSS 0.80fF
C18472 a_12345_36924# VSS 1.62fF
C18473 a_11317_36924# VSS 3.30fF
C18474 a_11149_36924# VSS 5.68fF
C18475 a_35244_32411# VSS 6.43fF
C18476 a_43776_30287# VSS 2.19fF
C18477 a_43533_30761# VSS 3.01fF
C18478 a_46815_37013# VSS 0.52fF
C18479 a_44811_36469# VSS 1.11fF
C18480 a_38737_37479# VSS 0.48fF
C18481 a_37680_37479# VSS 0.45fF
C18482 a_38651_37737# VSS 0.32fF
C18483 a_39045_37692# VSS 2.89fF
C18484 a_37739_37737# VSS 0.32fF
C18485 a_36617_37691# VSS 3.00fF
C18486 a_33033_37479# VSS 0.49fF
C18487 a_32947_37737# VSS 0.32fF
C18488 a_33341_37692# VSS 3.00fF
C18489 a_33007_37683# VSS 1.45fF
C18490 a_30457_37479# VSS 0.47fF
C18491 a_30371_37737# VSS 0.31fF
C18492 a_30765_37692# VSS 2.99fF
C18493 a_28020_37479# VSS 0.46fF
C18494 a_28079_37737# VSS 0.33fF
C18495 a_26957_37691# VSS 3.30fF
C18496 a_24015_36911# VSS 0.36fF
C18497 a_21219_36885# VSS 1.42fF
C18498 a_22085_37479# VSS 0.47fF
C18499 a_21999_37737# VSS 0.30fF
C18500 a_22393_37692# VSS 2.88fF
C18501 a_22059_37683# VSS 2.38fF
C18502 a_19509_37479# VSS 0.42fF
C18503 a_19928_37253# VSS 1.77fF
C18504 a_19423_37737# VSS 0.31fF
C18505 a_19817_37692# VSS 2.88fF
C18506 a_15737_37479# VSS 0.43fF
C18507 a_16981_37462# VSS 1.94fF
C18508 a_16045_37692# VSS 2.90fF
C18509 a_14712_37429# VSS 1.45fF
C18510 a_14719_37737# VSS 0.64fF
C18511 a_14600_37607# VSS 2.03fF
C18512 a_12513_36924# VSS 1.53fF
C18513 a_10677_37479# VSS 0.48fF
C18514 a_7355_37013# VSS 0.42fF
C18515 a_6099_37039# VSS 0.40fF
C18516 a_2467_35925# VSS 0.38fF
C18517 cgen.dlycontrol2_in[0] VSS 3.80fF
C18518 a_4031_37191# VSS 0.32fF
C18519 a_13597_37571# VSS 2.89fF
C18520 a_13357_37429# VSS 1.31fF
C18521 a_11921_37462# VSS 3.97fF
C18522 a_10591_37737# VSS 0.33fF
C18523 a_10985_37692# VSS 2.93fF
C18524 a_10651_37683# VSS 0.88fF
C18525 a_45187_38129# VSS 0.82fF
C18526 a_40532_38341# VSS 0.48fF
C18527 a_37463_38007# VSS 0.32fF
C18528 a_39981_37462# VSS 1.28fF
C18529 a_39469_38053# VSS 2.89fF
C18530 a_37776_37479# VSS 1.58fF
C18531 a_37404_38341# VSS 0.49fF
C18532 a_34887_38007# VSS 0.30fF
C18533 a_36161_37462# VSS 2.45fF
C18534 a_36341_38053# VSS 3.14fF
C18535 a_34924_37253# VSS 1.59fF
C18536 a_34828_38341# VSS 0.47fF
C18537 a_34277_37462# VSS 1.28fF
C18538 a_33765_38053# VSS 2.92fF
C18539 a_30431_37683# VSS 1.44fF
C18540 a_31976_38341# VSS 0.45fF
C18541 a_31701_37462# VSS 1.24fF
C18542 a_30913_38053# VSS 2.93fF
C18543 a_29220_37253# VSS 1.55fF
C18544 a_28116_37479# VSS 1.70fF
C18545 a_27795_38007# VSS 0.33fF
C18546 a_26515_38007# VSS 0.31fF
C18547 a_27881_38341# VSS 0.45fF
C18548 a_28189_37981# VSS 3.01fF
C18549 a_26456_38341# VSS 0.47fF
C18550 a_23847_38007# VSS 0.30fF
C18551 a_26501_37462# VSS 1.30fF
C18552 a_25393_38053# VSS 2.95fF
C18553 a_23788_38341# VSS 0.47fF
C18554 a_23329_37462# VSS 1.19fF
C18555 a_22725_38053# VSS 2.87fF
C18556 a_20752_38341# VSS 0.43fF
C18557 a_18143_38007# VSS 0.30fF
C18558 a_20848_38341# VSS 1.47fF
C18559 a_19689_38053# VSS 2.90fF
C18560 a_19233_38215# VSS 1.45fF
C18561 a_18084_38341# VSS 0.48fF
C18562 a_18180_38341# VSS 1.37fF
C18563 a_17021_38053# VSS 2.88fF
C18564 a_14773_38306# VSS 1.43fF
C18565 a_13529_38341# VSS 0.47fF
C18566 a_13837_37981# VSS 2.85fF
C18567 a_13503_37981# VSS 1.42fF
C18568 a_12197_38306# VSS 2.15fF
C18569 a_10867_38007# VSS 0.32fF
C18570 a_6403_37252# VSS 0.38fF
C18571 a_4127_37013# VSS 0.57fF
C18572 a_10953_38341# VSS 0.48fF
C18573 a_11261_37981# VSS 2.90fF
C18574 a_47357_38127# VSS 0.66fF
C18575 a_45325_38127# VSS 0.57fF
C18576 vcm.sky130_fd_sc_hd__buf_4_3.X VSS 0.69fF
C18577 vcm.sky130_fd_sc_hd__buf_4_2.X VSS 1.28fF
C18578 a_77980_38962# VSS 0.47fF
C18579 a_77428_38962# VSS 0.45fF
C18580 vcm.sky130_fd_sc_hd__buf_4_2.A VSS 0.47fF
C18581 a_45866_38279# VSS 0.66fF
C18582 a_47223_38671# VSS 0.48fF
C18583 a_39197_38567# VSS 0.44fF
C18584 a_38711_37683# VSS 2.68fF
C18585 a_39505_38780# VSS 2.84fF
C18586 a_22153_37179# VSS 2.01fF
C18587 a_36253_38567# VSS 0.51fF
C18588 a_36167_38825# VSS 0.35fF
C18589 a_36561_38780# VSS 3.08fF
C18590 a_33033_38567# VSS 0.48fF
C18591 a_31976_38567# VSS 0.44fF
C18592 a_32947_38825# VSS 0.32fF
C18593 a_33341_38780# VSS 2.94fF
C18594 a_32035_38825# VSS 0.31fF
C18595 a_28020_38567# VSS 0.49fF
C18596 a_30913_38779# VSS 2.92fF
C18597 a_28079_38825# VSS 0.33fF
C18598 a_26957_38779# VSS 3.12fF
C18599 a_23604_38567# VSS 0.43fF
C18600 a_23663_38825# VSS 0.30fF
C18601 a_20568_38567# VSS 0.48fF
C18602 a_23700_38567# VSS 1.39fF
C18603 a_22541_38779# VSS 2.92fF
C18604 a_20627_38825# VSS 0.31fF
C18605 a_17440_38567# VSS 0.45fF
C18606 a_19505_38779# VSS 2.93fF
C18607 a_17499_38825# VSS 0.31fF
C18608 a_14864_38567# VSS 0.48fF
C18609 a_17536_38567# VSS 1.64fF
C18610 a_16377_38779# VSS 2.82fF
C18611 a_14923_38825# VSS 0.31fF
C18612 a_10927_37981# VSS 1.36fF
C18613 a_13801_38779# VSS 2.84fF
C18614 a_12693_38543# VSS 0.59fF
C18615 a_6061_38377# VSS 0.55fF
C18616 a_2563_34837# VSS 0.88fF
C18617 a_3325_36495# VSS 1.46fF
C18618 cgen.dlycontrol2_in[1] VSS 3.09fF
C18619 a_4535_38377# VSS 0.40fF
C18620 a_11113_38659# VSS 0.69fF
C18621 a_11041_38772# VSS 3.09fF
C18622 a_44515_38645# VSS 0.56fF
C18623 vcm.sky130_fd_sc_hd__dlymetal6s6s_1_5.X VSS 0.52fF
C18624 a_54790_39198# VSS 0.52fF
C18625 vcm.sky130_fd_sc_hd__nand2_1_1.Y VSS 0.31fF
C18626 a_44789_39215# VSS 0.36fF
C18627 a_40532_39429# VSS 0.43fF
C18628 a_37463_39095# VSS 0.30fF
C18629 a_39469_39141# VSS 2.89fF
C18630 a_37404_39429# VSS 0.45fF
C18631 a_34887_39095# VSS 0.30fF
C18632 a_37497_38550# VSS 1.52fF
C18633 a_36341_39141# VSS 3.15fF
C18634 a_34828_39429# VSS 0.47fF
C18635 a_34277_38550# VSS 1.28fF
C18636 a_33765_39141# VSS 2.87fF
C18637 a_32072_38567# VSS 1.59fF
C18638 a_29159_37607# VSS 0.64fF
C18639 a_10873_38517# VSS 2.71fF
C18640 a_27603_34191# VSS 0.60fF
C18641 a_29768_39429# VSS 0.43fF
C18642 a_29864_39429# VSS 1.28fF
C18643 a_28705_39141# VSS 2.96fF
C18644 a_28116_38567# VSS 1.33fF
C18645 a_25755_38695# VSS 0.44fF
C18646 a_26180_39429# VSS 0.48fF
C18647 a_26276_39429# VSS 1.23fF
C18648 a_25117_39141# VSS 2.95fF
C18649 a_23420_39429# VSS 0.47fF
C18650 a_22085_38550# VSS 1.36fF
C18651 a_22357_39141# VSS 2.92fF
C18652 a_20752_39429# VSS 0.43fF
C18653 a_20848_39429# VSS 1.41fF
C18654 a_19689_39141# VSS 3.02fF
C18655 a_18176_39429# VSS 0.44fF
C18656 a_18272_39429# VSS 1.47fF
C18657 a_17113_39141# VSS 2.81fF
C18658 a_14773_39394# VSS 1.37fF
C18659 a_13529_39429# VSS 0.46fF
C18660 a_13837_39069# VSS 2.80fF
C18661 a_13503_39069# VSS 1.83fF
C18662 a_2847_38975# VSS 0.64fF
C18663 a_1591_38677# VSS 0.51fF
C18664 a_12513_39100# VSS 1.34fF
C18665 a_12585_39355# VSS 0.74fF
C18666 comp.adc_inverter_1.in VSS 2.75fF
C18667 a_46947_39215# VSS 0.94fF
C18668 a_46705_38671# VSS 0.57fF
C18669 a_52398_39208# VSS 0.77fF
C18670 clk_vcm VSS 3.33fF
C18671 vcm.sky130_fd_sc_hd__buf_4_3.A VSS 0.99fF
C18672 vcm.sky130_fd_sc_hd__nand2_1_0.Y VSS 0.44fF
C18673 comp.adc_nor_latch_0.QN VSS 0.85fF
C18674 comp.adc_nor_latch_0.NOR_1/A VSS 0.93fF
C18675 a_38876_39655# VSS 0.48fF
C18676 a_45019_38645# VSS 4.20fF
C18677 a_46523_39733# VSS 0.92fF
C18678 a_38935_39913# VSS 0.33fF
C18679 a_35012_39655# VSS 0.43fF
C18680 a_36227_38771# VSS 1.62fF
C18681 a_38972_39655# VSS 1.27fF
C18682 a_37813_39867# VSS 3.08fF
C18683 a_35071_39913# VSS 0.32fF
C18684 a_31976_39655# VSS 0.48fF
C18685 a_33007_38771# VSS 1.37fF
C18686 a_35108_39655# VSS 1.50fF
C18687 a_33949_39867# VSS 2.93fF
C18688 a_32035_39913# VSS 0.32fF
C18689 a_30913_39867# VSS 2.91fF
C18690 a_28020_39655# VSS 0.48fF
C18691 a_23821_35279# VSS 1.97fF
C18692 a_29159_39783# VSS 1.56fF
C18693 a_12345_39100# VSS 1.67fF
C18694 a_28079_39913# VSS 0.32fF
C18695 a_26957_39867# VSS 3.15fF
C18696 a_23604_39655# VSS 0.44fF
C18697 a_23663_39913# VSS 0.30fF
C18698 a_21028_39655# VSS 0.44fF
C18699 a_23700_39655# VSS 1.47fF
C18700 a_22541_39867# VSS 2.95fF
C18701 a_21087_39913# VSS 0.30fF
C18702 a_19509_39638# VSS 1.57fF
C18703 a_21124_39655# VSS 1.38fF
C18704 a_19965_39867# VSS 2.81fF
C18705 a_16612_39655# VSS 0.47fF
C18706 a_16671_39913# VSS 0.31fF
C18707 a_15549_39867# VSS 2.84fF
C18708 a_12228_39605# VSS 1.86fF
C18709 a_1895_38842# VSS 0.69fF
C18710 a_4533_38279# VSS 2.27fF
C18711 a_2283_39189# VSS 0.37fF
C18712 comp.adc_comp_circuit_0.adc_comp_buffer_1.in VSS 1.30fF
C18713 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_0.nmoscap_top VSS 91.52fF
C18714 comp.adc_inverter_1.out VSS 1.54fF
C18715 comp.adc_nor_latch_0.R VSS 0.96fF
C18716 comp.adc_comp_circuit_0.adc_comp_buffer_0.in VSS 1.10fF
C18717 a_54790_39936# VSS 0.36fF
C18718 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_bot VSS 740.70fF
C18719 vcm.adc_noise_decoup_cell1_3[7|4].mimcap_top VSS 199.81fF
C18720 vcm.adc_noise_decoup_cell1_1[7|4].mimcap_top VSS 1474.07fF
C18721 vcm.sky130_fd_sc_hd__buf_4_1.X VSS 0.94fF
C18722 a_40628_39429# VSS 1.58fF
C18723 a_39387_40183# VSS 0.31fF
C18724 a_39473_40517# VSS 0.44fF
C18725 a_39781_40157# VSS 2.99fF
C18726 a_12309_38659# VSS 3.43fF
C18727 a_34828_40517# VSS 0.47fF
C18728 a_33765_40229# VSS 2.96fF
C18729 a_29163_38545# VSS 0.53fF
C18730 a_29735_40183# VSS 0.30fF
C18731 a_29676_40517# VSS 0.47fF
C18732 a_26423_40183# VSS 0.30fF
C18733 a_29772_40517# VSS 1.17fF
C18734 a_28613_40229# VSS 3.01fF
C18735 a_28116_39655# VSS 1.23fF
C18736 a_26364_40517# VSS 0.47fF
C18737 a_26460_40517# VSS 1.23fF
C18738 a_25301_40229# VSS 2.92fF
C18739 a_23788_40517# VSS 0.43fF
C18740 a_23884_40517# VSS 1.42fF
C18741 a_22725_40229# VSS 2.87fF
C18742 a_20476_40517# VSS 0.43fF
C18743 a_19413_40229# VSS 2.93fF
C18744 a_17441_40482# VSS 1.01fF
C18745 a_16111_40183# VSS 0.31fF
C18746 a_16197_40517# VSS 0.47fF
C18747 a_16505_40157# VSS 2.94fF
C18748 a_15048_40517# VSS 0.46fF
C18749 a_15093_39638# VSS 1.12fF
C18750 a_13985_40229# VSS 2.88fF
C18751 a_11773_39087# VSS 1.98fF
C18752 a_12969_40175# VSS 0.43fF
C18753 a_5687_38279# VSS 0.49fF
C18754 a_11565_39061# VSS 0.38fF
C18755 a_12585_40443# VSS 0.51fF
C18756 a_11339_39319# VSS 0.70fF
C18757 a_46897_40303# VSS 0.71fF
C18758 a_77980_40594# VSS 0.47fF
C18759 vcm.sky130_fd_sc_hd__nand2_1_1.A VSS 1.36fF
C18760 a_77428_40594# VSS 0.45fF
C18761 vcm.sky130_fd_sc_hd__buf_4_0.A VSS 0.46fF
C18762 vcm.sky130_fd_sc_hd__dlymetal6s6s_1_3.X VSS 0.52fF
C18763 vcm.sky130_fd_sc_hd__buf_4_0.X VSS 1.63fF
C18764 a_44444_32233# VSS 3.33fF
C18765 a_45246_41167# VSS 0.73fF
C18766 a_39105_40743# VSS 0.48fF
C18767 a_32988_40743# VSS 0.48fF
C18768 a_39019_41001# VSS 0.32fF
C18769 a_44382_41167# VSS 0.50fF
C18770 a_39413_40956# VSS 2.92fF
C18771 a_33047_41001# VSS 0.33fF
C18772 a_31469_40726# VSS 1.40fF
C18773 a_33084_40743# VSS 1.34fF
C18774 a_31925_40955# VSS 2.96fF
C18775 a_27836_40743# VSS 0.49fF
C18776 a_28975_40871# VSS 0.59fF
C18777 a_13909_39605# VSS 1.89fF
C18778 a_27895_41001# VSS 0.33fF
C18779 a_26773_40955# VSS 3.07fF
C18780 a_25671_40719# VSS 0.41fF
C18781 a_22684_40743# VSS 0.48fF
C18782 a_22743_41001# VSS 0.32fF
C18783 a_24667_40719# VSS 0.38fF
C18784 a_22269_40391# VSS 1.28fF
C18785 a_21621_40955# VSS 2.82fF
C18786 a_20605_40719# VSS 0.81fF
C18787 a_20221_40835# VSS 2.78fF
C18788 a_19409_40719# VSS 1.13fF
C18789 a_17900_40743# VSS 0.45fF
C18790 a_17959_41001# VSS 0.33fF
C18791 a_16171_40157# VSS 1.33fF
C18792 a_14533_39631# VSS 0.99fF
C18793 a_18975_40871# VSS 1.02fF
C18794 a_17996_40743# VSS 1.56fF
C18795 a_16837_40955# VSS 2.97fF
C18796 a_13345_40743# VSS 0.43fF
C18797 a_14589_40726# VSS 2.30fF
C18798 a_13653_40956# VSS 2.91fF
C18799 a_12235_39913# VSS 0.64fF
C18800 a_7079_40277# VSS 0.68fF
C18801 a_6127_40516# VSS 0.71fF
C18802 a_5823_40303# VSS 0.44fF
C18803 a_5233_40553# VSS 0.93fF
C18804 a_2839_38101# VSS 2.42fF
C18805 cgen.dlycontrol2_in[2] VSS 2.53fF
C18806 a_4705_39759# VSS 0.48fF
C18807 a_3295_40277# VSS 0.42fF
C18808 a_44382_40847# VSS 0.63fF
C18809 a_35312_31599# VSS 3.51fF
C18810 comp.adc_comp_circuit_0.adc_noise_decoup_cell2_1.nmoscap_top VSS 88.59fF
C18811 a_39387_41271# VSS 0.33fF
C18812 a_34887_41271# VSS 0.31fF
C18813 a_39473_41605# VSS 0.45fF
C18814 a_39781_41245# VSS 2.98fF
C18815 a_34828_41605# VSS 0.47fF
C18816 a_33765_41317# VSS 2.98fF
C18817 a_31793_41570# VSS 2.42fF
C18818 a_30463_41271# VSS 0.32fF
C18819 a_30549_41605# VSS 0.48fF
C18820 a_30857_41245# VSS 2.99fF
C18821 a_27887_41271# VSS 0.34fF
C18822 a_26515_41271# VSS 0.33fF
C18823 a_27973_41605# VSS 0.50fF
C18824 a_28281_41245# VSS 3.12fF
C18825 a_26456_41605# VSS 0.48fF
C18826 a_23939_41271# VSS 0.31fF
C18827 a_26317_40726# VSS 1.29fF
C18828 a_25393_41317# VSS 3.00fF
C18829 a_23880_41605# VSS 0.48fF
C18830 a_20811_41271# VSS 0.30fF
C18831 a_22817_41317# VSS 3.06fF
C18832 a_20752_41605# VSS 0.44fF
C18833 a_18235_41271# VSS 0.33fF
C18834 a_19689_41317# VSS 2.91fF
C18835 a_18176_41605# VSS 0.49fF
C18836 a_15107_41271# VSS 0.31fF
C18837 a_17113_41317# VSS 2.99fF
C18838 a_15048_41605# VSS 0.48fF
C18839 a_13985_41317# VSS 2.93fF
C18840 a_12197_41570# VSS 1.23fF
C18841 a_10867_41271# VSS 0.33fF
C18842 a_3659_39733# VSS 0.56fF
C18843 a_3325_40847# VSS 0.73fF
C18844 a_2847_41151# VSS 0.38fF
C18845 a_2411_33749# VSS 6.65fF
C18846 a_1591_40853# VSS 0.52fF
C18847 a_10953_41605# VSS 0.48fF
C18848 a_11261_41245# VSS 2.99fF
C18849 a_10927_41245# VSS 0.58fF
C18850 a_40256_41831# VSS 0.45fF
C18851 a_40315_42089# VSS 0.31fF
C18852 a_37680_41831# VSS 0.50fF
C18853 a_46753_41935# VSS 1.39fF
C18854 a_32405_32463# VSS 2.22fF
C18855 a_40352_41831# VSS 1.73fF
C18856 a_39193_42043# VSS 2.98fF
C18857 a_37739_42089# VSS 0.35fF
C18858 a_34552_41831# VSS 0.49fF
C18859 a_34924_41605# VSS 1.76fF
C18860 a_11113_40835# VSS 1.69fF
C18861 a_36617_42043# VSS 3.11fF
C18862 a_34611_42089# VSS 0.31fF
C18863 a_31976_41831# VSS 0.49fF
C18864 a_30523_41245# VSS 1.44fF
C18865 a_33309_41479# VSS 1.65fF
C18866 a_33489_42043# VSS 3.06fF
C18867 a_32035_42089# VSS 0.32fF
C18868 a_28940_41831# VSS 0.46fF
C18869 a_29217_41570# VSS 1.59fF
C18870 a_30913_42043# VSS 3.04fF
C18871 a_28999_42089# VSS 0.32fF
C18872 a_26272_41831# VSS 0.45fF
C18873 a_27421_41814# VSS 1.76fF
C18874 a_29036_41831# VSS 1.63fF
C18875 a_27877_42043# VSS 3.06fF
C18876 a_26331_42089# VSS 0.32fF
C18877 a_21981_34191# VSS 1.66fF
C18878 a_10767_39087# VSS 1.14fF
C18879 a_25209_42043# VSS 2.99fF
C18880 a_12116_39783# VSS 0.88fF
C18881 a_20337_41831# VSS 0.43fF
C18882 a_17900_41831# VSS 0.45fF
C18883 a_20572_40517# VSS 1.64fF
C18884 a_20645_42044# VSS 3.00fF
C18885 a_14149_39747# VSS 2.56fF
C18886 a_17959_42089# VSS 0.32fF
C18887 a_15324_41831# VSS 0.45fF
C18888 a_16837_42043# VSS 3.03fF
C18889 a_15383_42089# VSS 0.31fF
C18890 a_15420_41831# VSS 1.36fF
C18891 a_14261_42043# VSS 2.93fF
C18892 a_10677_41831# VSS 0.48fF
C18893 a_11921_41814# VSS 1.36fF
C18894 a_10591_42089# VSS 0.32fF
C18895 a_10985_42044# VSS 3.02fF
C18896 a_10651_42035# VSS 1.42fF
C18897 a_39079_40947# VSS 1.59fF
C18898 a_38927_42359# VSS 0.31fF
C18899 a_37923_42359# VSS 0.31fF
C18900 a_39013_42693# VSS 0.44fF
C18901 a_39321_42333# VSS 2.87fF
C18902 a_38737_41814# VSS 1.44fF
C18903 a_37864_42693# VSS 0.44fF
C18904 a_36801_42405# VSS 2.96fF
C18905 a_33223_42359# VSS 0.32fF
C18906 a_33309_42693# VSS 0.48fF
C18907 a_33617_42333# VSS 2.94fF
C18908 a_31923_42367# VSS 0.52fF
C18909 a_12116_40871# VSS 2.69fF
C18910 a_27947_41245# VSS 1.67fF
C18911 a_27519_42359# VSS 0.34fF
C18912 a_27605_42693# VSS 0.47fF
C18913 a_27913_42333# VSS 2.94fF
C18914 a_25319_42359# VSS 0.31fF
C18915 a_25260_42693# VSS 0.48fF
C18916 a_10873_40693# VSS 2.69fF
C18917 a_11041_40948# VSS 3.00fF
C18918 a_24937_41479# VSS 1.42fF
C18919 a_24197_42405# VSS 2.79fF
C18920 a_23741_42567# VSS 1.31fF
C18921 a_20752_42693# VSS 0.47fF
C18922 a_18235_42359# VSS 0.31fF
C18923 a_21815_42351# VSS 0.37fF
C18924 a_19689_42405# VSS 3.03fF
C18925 a_18176_42693# VSS 0.44fF
C18926 a_18272_42693# VSS 1.50fF
C18927 a_17113_42405# VSS 2.92fF
C18928 a_14497_42658# VSS 1.57fF
C18929 a_13167_42359# VSS 0.31fF
C18930 a_13253_42693# VSS 0.47fF
C18931 a_13561_42333# VSS 2.88fF
C18932 a_13227_42333# VSS 1.39fF
C18933 a_6369_39465# VSS 0.48fF
C18934 a_6619_41909# VSS 0.36fF
C18935 a_5558_41935# VSS 0.30fF
C18936 a_4984_41935# VSS 0.37fF
C18937 a_4432_42313# VSS 0.36fF
C18938 a_4149_41941# VSS 0.34fF
C18939 a_3983_41941# VSS 0.50fF
C18940 cgen.dlycontrol2_in[3] VSS 1.33fF
C18941 a_10949_42364# VSS 0.41fF
C18942 a_11021_42619# VSS 0.56fF
C18943 a_10781_42364# VSS 2.82fF
C18944 a_40256_42919# VSS 0.49fF
C18945 a_44774_40821# VSS 1.08fF
C18946 a_40315_43177# VSS 0.31fF
C18947 a_37680_42919# VSS 0.49fF
C18948 a_37960_42693# VSS 1.48fF
C18949 a_39193_43131# VSS 2.90fF
C18950 a_37739_43177# VSS 0.33fF
C18951 a_34552_42919# VSS 0.44fF
C18952 a_36345_42567# VSS 1.73fF
C18953 a_36617_43131# VSS 3.08fF
C18954 a_34611_43177# VSS 0.30fF
C18955 a_31976_42919# VSS 0.44fF
C18956 a_34553_42658# VSS 1.55fF
C18957 a_33489_43131# VSS 2.99fF
C18958 a_32035_43177# VSS 0.30fF
C18959 a_28848_42919# VSS 0.49fF
C18960 a_32072_42919# VSS 1.38fF
C18961 a_30913_43131# VSS 2.86fF
C18962 a_28907_43177# VSS 0.32fF
C18963 a_27329_42902# VSS 1.61fF
C18964 a_27785_43131# VSS 3.05fF
C18965 a_24753_42919# VSS 0.43fF
C18966 a_23604_42919# VSS 0.43fF
C18967 a_25997_42902# VSS 1.49fF
C18968 a_21028_42919# VSS 0.44fF
C18969 a_25061_43132# VSS 2.87fF
C18970 a_11389_40443# VSS 1.97fF
C18971 a_23700_42919# VSS 1.57fF
C18972 a_22541_43131# VSS 2.88fF
C18973 a_21087_43177# VSS 0.30fF
C18974 a_19965_43131# VSS 2.87fF
C18975 a_16381_42919# VSS 0.47fF
C18976 a_17625_42902# VSS 1.38fF
C18977 a_16689_43132# VSS 2.88fF
C18978 a_16355_43123# VSS 1.48fF
C18979 a_13805_42919# VSS 0.46fF
C18980 a_15049_42902# VSS 1.72fF
C18981 a_14113_43132# VSS 2.91fF
C18982 a_12658_42895# VSS 1.11fF
C18983 a_7263_42453# VSS 0.47fF
C18984 a_6007_42479# VSS 0.42fF
C18985 a_4253_42729# VSS 0.41fF
C18986 cgen.dlycontrol2_in[4] VSS 2.27fF
C18987 a_11021_43011# VSS 1.12fF
C18988 a_10949_43124# VSS 1.39fF
C18989 a_11910_43047# VSS 0.38fF
C18990 a_44739_43567# VSS 0.46fF
C18991 a_40532_43781# VSS 0.44fF
C18992 a_40349_40726# VSS 1.59fF
C18993 a_39469_43493# VSS 2.84fF
C18994 a_39013_43655# VSS 1.90fF
C18995 a_30543_40721# VSS 1.51fF
C18996 a_35656_43781# VSS 0.44fF
C18997 a_35752_43781# VSS 1.66fF
C18998 a_34593_43493# VSS 2.85fF
C18999 a_33283_42333# VSS 1.30fF
C19000 a_24833_40719# VSS 1.29fF
C19001 a_31095_42367# VSS 0.39fF
C19002 a_30044_43781# VSS 0.46fF
C19003 a_26515_43447# VSS 0.30fF
C19004 a_30140_43781# VSS 1.23fF
C19005 a_28981_43493# VSS 2.94fF
C19006 a_28525_43655# VSS 1.35fF
C19007 a_20438_35431# VSS 0.92fF
C19008 a_26456_43781# VSS 0.44fF
C19009 a_11497_40719# VSS 3.84fF
C19010 a_25393_43493# VSS 2.82fF
C19011 a_23420_43781# VSS 0.45fF
C19012 a_22361_41479# VSS 1.32fF
C19013 a_22357_43493# VSS 2.91fF
C19014 a_20848_41605# VSS 1.57fF
C19015 a_12228_40693# VSS 1.69fF
C19016 a_20016_43781# VSS 0.48fF
C19017 cgen.start_conv_in VSS 5.64fF
C19018 a_19233_41479# VSS 1.67fF
C19019 a_18953_43493# VSS 2.96fF
C19020 a_17996_41831# VSS 1.38fF
C19021 a_17902_43439# VSS 0.41fF
C19022 a_15921_38550# VSS 1.25fF
C19023 a_13443_43447# VSS 0.31fF
C19024 a_13529_43781# VSS 0.48fF
C19025 a_17154_43671# VSS 0.50fF
C19026 a_12069_38517# VSS 2.61fF
C19027 a_12237_38772# VSS 0.68fF
C19028 a_13837_43421# VSS 2.91fF
C19029 a_13503_43421# VSS 1.44fF
C19030 a_10867_43447# VSS 0.31fF
C19031 a_6311_42692# VSS 0.32fF
C19032 a_6554_43255# VSS 0.33fF
C19033 a_2021_26677# VSS 2.02fF
C19034 a_3879_42997# VSS 0.51fF
C19035 a_2847_43327# VSS 0.38fF
C19036 a_1591_43029# VSS 0.51fF
C19037 a_1586_33927# VSS 2.98fF
C19038 cgen.dlycontrol4_in[2] VSS 5.14fF
C19039 a_10953_43781# VSS 0.47fF
C19040 a_11261_43421# VSS 2.88fF
C19041 cgen.dlycontrol4_in[1] VSS 4.51fF
C19042 a_34552_44007# VSS 0.48fF
C19043 a_44733_44431# VSS 0.34fF
C19044 a_30819_40191# VSS 0.74fF
C19045 a_33395_43455# VSS 1.31fF
C19046 a_34611_44265# VSS 0.32fF
C19047 a_31976_44007# VSS 0.48fF
C19048 a_11113_39747# VSS 1.71fF
C19049 a_33489_44219# VSS 2.95fF
C19050 a_32035_44265# VSS 0.33fF
C19051 a_28572_44007# VSS 0.49fF
C19052 a_30913_44219# VSS 2.90fF
C19053 a_29627_43983# VSS 0.84fF
C19054 a_28631_44265# VSS 0.32fF
C19055 a_26552_43781# VSS 1.45fF
C19056 cgen.dlycontrol4_in[0] VSS 13.41fF
C19057 a_27509_44219# VSS 3.15fF
C19058 a_12197_43746# VSS 1.56fF
C19059 a_23512_44007# VSS 0.48fF
C19060 a_14773_43746# VSS 1.76fF
C19061 a_23571_44265# VSS 0.30fF
C19062 a_20936_44007# VSS 0.44fF
C19063 a_21124_42919# VSS 1.40fF
C19064 a_10873_39605# VSS 2.37fF
C19065 a_11041_39860# VSS 4.29fF
C19066 a_11149_40188# VSS 6.13fF
C19067 a_11317_40188# VSS 2.88fF
C19068 a_22085_42902# VSS 2.15fF
C19069 a_22449_44219# VSS 2.89fF
C19070 a_20995_44265# VSS 0.30fF
C19071 a_17900_44007# VSS 0.45fF
C19072 a_19873_44219# VSS 2.92fF
C19073 a_17959_44265# VSS 0.32fF
C19074 a_15324_44007# VSS 0.44fF
C19075 a_16837_44219# VSS 2.88fF
C19076 a_15383_44265# VSS 0.30fF
C19077 a_15420_44007# VSS 1.46fF
C19078 a_14261_44219# VSS 2.86fF
C19079 a_10677_44007# VSS 0.43fF
C19080 a_3983_43567# VSS 0.47fF
C19081 a_2867_43541# VSS 0.45fF
C19082 a_1927_43541# VSS 0.45fF
C19083 a_10927_43421# VSS 1.56fF
C19084 a_10985_44220# VSS 2.80fF
C19085 a_10781_42869# VSS 3.16fF
C19086 a_32219_44535# VSS 0.31fF
C19087 a_32160_44869# VSS 0.44fF
C19088 a_29367_44535# VSS 0.30fF
C19089 a_37731_44527# VSS 0.50fF
C19090 a_36854_44527# VSS 0.31fF
C19091 a_35290_44527# VSS 0.49fF
C19092 a_34002_44527# VSS 0.40fF
C19093 a_31978_43439# VSS 0.78fF
C19094 a_32256_44869# VSS 1.49fF
C19095 a_31097_44581# VSS 3.15fF
C19096 a_30641_44743# VSS 2.42fF
C19097 a_29308_44869# VSS 0.44fF
C19098 a_26331_44535# VSS 0.32fF
C19099 a_29404_44869# VSS 1.44fF
C19100 a_28245_44581# VSS 3.03fF
C19101 a_27789_44743# VSS 1.92fF
C19102 a_26272_44869# VSS 0.48fF
C19103 a_24937_43655# VSS 1.40fF
C19104 a_25209_44581# VSS 3.03fF
C19105 a_23604_44869# VSS 0.43fF
C19106 a_20811_44535# VSS 0.31fF
C19107 a_23700_44869# VSS 1.73fF
C19108 a_22541_44581# VSS 3.07fF
C19109 a_21032_44007# VSS 1.64fF
C19110 a_20752_44869# VSS 0.47fF
C19111 a_17867_44535# VSS 0.32fF
C19112 a_19417_43990# VSS 2.28fF
C19113 a_19689_44581# VSS 3.03fF
C19114 a_17996_44007# VSS 1.83fF
C19115 a_17808_44869# VSS 0.48fF
C19116 a_15107_44535# VSS 0.31fF
C19117 a_16657_42567# VSS 2.29fF
C19118 a_16745_44581# VSS 3.08fF
C19119 a_13779_43123# VSS 1.41fF
C19120 a_15048_44869# VSS 0.47fF
C19121 a_13805_43990# VSS 2.32fF
C19122 a_13985_44581# VSS 3.08fF
C19123 a_12196_44869# VSS 0.43fF
C19124 cgen.dlycontrol4_in[3] VSS 6.73fF
C19125 a_3325_43023# VSS 0.88fF
C19126 cgen.dlycontrol4_in[4] VSS 5.28fF
C19127 a_12292_44869# VSS 1.74fF
C19128 a_11133_44581# VSS 2.99fF
C19129 a_10651_44211# VSS 1.51fF
C19130 a_5747_44655# VSS 0.33fF
C19131 a_44966_43255# VSS 1.35fF
C19132 a_45064_44807# VSS 0.30fF
C19133 a_6800_44629# VSS 0.35fF
C19134 cgen.dlycontrol3_in[0] VSS 2.17fF
C19135 a_6141_44629# VSS 0.84fF
C19136 a_4257_34319# VSS 2.00fF
C19137 a_2659_35015# VSS 3.83fF
C19138 a_47026_45519# VSS 0.31fF
C19139 a_43720_32143# VSS 1.88fF
C19140 cgen.dlycontrol4_in[5] VSS 3.67fF
C19141 a_5921_44629# VSS 0.37fF
C19142 a_2939_45503# VSS 0.68fF
C19143 a_1683_45205# VSS 0.50fF
C19144 a_44635_46025# VSS 0.40fF
C19145 a_46968_45743# VSS 0.55fF
C19146 a_47290_45717# VSS 0.63fF
C19147 a_47147_44655# VSS 0.45fF
C19148 a_4313_44111# VSS 0.47fF
C19149 dummypin[7] VSS 0.69fF
C19150 adc_top_88.HI VSS 0.34fF
C19151 nmat.col[31] VSS 12.10fF
C19152 a_46027_44905# VSS 0.76fF
C19153 a_7109_29423# VSS 10.00fF
C19154 a_40741_46565# VSS 0.35fF
C19155 a_40467_46261# VSS 0.37fF
C19156 nmat.rowon_n[14] VSS 8.37fF
C19157 a_13091_18535# VSS 2.68fF
C19158 a_16926_46261# VSS 0.42fF
C19159 a_14427_46519# VSS 0.32fF
C19160 a_1987_45370# VSS 0.34fF
C19161 a_2559_46261# VSS 0.31fF
C19162 a_40837_46261# VSS 11.06fF
C19163 a_47975_46831# VSS 0.40fF
C19164 a_36532_46805# VSS 0.92fF
C19165 a_42024_46805# VSS 0.65fF
C19166 a_41926_46983# VSS 0.56fF
C19167 a_37519_46983# VSS 0.33fF
C19168 a_35068_46805# VSS 0.32fF
C19169 a_32827_46805# VSS 0.54fF
C19170 a_1781_9308# VSS 13.20fF
C19171 a_27411_46805# VSS 0.68fF
C19172 a_26155_46831# VSS 0.46fF
C19173 a_25681_46831# VSS 0.61fF
C19174 a_18869_46831# VSS 0.42fF
C19175 a_12079_9615# VSS 6.82fF
C19176 a_13091_7655# VSS 5.03fF
C19177 a_14379_46287# VSS 0.40fF
C19178 a_25189_46287# VSS 0.40fF
C19179 a_21797_47081# VSS 0.31fF
C19180 a_21837_46983# VSS 0.38fF
C19181 nmat.rowon_n[12] VSS 10.49fF
C19182 a_18521_46837# VSS 0.34fF
C19183 a_17478_46805# VSS 0.40fF
C19184 a_16552_46805# VSS 0.40fF
C19185 a_6747_46831# VSS 1.01fF
C19186 cgen.dlycontrol3_in[1] VSS 3.03fF
C19187 a_11823_46973# VSS 0.53fF
C19188 a_11071_46805# VSS 0.66fF
C19189 a_6830_44655# VSS 0.57fF
C19190 a_4955_40277# VSS 2.42fF
C19191 a_5455_46831# VSS 0.50fF
C19192 a_5173_45993# VSS 0.31fF
C19193 a_5221_45199# VSS 0.44fF
C19194 a_4979_38127# VSS 0.85fF
C19195 a_29937_31055# VSS 5.26fF
C19196 a_45112_47607# VSS 0.74fF
C19197 a_44976_47349# VSS 0.42fF
C19198 a_40105_47375# VSS 3.12fF
C19199 a_39647_47679# VSS 0.60fF
C19200 a_38569_46831# VSS 0.32fF
C19201 a_38391_47381# VSS 0.43fF
C19202 a_35186_47375# VSS 3.51fF
C19203 a_34850_47695# VSS 0.71fF
C19204 a_33986_47695# VSS 0.49fF
C19205 a_33986_47375# VSS 0.41fF
C19206 a_31105_46805# VSS 0.51fF
C19207 a_32371_47349# VSS 0.32fF
C19208 a_31675_47695# VSS 8.87fF
C19209 a_29711_47679# VSS 0.68fF
C19210 a_28639_47081# VSS 0.30fF
C19211 a_28455_47381# VSS 0.43fF
C19212 a_23823_47679# VSS 0.65fF
C19213 a_22567_47381# VSS 0.45fF
C19214 a_20316_47607# VSS 0.32fF
C19215 a_19441_47491# VSS 0.32fF
C19216 a_18660_47607# VSS 0.33fF
C19217 a_18083_47593# VSS 0.63fF
C19218 a_17927_47349# VSS 0.32fF
C19219 a_14379_6567# VSS 5.11fF
C19220 a_17012_47349# VSS 0.39fF
C19221 a_12604_47080# VSS 0.87fF
C19222 a_9839_47679# VSS 0.41fF
C19223 a_8453_46287# VSS 0.39fF
C19224 a_8583_47381# VSS 0.49fF
C19225 a_5566_44905# VSS 0.34fF
C19226 a_3987_47375# VSS 0.36fF
C19227 a_3793_47479# VSS 0.31fF
C19228 a_1775_47375# VSS 0.62fF
C19229 a_45201_47919# VSS 0.36fF
C19230 a_36956_47919# VSS 0.50fF
C19231 a_35730_47919# VSS 0.72fF
C19232 a_32687_46607# VSS 6.59fF
C19233 a_31767_47919# VSS 0.39fF
C19234 a_25466_47919# VSS 0.72fF
C19235 a_24602_47919# VSS 0.49fF
C19236 a_43267_47081# VSS 0.55fF
C19237 a_13643_29415# VSS 2.86fF
C19238 a_47407_47919# VSS 0.46fF
C19239 a_46487_47919# VSS 0.43fF
C19240 a_41663_47893# VSS 0.47fF
C19241 a_40047_47919# VSS 0.43fF
C19242 a_35786_47893# VSS 0.44fF
C19243 a_31152_48071# VSS 0.62fF
C19244 a_30999_48071# VSS 1.43fF
C19245 a_24602_48169# VSS 0.50fF
C19246 a_15899_47939# VSS 1.84fF
C19247 a_19541_28879# VSS 3.94fF
C19248 a_22895_47893# VSS 0.31fF
C19249 a_20879_47893# VSS 0.44fF
C19250 a_19647_48052# VSS 0.34fF
C19251 a_19491_47893# VSS 0.33fF
C19252 a_3983_47919# VSS 0.33fF
C19253 a_8079_46519# VSS 0.80fF
C19254 a_4579_47919# VSS 1.76fF
C19255 a_11547_48061# VSS 0.40fF
C19256 a_10795_47893# VSS 0.64fF
C19257 a_2935_38279# VSS 2.76fF
C19258 a_4128_46983# VSS 1.66fF
C19259 a_3978_48071# VSS 0.65fF
C19260 a_44697_48783# VSS 1.20fF
C19261 a_43315_48437# VSS 2.01fF
C19262 a_33423_47695# VSS 8.04fF
C19263 a_33839_46805# VSS 1.57fF
C19264 a_40949_48437# VSS 0.42fF
C19265 a_39647_48767# VSS 0.37fF
C19266 a_38391_48469# VSS 0.46fF
C19267 a_14887_46377# VSS 6.67fF
C19268 a_29076_48695# VSS 1.68fF
C19269 a_28901_48437# VSS 0.54fF
C19270 a_28629_48437# VSS 0.49fF
C19271 a_21063_48723# VSS 0.37fF
C19272 a_19399_48437# VSS 0.31fF
C19273 a_17397_48463# VSS 0.66fF
C19274 a_17927_48437# VSS 0.31fF
C19275 a_17049_48579# VSS 0.30fF
C19276 a_13688_47893# VSS 0.57fF
C19277 a_11067_30287# VSS 12.96fF
C19278 a_13275_48783# VSS 6.31fF
C19279 a_9871_48463# VSS 0.43fF
C19280 a_5411_48695# VSS 0.52fF
C19281 a_4167_48463# VSS 0.45fF
C19282 a_1769_14735# VSS 6.96fF
C19283 a_1739_47893# VSS 2.96fF
C19284 cgen.dlycontrol3_in[3] VSS 2.92fF
C19285 cgen.dlycontrol3_in[2] VSS 3.40fF
C19286 a_30111_47911# VSS 4.46fF
C19287 a_38695_48634# VSS 0.69fF
C19288 a_6283_31591# VSS 14.62fF
C19289 a_27020_49007# VSS 0.49fF
C19290 a_25794_49007# VSS 0.70fF
C19291 a_21279_48999# VSS 1.52fF
C19292 nmat.col[15] VSS 9.20fF
C19293 a_21215_48071# VSS 2.20fF
C19294 a_7578_48553# VSS 0.41fF
C19295 a_4263_49007# VSS 0.49fF
C19296 a_47591_49007# VSS 0.44fF
C19297 a_45450_48695# VSS 0.90fF
C19298 a_45370_48169# VSS 0.42fF
C19299 a_44774_48695# VSS 0.45fF
C19300 a_44870_48437# VSS 0.59fF
C19301 a_38793_49007# VSS 0.34fF
C19302 a_33467_46261# VSS 4.88fF
C19303 a_33957_48437# VSS 0.76fF
C19304 a_36265_48981# VSS 0.44fF
C19305 a_32871_49007# VSS 0.52fF
C19306 a_25850_48981# VSS 0.40fF
C19307 a_23971_49140# VSS 0.48fF
C19308 a_21923_47919# VSS 0.38fF
C19309 a_21883_48981# VSS 0.33fF
C19310 a_19487_49159# VSS 0.31fF
C19311 a_18359_49140# VSS 0.88fF
C19312 a_18203_48981# VSS 0.34fF
C19313 a_16219_49007# VSS 0.44fF
C19314 a_6467_29415# VSS 6.16fF
C19315 a_9135_49257# VSS 0.34fF
C19316 a_8907_48437# VSS 1.22fF
C19317 a_8267_49159# VSS 0.68fF
C19318 a_6895_48981# VSS 0.40fF
C19319 a_5639_49007# VSS 0.42fF
C19320 a_4075_49007# VSS 0.46fF
C19321 a_46487_49871# VSS 0.48fF
C19322 a_41731_49525# VSS 7.32fF
C19323 a_37820_30485# VSS 5.19fF
C19324 a_40415_49551# VSS 0.41fF
C19325 a_37471_49551# VSS 0.52fF
C19326 a_33281_49551# VSS 0.67fF
C19327 a_32411_49559# VSS 0.31fF
C19328 pmat.col[11] VSS 6.41fF
C19329 a_9411_2215# VSS 12.22fF
C19330 a_25802_48169# VSS 0.95fF
C19331 a_25839_49783# VSS 1.42fF
C19332 a_24270_49783# VSS 0.30fF
C19333 a_20619_49551# VSS 0.52fF
C19334 a_18947_49811# VSS 0.49fF
C19335 a_15839_49525# VSS 0.44fF
C19336 nmat.sw VSS 18.78fF
C19337 a_11948_49783# VSS 1.39fF
C19338 dummypin[6] VSS 0.88fF
C19339 adc_top_87.HI VSS 0.37fF
C19340 pmat.col[23] VSS 6.32fF
C19341 pmat.col[15] VSS 6.63fF
C19342 pmat.col[8] VSS 6.33fF
C19343 a_19283_49783# VSS 2.63fF
C19344 a_22499_49783# VSS 3.15fF
C19345 a_20475_49783# VSS 1.49fF
C19346 a_12044_49641# VSS 0.60fF
C19347 a_11067_49871# VSS 6.45fF
C19348 a_47211_50069# VSS 0.54fF
C19349 a_46211_50095# VSS 0.41fF
C19350 a_38851_28327# VSS 6.73fF
C19351 a_25695_28111# VSS 8.63fF
C19352 a_10883_3303# VSS 15.32fF
C19353 a_34948_50069# VSS 0.34fF
C19354 a_24775_50095# VSS 0.42fF
C19355 a_21371_50087# VSS 4.83fF
C19356 a_23971_50228# VSS 0.38fF
C19357 a_18487_50069# VSS 0.54fF
C19358 a_15747_50069# VSS 0.38fF
C19359 a_14287_50345# VSS 0.35fF
C19360 a_14249_49525# VSS 0.48fF
C19361 a_7373_49007# VSS 0.68fF
C19362 a_11803_49551# VSS 0.63fF
C19363 a_11455_50237# VSS 0.43fF
C19364 a_10703_50069# VSS 0.64fF
C19365 a_4627_50095# VSS 0.41fF
C19366 a_2847_50069# VSS 0.48fF
C19367 a_1895_50308# VSS 0.45fF
C19368 a_1591_50095# VSS 0.50fF
C19369 pmat.col[26] VSS 6.28fF
C19370 pmat.col[21] VSS 6.17fF
C19371 _1183_.A2 VSS 20.98fF
C19372 a_25879_31591# VSS 9.26fF
C19373 pmat.col[16] VSS 6.15fF
C19374 a_35224_50613# VSS 0.32fF
C19375 a_30663_50087# VSS 10.83fF
C19376 a_22199_30287# VSS 5.50fF
C19377 a_28131_50069# VSS 1.26fF
C19378 a_28049_50613# VSS 0.33fF
C19379 pmat.col[5] VSS 6.73fF
C19380 a_22343_50613# VSS 0.32fF
C19381 a_21395_50857# VSS 1.04fF
C19382 a_17163_50857# VSS 0.59fF
C19383 a_15655_50613# VSS 0.41fF
C19384 a_11711_50959# VSS 5.76fF
C19385 a_4075_31591# VSS 8.06fF
C19386 a_4927_50613# VSS 0.52fF
C19387 cgen.dlycontrol3_in[4] VSS 1.65fF
C19388 pmat.col[29] VSS 6.29fF
C19389 a_26891_28327# VSS 8.78fF
C19390 a_30571_50959# VSS 10.64fF
C19391 pmat.col[19] VSS 6.20fF
C19392 a_28915_50959# VSS 6.08fF
C19393 pmat.col[10] VSS 6.15fF
C19394 pmat.col[7] VSS 6.16fF
C19395 a_38575_50639# VSS 0.36fF
C19396 a_17139_30503# VSS 8.09fF
C19397 a_21647_51183# VSS 0.47fF
C19398 a_20411_51157# VSS 0.34fF
C19399 a_19675_51157# VSS 0.36fF
C19400 a_18429_51189# VSS 0.34fF
C19401 a_17033_51183# VSS 0.46fF
C19402 a_17559_51157# VSS 0.34fF
C19403 a_1769_13103# VSS 3.94fF
C19404 a_9319_50639# VSS 0.30fF
C19405 a_13091_50095# VSS 0.37fF
C19406 a_12559_51325# VSS 0.44fF
C19407 a_11807_51157# VSS 0.60fF
C19408 a_10205_51433# VSS 0.31fF
C19409 a_9184_51335# VSS 0.33fF
C19410 a_2983_48071# VSS 2.04fF
C19411 a_4399_51157# VSS 1.30fF
C19412 pmat.col[28] VSS 6.32fF
C19413 a_15667_27239# VSS 10.96fF
C19414 pmat.col[24] VSS 6.22fF
C19415 pmat.col[17] VSS 6.05fF
C19416 pmat.col[14] VSS 6.31fF
C19417 pmat.col[12] VSS 6.62fF
C19418 pmat.col[0] VSS 6.99fF
C19419 a_31631_51701# VSS 0.30fF
C19420 a_24407_31375# VSS 11.15fF
C19421 a_21739_29415# VSS 13.95fF
C19422 a_18823_50247# VSS 1.48fF
C19423 a_20776_51959# VSS 0.33fF
C19424 a_19948_51959# VSS 0.32fF
C19425 a_18547_51565# VSS 3.63fF
C19426 a_16083_50069# VSS 3.47fF
C19427 a_18568_51959# VSS 0.33fF
C19428 a_14825_50095# VSS 0.35fF
C19429 a_14491_51969# VSS 0.40fF
C19430 a_13739_51701# VSS 0.66fF
C19431 a_12263_50959# VSS 12.66fF
C19432 a_9427_50095# VSS 0.86fF
C19433 a_9463_50877# VSS 1.10fF
C19434 a_9335_51727# VSS 0.35fF
C19435 a_9919_51959# VSS 0.44fF
C19436 a_7907_52031# VSS 0.38fF
C19437 a_6651_51733# VSS 0.38fF
C19438 a_2389_45859# VSS 3.26fF
C19439 a_4403_51701# VSS 0.33fF
C19440 a_2715_51969# VSS 0.44fF
C19441 a_2195_51701# VSS 0.39fF
C19442 pmat.col[27] VSS 6.27fF
C19443 pmat.col[22] VSS 6.20fF
C19444 pmat.col[20] VSS 6.22fF
C19445 pmat.col[18] VSS 6.29fF
C19446 pmat.col[13] VSS 6.20fF
C19447 pmat.col[1] VSS 8.29fF
C19448 pmat.col[9] VSS 6.27fF
C19449 pmat.col[6] VSS 6.16fF
C19450 a_5363_33551# VSS 8.43fF
C19451 pmat.col[3] VSS 6.18fF
C19452 pmat.col[4] VSS 6.27fF
C19453 pmat.col[2] VSS 6.20fF
C19454 a_19584_52423# VSS 1.42fF
C19455 a_16800_47213# VSS 1.30fF
C19456 a_47449_52271# VSS 0.59fF
C19457 a_37709_52245# VSS 0.30fF
C19458 a_34942_51701# VSS 1.27fF
C19459 a_34705_51959# VSS 3.25fF
C19460 _1184_.A2 VSS 14.90fF
C19461 a_16311_28327# VSS 17.95fF
C19462 ANTENNA__1195__A1.DIODE VSS 21.62fF
C19463 ANTENNA__1395__B1.DIODE VSS 18.48fF
C19464 a_13459_28111# VSS 17.35fF
C19465 ANTENNA__1196__A2.DIODE VSS 19.18fF
C19466 a_19488_52423# VSS 0.32fF
C19467 a_10245_51335# VSS 0.54fF
C19468 a_8385_51727# VSS 1.56fF
C19469 a_5785_48463# VSS 0.57fF
C19470 cgen.enable_dlycontrol_in VSS 7.52fF
C19471 pmat.col[30] VSS 6.21fF
C19472 pmat.col[25] VSS 6.45fF
C19473 a_13091_28327# VSS 19.11fF
C19474 a_18243_28327# VSS 10.19fF
C19475 _1192_.A2 VSS 21.10fF
C19476 _1192_.B1 VSS 27.46fF
C19477 _1194_.B1 VSS 25.93fF
C19478 ANTENNA__1395__A2.DIODE VSS 12.60fF
C19479 a_11067_27239# VSS 12.11fF
C19480 nmat.en_bit_n[1] VSS 5.59fF
C19481 a_24591_28327# VSS 9.47fF
C19482 ANTENNA__1197__B.DIODE VSS 15.96fF
C19483 ANTENNA__1184__B1.DIODE VSS 17.11fF
C19484 ANTENNA__1187__B1.DIODE VSS 13.01fF
C19485 a_24867_53135# VSS 9.26fF
C19486 _1187_.A2 VSS 31.48fF
C19487 a_23395_53135# VSS 5.25fF
C19488 ANTENNA__1190__A1.DIODE VSS 28.03fF
C19489 ANTENNA__1190__B1.DIODE VSS 19.06fF
C19490 a_20583_53080# VSS 0.38fF
C19491 pmat.rowoff_n[2] VSS 2.04fF
C19492 pmat.rowoff_n[1] VSS 3.29fF
C19493 pmat.rowoff_n[3] VSS 1.32fF
C19494 a_19579_52789# VSS 0.33fF
C19495 a_18777_51183# VSS 0.30fF
C19496 a_18199_52789# VSS 0.55fF
C19497 a_16113_52271# VSS 0.37fF
C19498 ANTENNA__1395__A1.DIODE VSS 13.92fF
C19499 _1194_.A2 VSS 26.69fF
C19500 ANTENNA__1197__A.DIODE VSS 19.79fF
C19501 a_13091_52047# VSS 5.40fF
C19502 a_5123_52423# VSS 1.11fF
C19503 a_2315_44124# VSS 2.77fF
C19504 a_2163_53057# VSS 0.50fF
C19505 a_1643_52789# VSS 0.38fF
C19506 pmat.col[31] VSS 13.28fF
C19507 a_14653_53458# VSS 2.17fF
C19508 a_9827_53379# VSS 0.71fF
C19509 a_4123_52789# VSS 0.46fF
C19510 a_2944_52789# VSS 0.45fF
C19511 _1519_.A VSS 13.89fF
C19512 a_12213_53359# VSS 0.61fF
C19513 a_9463_53511# VSS 0.76fF
C19514 a_10641_52815# VSS 0.95fF
C19515 a_9367_53511# VSS 0.31fF
C19516 a_7163_53333# VSS 0.46fF
C19517 _1196_.B1 VSS 31.09fF
C19518 a_12003_52815# VSS 0.92fF
C19519 a_9871_53903# VSS 0.33fF
C19520 a_8735_54207# VSS 0.44fF
C19521 a_7479_53909# VSS 0.41fF
C19522 a_6559_53903# VSS 0.42fF
C19523 a_6553_53047# VSS 0.98fF
C19524 a_4259_31375# VSS 6.57fF
C19525 a_3707_53903# VSS 0.55fF
C19526 a_1591_52815# VSS 1.05fF
C19527 _1179_.X VSS 20.08fF
C19528 a_82787_54421# VSS 0.57fF
C19529 ANTENNA_fanout52_A.DIODE VSS 13.08fF
C19530 a_82815_54965# VSS 0.43fF
C19531 dummypin[5] VSS 0.86fF
C19532 adc_top_86.HI VSS 0.34fF
C19533 a_3199_53877# VSS 0.61fF
C19534 a_12895_53359# VSS 0.39fF
C19535 a_9213_53903# VSS 0.85fF
C19536 a_51202_55126# VSS 0.37fF
C19537 inp_analog VSS 5.29fF
C19538 a_36234_55126# VSS 0.40fF
C19539 pmat.en_bit_n[0] VSS 4.75fF
C19540 a_35230_55126# VSS 0.39fF
C19541 pmat.en_bit_n[2] VSS 5.65fF
C19542 a_34226_55126# VSS 0.39fF
C19543 pmat.en_bit_n[1] VSS 1.15fF
C19544 a_20170_55126# VSS 0.41fF
C19545 pmat.en_C0_n VSS 1.17fF
C19546 a_18162_55166# VSS 6.70fF
C19547 a_18546_55168# VSS 4.48fF
C19548 pmat.sw VSS 17.71fF
C19549 a_14163_55295# VSS 0.40fF
C19550 a_12907_54997# VSS 0.42fF
C19551 a_4587_53505# VSS 0.51fF
C19552 a_5329_54965# VSS 0.35fF
C19553 a_4243_54991# VSS 0.39fF
C19554 a_3970_55311# VSS 0.35fF
C19555 a_2163_55233# VSS 0.54fF
C19556 a_1643_54965# VSS 0.39fF
C19557 a_1586_50247# VSS 7.40fF
C19558 a_6559_33767# VSS 6.92fF
C19559 a_5955_55223# VSS 0.58fF
C19560 a_10497_54697# VSS 0.97fF
C19561 a_10955_55687# VSS 0.50fF
C19562 a_10409_53903# VSS 0.61fF
C19563 a_2787_55535# VSS 0.55fF
C19564 a_1591_54991# VSS 0.83fF
C19565 a_2840_55509# VSS 0.32fF
C19566 a_18162_56170# VSS 5.02fF
C19567 a_18546_56172# VSS 3.53fF
C19568 pmat.rowoff_n[0] VSS 1.28fF
C19569 pmat.row_n[0] VSS 14.33fF
C19570 a_11711_56079# VSS 0.55fF
C19571 a_11202_55687# VSS 0.85fF
C19572 a_10595_53361# VSS 0.68fF
C19573 a_11444_55535# VSS 0.36fF
C19574 a_9581_56079# VSS 1.90fF
C19575 a_9103_56383# VSS 0.54fF
C19576 a_8013_56085# VSS 0.32fF
C19577 a_7847_56085# VSS 0.53fF
C19578 a_5245_56053# VSS 0.33fF
C19579 a_3967_56311# VSS 0.37fF
C19580 a_1644_56053# VSS 0.31fF
C19581 pmat.rowon_n[0] VSS 11.46fF
C19582 a_2411_43301# VSS 12.47fF
C19583 a_11902_56775# VSS 0.65fF
C19584 a_18162_57174# VSS 4.96fF
C19585 pmat.rowon_n[1] VSS 4.15fF
C19586 a_18546_57176# VSS 3.50fF
C19587 a_4535_56623# VSS 0.33fF
C19588 a_2163_56765# VSS 0.55fF
C19589 a_1643_56597# VSS 0.39fF
C19590 a_12613_57141# VSS 0.61fF
C19591 a_8507_57487# VSS 0.32fF
C19592 a_8749_57141# VSS 0.92fF
C19593 a_8477_57141# VSS 0.31fF
C19594 a_2944_56872# VSS 0.35fF
C19595 a_5211_57172# VSS 1.31fF
C19596 a_3514_57167# VSS 0.32fF
C19597 a_1591_56623# VSS 0.65fF
C19598 dummypin[4] VSS 0.81fF
C19599 a_18162_58178# VSS 4.95fF
C19600 pmat.rowon_n[2] VSS 4.05fF
C19601 a_18546_58180# VSS 3.50fF
C19602 a_7521_47081# VSS 1.02fF
C19603 a_6835_51183# VSS 0.79fF
C19604 a_5528_57685# VSS 0.84fF
C19605 a_3770_57399# VSS 0.61fF
C19606 pmat.row_n[1] VSS 13.23fF
C19607 a_12967_58559# VSS 0.48fF
C19608 a_1957_43567# VSS 11.32fF
C19609 a_11711_58261# VSS 0.42fF
C19610 a_9577_58229# VSS 0.36fF
C19611 a_4719_58255# VSS 0.48fF
C19612 a_4719_30287# VSS 3.93fF
C19613 a_4720_58487# VSS 0.43fF
C19614 a_3484_58229# VSS 0.44fF
C19615 a_1823_58237# VSS 1.88fF
C19616 pmat.row_n[2] VSS 16.10fF
C19617 a_12447_16143# VSS 11.60fF
C19618 a_18162_59182# VSS 4.95fF
C19619 a_18546_59184# VSS 3.50fF
C19620 pmat.rowoff_n[6] VSS 1.37fF
C19621 a_3746_58487# VSS 5.05fF
C19622 a_6927_30503# VSS 6.61fF
C19623 a_3938_58229# VSS 1.24fF
C19624 a_6559_57167# VSS 0.90fF
C19625 a_2944_59048# VSS 0.50fF
C19626 a_2163_58941# VSS 0.48fF
C19627 a_1923_53055# VSS 2.87fF
C19628 a_1643_58773# VSS 0.38fF
C19629 pmat.rowoff_n[5] VSS 1.16fF
C19630 a_9963_13967# VSS 10.55fF
C19631 pmat.rowon_n[3] VSS 12.94fF
C19632 a_5341_59317# VSS 0.35fF
C19633 a_4956_59317# VSS 0.33fF
C19634 a_3956_59317# VSS 0.80fF
C19635 a_3175_59585# VSS 0.56fF
C19636 a_2655_59317# VSS 0.37fF
C19637 a_1591_31599# VSS 3.51fF
C19638 a_18162_60186# VSS 4.97fF
C19639 a_18546_60188# VSS 3.50fF
C19640 a_10515_13967# VSS 11.99fF
C19641 pmat.rowoff_n[11] VSS 1.11fF
C19642 a_1769_47919# VSS 4.08fF
C19643 a_5682_56311# VSS 2.30fF
C19644 a_4043_59861# VSS 0.57fF
C19645 a_1591_58799# VSS 1.15fF
C19646 a_1644_59861# VSS 0.30fF
C19647 pmat.row_n[3] VSS 13.53fF
C19648 pmat.rowon_n[4] VSS 3.89fF
C19649 a_12155_60751# VSS 0.61fF
C19650 a_11711_60751# VSS 0.53fF
C19651 a_11007_58229# VSS 2.63fF
C19652 a_10878_58487# VSS 1.59fF
C19653 a_9240_60751# VSS 0.31fF
C19654 a_8599_60751# VSS 0.34fF
C19655 a_8841_60405# VSS 0.48fF
C19656 a_8569_60405# VSS 0.33fF
C19657 a_4843_54826# VSS 1.63fF
C19658 a_3891_60431# VSS 0.52fF
C19659 adc_top_85.HI VSS 0.36fF
C19660 a_18162_61190# VSS 4.95fF
C19661 pmat.rowon_n[5] VSS 3.99fF
C19662 a_18546_61192# VSS 3.50fF
C19663 pmat.row_n[4] VSS 16.24fF
C19664 pmat.rowoff_n[9] VSS 1.21fF
C19665 a_9135_60967# VSS 7.49fF
C19666 a_2263_43719# VSS 11.99fF
C19667 a_10195_59861# VSS 0.34fF
C19668 a_4041_61225# VSS 0.34fF
C19669 a_4081_61127# VSS 0.60fF
C19670 a_1823_60949# VSS 0.62fF
C19671 a_11435_58791# VSS 11.53fF
C19672 a_11067_16359# VSS 10.98fF
C19673 a_8193_61493# VSS 0.58fF
C19674 a_7808_61493# VSS 0.33fF
C19675 a_5535_57993# VSS 1.89fF
C19676 a_5731_58951# VSS 1.06fF
C19677 a_2163_61761# VSS 0.50fF
C19678 a_1643_61493# VSS 0.39fF
C19679 _1224_.X VSS 26.44fF
C19680 a_82863_64213# VSS 1.06fF
C19681 dummypin[3] VSS 0.91fF
C19682 adc_top_84.HI VSS 0.34fF
C19683 a_18162_62194# VSS 4.97fF
C19684 pmat.rowon_n[6] VSS 3.80fF
C19685 a_18546_62196# VSS 3.50fF
C19686 a_10239_14183# VSS 11.56fF
C19687 pmat.row_n[5] VSS 13.96fF
C19688 a_2944_61493# VSS 1.00fF
C19689 a_12107_62037# VSS 0.48fF
C19690 a_10190_60663# VSS 2.19fF
C19691 a_10286_60405# VSS 0.62fF
C19692 a_7457_62037# VSS 0.57fF
C19693 a_5784_52423# VSS 1.60fF
C19694 a_4317_62215# VSS 0.69fF
C19695 a_4220_62037# VSS 0.36fF
C19696 pmat.rowoff_n[4] VSS 11.88fF
C19697 a_13656_62927# VSS 0.32fF
C19698 a_12429_62607# VSS 0.49fF
C19699 a_12985_62581# VSS 0.30fF
C19700 a_12081_62723# VSS 0.32fF
C19701 a_10391_62911# VSS 0.63fF
C19702 a_9135_62613# VSS 0.45fF
C19703 a_7212_62607# VSS 0.41fF
C19704 a_6175_60039# VSS 1.14fF
C19705 a_4025_54965# VSS 4.05fF
C19706 a_5357_62779# VSS 0.95fF
C19707 a_3305_62607# VSS 0.30fF
C19708 a_3345_62839# VSS 0.89fF
C19709 a_2215_47375# VSS 3.59fF
C19710 a_1591_61519# VSS 0.74fF
C19711 a_1644_62581# VSS 0.30fF
C19712 a_18162_63198# VSS 4.95fF
C19713 a_18546_63200# VSS 3.50fF
C19714 pmat.rowoff_n[10] VSS 1.12fF
C19715 a_12076_62839# VSS 0.38fF
C19716 a_4509_62037# VSS 0.52fF
C19717 a_3784_62607# VSS 0.54fF
C19718 a_7563_63303# VSS 0.54fF
C19719 a_7364_63303# VSS 0.78fF
C19720 a_2467_63125# VSS 0.61fF
C19721 a_18162_64202# VSS 4.95fF
C19722 a_18546_64204# VSS 3.50fF
C19723 pmat.row_n[6] VSS 13.25fF
C19724 a_10515_61839# VSS 7.14fF
C19725 a_11067_64015# VSS 8.75fF
C19726 a_4266_63303# VSS 1.04fF
C19727 a_7797_63151# VSS 0.59fF
C19728 a_8656_63811# VSS 0.31fF
C19729 a_8695_63937# VSS 0.61fF
C19730 a_8175_63669# VSS 0.39fF
C19731 a_6568_59887# VSS 0.45fF
C19732 a_5065_63669# VSS 0.40fF
C19733 a_4680_63669# VSS 0.34fF
C19734 a_2847_63999# VSS 0.41fF
C19735 a_1591_63701# VSS 0.40fF
C19736 a_10515_15055# VSS 10.55fF
C19737 nmat.rowon_n[7] VSS 15.42fF
C19738 a_10055_31591# VSS 10.62fF
C19739 pmat.rowoff_n[7] VSS 10.21fF
C19740 a_1823_64213# VSS 0.92fF
C19741 a_1644_64213# VSS 0.30fF
C19742 a_18162_65206# VSS 4.97fF
C19743 pmat.rowon_n[9] VSS 3.99fF
C19744 a_18546_65208# VSS 3.50fF
C19745 a_11203_62037# VSS 0.39fF
C19746 a_13979_65087# VSS 0.38fF
C19747 a_12723_64789# VSS 0.47fF
C19748 a_11713_64899# VSS 0.32fF
C19749 a_10049_60663# VSS 2.52fF
C19750 a_10707_64783# VSS 0.32fF
C19751 a_10569_64489# VSS 0.40fF
C19752 a_9287_65087# VSS 0.44fF
C19753 a_8031_64789# VSS 0.52fF
C19754 a_4128_64391# VSS 6.19fF
C19755 a_3751_64757# VSS 0.47fF
C19756 pmat.row_n[7] VSS 18.61fF
C19757 pmat.rowon_n[7] VSS 15.72fF
C19758 pmat.row_n[8] VSS 17.39fF
C19759 pmat.row_n[9] VSS 16.27fF
C19760 a_5462_62215# VSS 3.55fF
C19761 a_5399_65479# VSS 1.46fF
C19762 a_2944_65576# VSS 0.52fF
C19763 a_2163_65469# VSS 0.43fF
C19764 a_1643_65301# VSS 0.39fF
C19765 _1154_.X VSS 37.18fF
C19766 a_82818_69135# VSS 1.98fF
C19767 _1154_.A VSS 18.48fF
C19768 dummypin[2] VSS 0.95fF
C19769 adc_top_83.HI VSS 0.34fF
C19770 a_18162_66210# VSS 4.97fF
C19771 pmat.rowon_n[10] VSS 4.22fF
C19772 a_18546_66212# VSS 3.50fF
C19773 a_14839_66103# VSS 1.96fF
C19774 pmat.rowon_n[8] VSS 9.10fF
C19775 a_5595_65301# VSS 0.63fF
C19776 a_6612_65845# VSS 0.45fF
C19777 a_3727_66113# VSS 0.64fF
C19778 a_3207_65845# VSS 0.37fF
C19779 a_1586_63927# VSS 9.99fF
C19780 a_1591_65327# VSS 1.93fF
C19781 a_10921_64786# VSS 0.66fF
C19782 a_13919_65871# VSS 0.51fF
C19783 a_12993_66415# VSS 0.37fF
C19784 a_14289_66421# VSS 0.32fF
C19785 a_12217_66389# VSS 1.04fF
C19786 a_18162_67214# VSS 4.95fF
C19787 a_18546_67216# VSS 3.50fF
C19788 pmat.rowoff_n[8] VSS 4.87fF
C19789 a_13973_66933# VSS 0.96fF
C19790 a_13432_62581# VSS 3.05fF
C19791 a_13763_67191# VSS 0.35fF
C19792 a_11797_60431# VSS 1.14fF
C19793 a_11883_62063# VSS 1.14fF
C19794 a_9643_66389# VSS 0.84fF
C19795 a_9552_67191# VSS 0.31fF
C19796 a_8819_67197# VSS 0.70fF
C19797 a_6612_66933# VSS 0.46fF
C19798 a_4298_67191# VSS 1.52fF
C19799 a_4037_66933# VSS 0.35fF
C19800 a_1823_66941# VSS 1.15fF
C19801 a_1644_66933# VSS 0.31fF
C19802 pmat.row_n[10] VSS 14.54fF
C19803 pmat.row_n[11] VSS 16.69fF
C19804 pmat.rowon_n[11] VSS 8.38fF
C19805 pmat.rowoff_n[13] VSS 1.17fF
C19806 a_4396_66933# VSS 0.54fF
C19807 a_3983_67503# VSS 0.60fF
C19808 a_14641_57711# VSS 0.77fF
C19809 a_11142_64783# VSS 0.79fF
C19810 a_9405_66627# VSS 1.11fF
C19811 a_7899_67477# VSS 0.50fF
C19812 a_5307_67655# VSS 1.27fF
C19813 a_4421_67477# VSS 0.37fF
C19814 a_4036_67477# VSS 0.36fF
C19815 a_2944_67752# VSS 0.96fF
C19816 a_2163_67645# VSS 0.55fF
C19817 a_1643_67477# VSS 0.37fF
C19818 a_18162_68218# VSS 4.95fF
C19819 pmat.rowon_n[12] VSS 4.15fF
C19820 a_18546_68220# VSS 3.50fF
C19821 a_9545_66567# VSS 0.78fF
C19822 a_12597_68279# VSS 0.96fF
C19823 a_12500_68021# VSS 0.33fF
C19824 a_7435_68021# VSS 0.61fF
C19825 a_5651_66975# VSS 8.83fF
C19826 a_3923_68021# VSS 2.16fF
C19827 pmat.rowoff_n[12] VSS 11.81fF
C19828 a_13718_68591# VSS 0.62fF
C19829 a_13575_68743# VSS 0.70fF
C19830 a_11837_68591# VSS 0.45fF
C19831 a_4985_51433# VSS 3.17fF
C19832 a_4075_68583# VSS 2.23fF
C19833 a_10991_68591# VSS 0.94fF
C19834 a_13279_68841# VSS 0.33fF
C19835 a_1823_68565# VSS 1.07fF
C19836 a_18162_69222# VSS 4.95fF
C19837 pmat.rowon_n[13] VSS 4.19fF
C19838 a_18546_69224# VSS 3.50fF
C19839 a_14287_69455# VSS 1.81fF
C19840 pmat.row_n[12] VSS 14.07fF
C19841 a_12789_68021# VSS 0.68fF
C19842 a_4583_68021# VSS 2.62fF
C19843 a_8538_69455# VSS 0.77fF
C19844 a_7674_69455# VSS 0.50fF
C19845 a_7674_69135# VSS 0.44fF
C19846 a_4298_69367# VSS 0.59fF
C19847 a_3508_69135# VSS 0.33fF
C19848 a_4037_69109# VSS 0.34fF
C19849 a_3029_69135# VSS 0.31fF
C19850 a_3069_69367# VSS 0.84fF
C19851 a_18162_70226# VSS 4.96fF
C19852 pmat.rowon_n[14] VSS 4.03fF
C19853 a_18546_70228# VSS 3.50fF
C19854 a_12719_69367# VSS 0.62fF
C19855 a_12152_66415# VSS 0.51fF
C19856 a_12067_67279# VSS 0.53fF
C19857 a_10864_68565# VSS 0.91fF
C19858 a_11487_69653# VSS 0.53fF
C19859 a_10391_69653# VSS 0.43fF
C19860 a_9301_69679# VSS 0.32fF
C19861 a_9139_68841# VSS 0.48fF
C19862 a_9135_69679# VSS 0.52fF
C19863 a_7730_69109# VSS 1.16fF
C19864 a_8439_69653# VSS 0.41fF
C19865 a_5497_62839# VSS 0.81fF
C19866 a_4719_69929# VSS 0.35fF
C19867 a_2419_69455# VSS 5.34fF
C19868 a_2944_69928# VSS 0.95fF
C19869 a_2163_69821# VSS 0.53fF
C19870 a_1643_69653# VSS 0.40fF
C19871 pmat.rowoff_n[14] VSS 1.19fF
C19872 a_14641_57167# VSS 0.82fF
C19873 a_14287_70543# VSS 1.62fF
C19874 pmat.row_n[14] VSS 17.05fF
C19875 a_8727_70197# VSS 0.36fF
C19876 a_1674_57711# VSS 7.68fF
C19877 a_5363_70543# VSS 5.12fF
C19878 a_3936_70197# VSS 0.46fF
C19879 a_3838_70455# VSS 0.42fF
C19880 a_2387_70483# VSS 0.48fF
C19881 a_1591_67503# VSS 0.54fF
C19882 pmat.row_n[13] VSS 14.77fF
C19883 a_1923_61759# VSS 10.17fF
C19884 a_18162_71230# VSS 4.97fF
C19885 a_18546_71232# VSS 3.53fF
C19886 a_4396_69109# VSS 0.70fF
C19887 a_3710_70455# VSS 0.44fF
C19888 a_12809_69679# VSS 0.54fF
C19889 a_5081_53135# VSS 4.64fF
C19890 a_4421_70741# VSS 0.35fF
C19891 a_4036_70741# VSS 0.40fF
C19892 a_13966_71631# VSS 0.73fF
C19893 a_13102_71631# VSS 0.52fF
C19894 a_13102_71311# VSS 0.63fF
C19895 a_11693_70767# VSS 0.39fF
C19896 a_8919_71615# VSS 0.46fF
C19897 a_7663_71317# VSS 0.55fF
C19898 a_4991_69831# VSS 6.33fF
C19899 a_4225_71311# VSS 0.34fF
C19900 a_2727_58470# VSS 2.57fF
C19901 a_4265_71543# VSS 0.44fF
C19902 a_1591_69679# VSS 1.19fF
C19903 a_1644_71285# VSS 0.32fF
C19904 pmat.rowon_n[15] VSS 4.37fF
C19905 a_51202_72194# VSS 0.48fF
C19906 a_50198_72194# VSS 0.40fF
C19907 pmat.col_n[31] VSS 15.23fF
C19908 a_49194_72194# VSS 0.40fF
C19909 pmat.col_n[30] VSS 9.53fF
C19910 a_48190_72194# VSS 0.39fF
C19911 pmat.col_n[29] VSS 8.93fF
C19912 a_47186_72194# VSS 0.39fF
C19913 pmat.col_n[28] VSS 9.08fF
C19914 a_46182_72194# VSS 0.39fF
C19915 pmat.col_n[27] VSS 8.65fF
C19916 a_45178_72194# VSS 0.40fF
C19917 pmat.col_n[26] VSS 8.63fF
C19918 a_44174_72194# VSS 0.39fF
C19919 pmat.col_n[25] VSS 8.73fF
C19920 a_43170_72194# VSS 0.39fF
C19921 pmat.col_n[24] VSS 8.44fF
C19922 a_42166_72194# VSS 0.39fF
C19923 pmat.col_n[23] VSS 8.58fF
C19924 a_41162_72194# VSS 0.40fF
C19925 pmat.col_n[22] VSS 8.41fF
C19926 a_40158_72194# VSS 0.39fF
C19927 pmat.col_n[21] VSS 8.83fF
C19928 a_39154_72194# VSS 0.39fF
C19929 pmat.col_n[20] VSS 8.36fF
C19930 a_38150_72194# VSS 0.39fF
C19931 pmat.col_n[19] VSS 9.03fF
C19932 a_37146_72194# VSS 0.40fF
C19933 pmat.col_n[18] VSS 8.52fF
C19934 a_36142_72194# VSS 0.39fF
C19935 pmat.col_n[17] VSS 8.04fF
C19936 a_35138_72194# VSS 0.39fF
C19937 pmat.col_n[16] VSS 8.01fF
C19938 a_34134_72194# VSS 0.40fF
C19939 pmat.col_n[15] VSS 8.18fF
C19940 a_33130_72194# VSS 0.40fF
C19941 pmat.col_n[14] VSS 8.50fF
C19942 a_32126_72194# VSS 0.39fF
C19943 pmat.col_n[13] VSS 8.50fF
C19944 a_31122_72194# VSS 0.39fF
C19945 pmat.col_n[12] VSS 8.57fF
C19946 a_30118_72194# VSS 0.40fF
C19947 pmat.col_n[11] VSS 8.44fF
C19948 a_29114_72194# VSS 0.40fF
C19949 pmat.col_n[10] VSS 8.51fF
C19950 a_28110_72194# VSS 0.39fF
C19951 pmat.col_n[9] VSS 8.37fF
C19952 a_27106_72194# VSS 0.39fF
C19953 pmat.col_n[8] VSS 8.63fF
C19954 a_26102_72194# VSS 0.40fF
C19955 pmat.col_n[7] VSS 8.39fF
C19956 a_25098_72194# VSS 0.40fF
C19957 pmat.col_n[6] VSS 8.39fF
C19958 a_24094_72194# VSS 0.39fF
C19959 pmat.col_n[5] VSS 8.44fF
C19960 a_23090_72194# VSS 0.39fF
C19961 pmat.col_n[4] VSS 8.39fF
C19962 a_22086_72194# VSS 0.40fF
C19963 pmat.col_n[3] VSS 8.57fF
C19964 a_21082_72194# VSS 0.40fF
C19965 pmat.col_n[2] VSS 8.44fF
C19966 a_20078_72194# VSS 0.39fF
C19967 pmat.col_n[1] VSS 8.17fF
C19968 a_19074_72194# VSS 0.39fF
C19969 a_18162_72234# VSS 5.70fF
C19970 pmat.row_n[15] VSS 17.26fF
C19971 a_3615_71631# VSS 9.68fF
C19972 a_13158_71285# VSS 1.20fF
C19973 a_5779_71285# VSS 1.65fF
C19974 a_2419_53351# VSS 9.65fF
C19975 a_2791_57703# VSS 6.19fF
C19976 a_13605_71017# VSS 0.39fF
C19977 a_12249_71311# VSS 0.47fF
C19978 a_12131_71829# VSS 0.34fF
C19979 a_11115_71285# VSS 0.90fF
C19980 a_11019_71543# VSS 0.68fF
C19981 a_9375_72007# VSS 1.08fF
C19982 a_9279_71829# VSS 1.20fF
C19983 a_8283_71829# VSS 0.57fF
C19984 a_6244_71829# VSS 0.41fF
C19985 a_3866_57399# VSS 2.38fF
C19986 a_2944_72104# VSS 0.67fF
C19987 a_2163_71997# VSS 0.40fF
C19988 a_1643_71829# VSS 0.40fF
C19989 pmat.col_n[0] VSS 8.57fF
C19990 pmat.sample VSS 12.47fF
C19991 a_18546_72236# VSS 8.97fF
C19992 pmat.sample_n VSS 17.04fF
C19993 a_13327_70741# VSS 1.65fF
C19994 a_14439_72703# VSS 0.39fF
C19995 a_13183_72405# VSS 0.46fF
C19996 a_4075_50087# VSS 6.49fF
C19997 a_5232_72373# VSS 0.31fF
C19998 a_3956_72373# VSS 0.99fF
C19999 a_3175_72641# VSS 0.56fF
C20000 a_2655_72373# VSS 0.36fF
C20001 pmat.rowoff_n[15] VSS 10.17fF
C20002 a_6451_67655# VSS 3.36fF
C20003 a_8491_47911# VSS 9.08fF
C20004 a_3339_70759# VSS 7.64fF
C20005 a_2879_57487# VSS 8.80fF
C20006 a_10699_72943# VSS 0.72fF
C20007 a_5687_71829# VSS 1.52fF
C20008 a_11271_73085# VSS 0.54fF
C20009 a_10751_72917# VSS 0.38fF
C20010 a_1591_71855# VSS 0.89fF
C20011 a_1644_72917# VSS 0.32fF
C20012 a_9103_73791# VSS 0.45fF
C20013 a_8013_73493# VSS 0.34fF
C20014 a_5403_67655# VSS 0.71fF
C20015 a_7847_73493# VSS 0.63fF
C20016 dummypin[1] VSS 1.00fF
C20017 adc_top_82.HI VSS 0.34fF
C20018 a_7099_74313# VSS 0.77fF
C20019 a_2407_49289# VSS 7.96fF
C20020 a_9831_74183# VSS 0.38fF
C20021 a_9655_74216# VSS 0.38fF
C20022 a_4697_74005# VSS 0.51fF
C20023 a_4409_74183# VSS 0.73fF
C20024 a_4312_74005# VSS 0.34fF
C20025 a_1899_35051# VSS 10.30fF
C20026 a_2163_74173# VSS 0.42fF
C20027 a_1643_74005# VSS 0.39fF
C20028 a_14071_74879# VSS 0.44fF
C20029 a_12981_74581# VSS 0.32fF
C20030 a_6292_65479# VSS 4.85fF
C20031 a_12815_74581# VSS 0.56fF
C20032 a_7111_74575# VSS 0.42fF
C20033 a_4351_55527# VSS 4.97fF
C20034 a_4048_74549# VSS 0.43fF
C20035 a_3228_74691# VSS 0.31fF
C20036 a_3267_74817# VSS 0.48fF
C20037 a_2747_74549# VSS 0.38fF
C20038 a_1823_74557# VSS 0.80fF
C20039 a_4259_73807# VSS 3.82fF
C20040 a_7092_74005# VSS 0.56fF
C20041 a_1591_74031# VSS 0.36fF
C20042 a_6787_47607# VSS 8.44fF
C20043 a_10697_75218# VSS 1.40fF
C20044 a_9581_73487# VSS 1.19fF
C20045 a_10515_75895# VSS 1.33fF
C20046 a_6051_74183# VSS 0.66fF
C20047 a_11397_76457# VSS 0.50fF
C20048 a_11023_76359# VSS 0.40fF
C20049 a_8539_76181# VSS 0.41fF
C20050 a_5497_73719# VSS 0.75fF
C20051 a_2149_45717# VSS 9.68fF
C20052 a_1823_76181# VSS 1.47fF
C20053 a_1644_76181# VSS 0.32fF
C20054 a_9287_77055# VSS 0.39fF
C20055 a_6292_69831# VSS 1.38fF
C20056 a_8031_76757# VSS 0.44fF
C20057 a_4123_76181# VSS 0.73fF
C20058 a_6975_76823# VSS 2.73fF
C20059 a_6795_76989# VSS 1.16fF
C20060 a_4429_76751# VSS 0.40fF
C20061 a_5047_76983# VSS 0.32fF
C20062 a_3951_77055# VSS 0.46fF
C20063 a_2999_76922# VSS 0.42fF
C20064 a_2695_76757# VSS 0.41fF
C20065 a_2099_76725# VSS 0.51fF
C20066 dummypin[0] VSS 0.97fF
C20067 a_7658_71543# VSS 3.62fF
C20068 a_10239_77295# VSS 1.13fF
C20069 a_6799_75637# VSS 0.68fF
C20070 a_6200_70919# VSS 1.57fF
C20071 a_10811_77437# VSS 0.56fF
C20072 a_3339_59879# VSS 11.12fF
C20073 a_10291_77269# VSS 0.41fF
C20074 a_6803_77269# VSS 0.42fF
C20075 a_1923_69823# VSS 8.59fF
C20076 a_5725_76207# VSS 0.39fF
C20077 a_5547_77295# VSS 0.44fF
C20078 a_1674_68047# VSS 5.64fF
C20079 adc_top_81.HI VSS 0.38fF
C20080 a_1823_77821# VSS 0.64fF
C20081 a_1644_77813# VSS 0.35fF
C20082 VDD VSS 22121.70fF
.ends

