* SPICE3 file created from adc_noise_decoup_cell2.ext - technology: sky130A

.subckt adc_noise_decoup_cell2 nmoscap_bot mimcap_bot mimcap_top nmoscap_top pwell
X0 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.576e+13p pd=7.64e+07u as=0p ps=0u w=1.84e+07u l=3.9e+06u
X1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=5.1e+06u w=1.89e+07u
C0 mimcap_top nmoscap_top 2.67fF
C1 nmoscap_top nmoscap_bot 142.82fF
C2 mimcap_top mimcap_bot 16.54fF
C3 mimcap_bot nmoscap_top 5.71fF
C4 mimcap_bot nmoscap_bot 6.30fF
C5 mimcap_top pwell 2.02fF
C6 nmoscap_top pwell 7.01fF
C7 nmoscap_bot pwell 6.37fF
.ends
