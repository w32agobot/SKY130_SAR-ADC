VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO emptybox_10_30
  CLASS BLOCK ;
  FOREIGN emptybox_10_30 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 30.000 ;
  OBS
      LAYER met1 ;
        RECT 0 0 10 30 ;
  END
END emptybox_10_30
END LIBRARY

