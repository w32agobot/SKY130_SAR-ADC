magic
tech sky130A
magscale 1 2
timestamp 1671464254
<< nwell >>
rect 0 506 1004 880
<< nmos >>
rect 232 212 262 296
rect 328 212 358 296
rect 536 252 566 336
rect 632 252 662 336
rect 728 252 758 336
<< pmos >>
rect 232 542 262 702
rect 328 542 358 702
rect 536 574 566 734
rect 632 574 662 734
rect 728 574 758 734
<< ndiff >>
rect 474 324 536 336
rect 170 256 232 296
rect 170 222 182 256
rect 216 222 232 256
rect 170 212 232 222
rect 262 284 328 296
rect 262 224 278 284
rect 312 224 328 284
rect 262 212 328 224
rect 358 284 420 296
rect 358 224 374 284
rect 408 224 420 284
rect 474 264 486 324
rect 520 264 536 324
rect 474 252 536 264
rect 566 324 632 336
rect 566 264 582 324
rect 616 264 632 324
rect 566 252 632 264
rect 662 324 728 336
rect 662 264 678 324
rect 712 264 728 324
rect 662 252 728 264
rect 758 324 820 336
rect 758 264 774 324
rect 808 264 820 324
rect 758 252 820 264
rect 358 212 420 224
<< pdiff >>
rect 474 722 536 734
rect 170 690 232 702
rect 170 554 182 690
rect 216 554 232 690
rect 170 542 232 554
rect 262 690 328 702
rect 262 554 278 690
rect 312 554 328 690
rect 262 542 328 554
rect 358 690 420 702
rect 358 554 374 690
rect 408 554 420 690
rect 474 586 486 722
rect 520 586 536 722
rect 474 574 536 586
rect 566 722 632 734
rect 566 586 582 722
rect 616 586 632 722
rect 566 574 632 586
rect 662 722 728 734
rect 662 586 678 722
rect 712 586 728 722
rect 662 574 728 586
rect 758 722 820 734
rect 758 586 774 722
rect 808 586 820 722
rect 758 574 820 586
rect 358 542 420 554
<< ndiffc >>
rect 182 222 216 256
rect 278 224 312 284
rect 374 224 408 284
rect 486 264 520 324
rect 582 264 616 324
rect 678 264 712 324
rect 774 264 808 324
<< pdiffc >>
rect 182 554 216 690
rect 278 554 312 690
rect 374 554 408 690
rect 486 586 520 722
rect 582 586 616 722
rect 678 586 712 722
rect 774 586 808 722
<< psubdiff >>
rect 570 148 628 182
rect 662 148 726 182
rect 760 148 792 182
<< nsubdiff >>
rect 302 838 806 844
rect 302 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 302 798 806 804
<< psubdiffcont >>
rect 628 148 662 182
rect 726 148 760 182
<< nsubdiffcont >>
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
<< poly >>
rect 212 818 280 828
rect 212 782 228 818
rect 264 782 280 818
rect 212 718 280 782
rect 536 734 566 760
rect 632 734 662 760
rect 728 734 758 760
rect 232 702 262 718
rect 328 702 358 728
rect 232 296 262 542
rect 328 508 358 542
rect 536 536 566 574
rect 632 548 662 574
rect 728 558 758 574
rect 494 516 566 536
rect 328 488 416 508
rect 328 450 370 488
rect 404 450 416 488
rect 328 328 416 450
rect 494 482 510 516
rect 544 482 566 516
rect 494 448 566 482
rect 608 526 676 548
rect 728 528 834 558
rect 608 492 624 526
rect 660 492 676 526
rect 608 480 676 492
rect 766 520 834 528
rect 766 486 782 520
rect 818 486 834 520
rect 766 476 834 486
rect 494 414 510 448
rect 544 414 566 448
rect 644 426 676 430
rect 494 398 566 414
rect 536 336 566 398
rect 608 410 676 426
rect 608 376 624 410
rect 660 376 676 410
rect 608 362 676 376
rect 632 336 662 362
rect 728 336 758 362
rect 328 296 358 328
rect 536 226 566 252
rect 632 226 662 252
rect 728 236 758 252
rect 728 220 888 236
rect 232 186 262 212
rect 328 186 358 212
rect 728 206 844 220
rect 834 186 844 206
rect 878 186 888 220
rect 834 170 888 186
<< polycont >>
rect 228 782 264 818
rect 370 450 404 488
rect 510 482 544 516
rect 624 492 660 526
rect 782 486 818 520
rect 510 414 544 448
rect 624 376 660 410
rect 844 186 878 220
<< locali >>
rect 34 922 182 1004
rect 34 888 48 922
rect 134 888 182 922
rect 34 882 182 888
rect 910 922 970 1004
rect 910 888 923 922
rect 958 888 970 922
rect 910 882 970 888
rect 34 704 148 882
rect 302 838 806 844
rect 228 818 264 834
rect 302 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 302 798 806 804
rect 228 772 264 782
rect 228 738 230 772
rect 374 722 520 738
rect 374 706 486 722
rect 34 630 48 704
rect 136 630 148 704
rect 34 338 148 630
rect 34 292 48 338
rect 130 292 148 338
rect 182 690 216 706
rect 182 340 216 554
rect 278 690 312 706
rect 278 330 312 554
rect 374 690 432 706
rect 408 672 432 690
rect 466 672 486 706
rect 408 586 486 672
rect 408 570 520 586
rect 582 722 616 798
rect 582 570 616 586
rect 678 722 712 762
rect 408 554 476 570
rect 678 560 712 586
rect 774 722 808 738
rect 774 570 808 586
rect 374 538 476 554
rect 370 488 404 504
rect 370 380 404 450
rect 370 340 404 346
rect 442 340 476 538
rect 608 492 624 526
rect 660 492 744 526
rect 510 448 544 482
rect 510 398 544 414
rect 608 410 644 424
rect 608 376 624 410
rect 660 376 676 410
rect 710 408 744 492
rect 782 520 818 536
rect 782 476 818 486
rect 856 408 970 882
rect 710 374 970 408
rect 34 106 148 292
rect 442 324 520 340
rect 442 300 486 324
rect 278 284 312 296
rect 182 256 216 272
rect 182 174 216 222
rect 278 208 312 224
rect 374 284 408 300
rect 374 208 408 224
rect 486 174 520 264
rect 582 326 616 340
rect 582 248 616 264
rect 678 324 712 340
rect 678 182 712 264
rect 774 326 808 340
rect 774 248 808 264
rect 856 338 970 374
rect 856 292 870 338
rect 956 292 970 338
rect 856 236 970 292
rect 840 220 970 236
rect 840 186 844 220
rect 878 186 970 220
rect 182 140 520 174
rect 570 148 628 182
rect 662 148 726 182
rect 760 148 792 182
rect 840 170 970 186
rect 856 108 970 170
rect 34 102 182 106
rect 34 68 48 102
rect 134 68 182 102
rect 34 0 182 68
rect 910 102 970 108
rect 910 68 922 102
rect 958 68 970 102
rect 910 0 970 68
<< viali >>
rect 48 888 134 922
rect 923 888 958 922
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
rect 230 738 264 772
rect 48 630 136 704
rect 48 292 130 338
rect 182 306 216 340
rect 432 672 466 706
rect 774 672 808 706
rect 370 346 404 380
rect 510 516 544 532
rect 510 498 544 516
rect 608 424 644 458
rect 782 442 818 476
rect 278 296 312 330
rect 374 234 408 268
rect 582 324 616 326
rect 582 292 616 324
rect 774 324 808 326
rect 774 292 808 324
rect 870 292 956 338
rect 628 148 662 182
rect 726 148 760 182
rect 48 68 134 102
rect 922 68 958 102
<< metal1 >>
rect 34 922 182 1004
rect 34 888 48 922
rect 134 888 182 922
rect 34 882 182 888
rect 910 922 970 1004
rect 910 888 923 922
rect 958 888 970 922
rect 910 882 970 888
rect 0 838 1004 854
rect 0 806 326 838
rect 0 798 196 806
rect 298 804 326 806
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 1004 838
rect 298 798 1004 804
rect 218 772 276 778
rect 218 770 230 772
rect 0 740 230 770
rect 218 738 230 740
rect 264 770 276 772
rect 264 740 1004 770
rect 264 738 276 740
rect 218 732 276 738
rect 34 704 148 712
rect 34 630 48 704
rect 136 630 148 704
rect 420 706 820 712
rect 420 672 432 706
rect 466 672 774 706
rect 808 672 820 706
rect 420 666 820 672
rect 34 624 148 630
rect 0 568 1004 596
rect 0 532 1004 540
rect 0 512 510 532
rect 496 498 510 512
rect 544 512 1004 532
rect 544 498 554 512
rect 496 486 554 498
rect 770 476 830 484
rect 594 458 656 464
rect 770 458 782 476
rect 0 430 608 458
rect 594 424 608 430
rect 644 442 782 458
rect 818 458 830 476
rect 818 442 1004 458
rect 644 430 1004 442
rect 644 424 656 430
rect 594 418 656 424
rect 0 390 416 402
rect 736 390 1004 402
rect 0 380 1004 390
rect 0 374 370 380
rect 358 346 370 374
rect 404 374 1004 380
rect 404 362 816 374
rect 404 346 416 362
rect 34 338 142 346
rect 34 292 48 338
rect 130 292 142 338
rect 170 340 228 346
rect 170 306 182 340
rect 216 306 228 340
rect 170 300 228 306
rect 34 286 142 292
rect 182 258 216 300
rect 266 288 272 340
rect 324 288 330 340
rect 358 334 416 346
rect 856 338 970 346
rect 570 326 820 334
rect 570 292 582 326
rect 616 292 774 326
rect 808 292 820 326
rect 368 268 416 290
rect 570 286 820 292
rect 856 292 870 338
rect 956 292 970 338
rect 856 286 970 292
rect 368 258 374 268
rect 0 234 374 258
rect 408 258 416 268
rect 408 234 1004 258
rect 0 220 1004 234
rect 0 182 1004 192
rect 0 148 628 182
rect 662 148 726 182
rect 760 148 1004 182
rect 0 136 1004 148
rect 34 102 182 108
rect 34 68 48 102
rect 134 68 182 102
rect 34 0 182 68
rect 910 102 970 108
rect 910 68 922 102
rect 958 68 970 102
rect 910 0 970 68
<< via1 >>
rect 272 330 324 340
rect 272 296 278 330
rect 278 296 312 330
rect 312 296 324 330
rect 272 288 324 296
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 770 972 810
rect 32 714 42 770
rect 98 714 330 770
rect 386 714 618 770
rect 674 714 906 770
rect 962 714 972 770
rect 32 674 972 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 32 608 972 618
rect 32 578 396 608
rect 32 522 42 578
rect 98 522 330 578
rect 386 522 396 578
rect 608 578 972 608
rect 32 482 396 522
rect 32 426 42 482
rect 98 426 330 482
rect 386 426 396 482
rect 460 460 544 544
rect 608 522 618 578
rect 674 522 906 578
rect 962 522 972 578
rect 608 482 972 522
rect 32 396 396 426
rect 608 426 618 482
rect 674 426 906 482
rect 962 426 972 482
rect 608 396 972 426
rect 32 386 972 396
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 340 330 386
rect 324 330 330 340
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 972 386
rect 32 290 272 330
rect 32 234 42 290
rect 98 288 272 290
rect 324 290 972 330
rect 324 288 330 290
rect 98 234 330 288
rect 386 234 618 290
rect 674 234 906 290
rect 962 234 972 290
rect 32 194 972 234
rect 32 138 42 194
rect 98 138 330 194
rect 386 138 618 194
rect 674 138 906 194
rect 962 138 972 194
rect 32 98 972 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 32 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 330 714 386 770
rect 618 714 674 770
rect 906 714 962 770
rect 42 618 98 674
rect 138 618 194 674
rect 234 618 290 674
rect 330 618 386 674
rect 426 618 482 674
rect 522 618 578 674
rect 618 618 674 674
rect 714 618 770 674
rect 810 618 866 674
rect 906 618 962 674
rect 42 522 98 578
rect 330 522 386 578
rect 42 426 98 482
rect 330 426 386 482
rect 618 522 674 578
rect 906 522 962 578
rect 618 426 674 482
rect 906 426 962 482
rect 42 330 98 386
rect 138 330 194 386
rect 234 340 290 386
rect 234 330 272 340
rect 272 330 290 340
rect 330 330 386 386
rect 426 330 482 386
rect 522 330 578 386
rect 618 330 674 386
rect 714 330 770 386
rect 810 330 866 386
rect 906 330 962 386
rect 42 234 98 290
rect 330 234 386 290
rect 618 234 674 290
rect 906 234 962 290
rect 42 138 98 194
rect 330 138 386 194
rect 618 138 674 194
rect 906 138 962 194
rect 42 42 98 98
rect 138 42 194 98
rect 234 42 290 98
rect 330 42 386 98
rect 426 42 482 98
rect 522 42 578 98
rect 618 42 674 98
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 612 866 680 900
rect 324 770 392 810
rect 36 680 104 714
rect 324 714 330 770
rect 386 714 392 770
rect 452 824 552 840
rect 452 756 468 824
rect 536 756 552 824
rect 452 740 552 756
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 770 680 810
rect 324 680 392 714
rect 612 714 618 770
rect 674 714 680 770
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 612 680 680 714
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 36 674 968 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 36 612 968 618
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 324 578 392 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 324 522 330 578
rect 386 522 392 578
rect 324 482 392 522
rect 36 392 104 426
rect 324 426 330 482
rect 386 426 392 482
rect 324 392 392 426
rect 612 578 680 612
rect 612 522 618 578
rect 674 522 680 578
rect 900 578 968 612
rect 612 482 680 522
rect 612 426 618 482
rect 674 426 680 482
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 612 392 680 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 968 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 36 324 968 330
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 324 290 392 324
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 324 234 330 290
rect 386 234 392 290
rect 612 290 680 324
rect 324 194 392 234
rect 36 104 104 138
rect 324 138 330 194
rect 386 138 392 194
rect 452 248 552 264
rect 452 180 468 248
rect 536 180 552 248
rect 452 164 552 180
rect 612 234 618 290
rect 674 234 680 290
rect 900 290 968 324
rect 612 194 680 234
rect 324 104 392 138
rect 612 138 618 194
rect 674 138 680 194
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 612 104 680 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 968 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 36 36 968 42
<< via3 >>
rect 180 756 248 824
rect 468 756 536 824
rect 756 756 824 824
rect 180 468 248 536
rect 756 468 824 536
rect 180 180 248 248
rect 468 180 536 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 472 840 532 934
rect 760 840 820 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 452 824 552 840
rect 452 820 468 824
rect 248 760 468 820
rect 248 756 264 760
rect 164 740 264 756
rect 452 756 468 760
rect 536 820 552 824
rect 740 824 840 840
rect 740 820 756 824
rect 536 760 756 820
rect 536 756 552 760
rect 452 740 552 756
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 184 552 244 740
rect 472 646 532 740
rect 760 552 820 740
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 532 264 536
rect 740 536 840 552
rect 740 532 756 536
rect 248 472 358 532
rect 646 472 756 532
rect 248 468 264 472
rect 164 452 264 468
rect 740 468 756 472
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 184 264 244 452
rect 472 264 532 358
rect 760 264 820 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 244 264 248
rect 452 248 552 264
rect 452 244 468 248
rect 248 184 468 244
rect 248 180 264 184
rect 164 164 264 180
rect 452 180 468 184
rect 536 244 552 248
rect 740 248 840 264
rect 740 244 756 248
rect 536 184 756 244
rect 536 180 552 184
rect 452 164 552 180
rect 740 180 756 184
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 184 70 244 164
rect 472 70 532 164
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 576 576 608 608
rect 544 544 576 576
rect 428 428 460 460
rect 416 396 428 428
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
flabel metal1 0 798 167 854 0 FreeSans 160 0 0 0 VDD
port 1 w power bidirectional
flabel metal1 837 798 1004 854 0 FreeSans 160 0 0 0 VDD
port 1 e power bidirectional
flabel metal1 0 136 1004 192 0 FreeSans 320 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal1 0 220 1004 258 0 FreeSans 320 0 0 0 vcom
port 3 nsew
flabel metal4 472 874 532 934 1 FreeSans 160 0 0 0 ctop
port 4 n
flabel metal1 34 0 182 108 5 FreeSans 320 0 0 0 col
port 5 s
flabel metal1 34 882 182 1004 1 FreeSans 320 0 0 0 col
port 5 n
flabel space 910 0 970 108 1 FreeSans 320 0 0 0 col_n
port 6 s
flabel space 910 882 970 1004 1 FreeSans 320 0 0 0 col_n
port 6 n
flabel metal1 0 430 171 458 0 FreeSans 160 0 0 0 row_n
port 7 w
flabel metal1 846 430 1004 458 0 FreeSans 160 0 0 0 row_n
port 7 e
flabel metal1 0 512 171 540 0 FreeSans 160 0 0 0 rowon_n
port 8 w
flabel metal1 849 512 1004 540 0 FreeSans 160 0 0 0 rowon_n
port 8 e
flabel metal1 0 374 171 402 0 FreeSans 160 0 0 0 sample
port 9 w
flabel metal1 846 374 1004 402 0 FreeSans 160 0 0 0 sample
port 9 e
flabel metal1 0 740 1004 770 0 FreeSans 160 0 0 0 sample_n
port 10 nsew
flabel metal1 0 568 171 596 7 FreeSans 160 0 0 0 off_n
port 11 w
flabel metal1 848 568 1004 596 3 FreeSans 160 0 0 0 off_n
port 11 e
rlabel metal2 500 972 500 972 1 cbot
<< end >>
