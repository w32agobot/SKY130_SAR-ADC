magic
tech sky130A
timestamp 1662981783
<< metal2 >>
rect 16 198 198 486
rect 304 198 486 486
rect 16 16 486 198
<< metal4 >>
rect 236 366 266 467
<< comment >>
rect 0 486 16 502
rect 486 486 502 502
rect 0 0 16 16
rect 486 0 502 16
<< end >>
