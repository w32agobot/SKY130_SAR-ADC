magic
tech sky130A
timestamp 1663074849
<< psubdiff >>
rect -2157 9110 -1950 9274
rect -2157 9093 -2143 9110
rect -1968 9093 -1950 9110
rect -2157 9070 -1950 9093
rect -2157 9053 -2143 9070
rect -1968 9053 -1950 9070
rect -2157 9030 -1950 9053
rect -2157 9013 -2143 9030
rect -1968 9013 -1950 9030
rect -2157 8990 -1950 9013
rect -2157 8973 -2143 8990
rect -1968 8973 -1950 8990
rect -2157 8950 -1950 8973
rect -2157 8933 -2143 8950
rect -1968 8933 -1950 8950
rect -2157 8910 -1950 8933
rect -2157 8893 -2143 8910
rect -1968 8893 -1950 8910
rect -2157 8870 -1950 8893
rect -2157 8853 -2143 8870
rect -1968 8853 -1950 8870
rect -2157 8830 -1950 8853
rect -2157 8813 -2143 8830
rect -1968 8813 -1950 8830
rect -2157 8790 -1950 8813
rect -2157 8773 -2143 8790
rect -1968 8773 -1950 8790
rect -2157 8750 -1950 8773
rect -2157 8733 -2143 8750
rect -1968 8733 -1950 8750
rect -2157 8710 -1950 8733
rect -2157 8693 -2143 8710
rect -1968 8693 -1950 8710
rect -2157 8670 -1950 8693
rect -2157 8653 -2143 8670
rect -1968 8653 -1950 8670
rect -2157 8630 -1950 8653
rect -2157 8613 -2143 8630
rect -1968 8613 -1950 8630
rect -2157 8590 -1950 8613
rect -2157 8573 -2143 8590
rect -1968 8573 -1950 8590
rect -2157 8550 -1950 8573
rect -2157 8533 -2143 8550
rect -1968 8533 -1950 8550
rect -2157 8510 -1950 8533
rect -2157 8493 -2143 8510
rect -1968 8493 -1950 8510
rect -2157 8470 -1950 8493
rect -2157 8453 -2143 8470
rect -1968 8453 -1950 8470
rect -2157 8430 -1950 8453
rect -2157 8413 -2143 8430
rect -1968 8413 -1950 8430
rect -2157 8390 -1950 8413
rect -2157 8373 -2143 8390
rect -1968 8373 -1950 8390
rect -2157 8350 -1950 8373
rect -2157 8333 -2143 8350
rect -1968 8333 -1950 8350
rect -2157 8310 -1950 8333
rect -2157 8293 -2143 8310
rect -1968 8293 -1950 8310
rect -2157 8270 -1950 8293
rect -2157 8253 -2143 8270
rect -1968 8253 -1950 8270
rect -2157 8230 -1950 8253
rect -2157 8213 -2143 8230
rect -1968 8213 -1950 8230
rect -2157 8190 -1950 8213
rect -2157 8173 -2143 8190
rect -1968 8173 -1950 8190
rect -2157 8150 -1950 8173
rect -2157 8133 -2143 8150
rect -1968 8133 -1950 8150
rect -2157 8110 -1950 8133
rect -2157 8093 -2143 8110
rect -1968 8093 -1950 8110
rect -2157 8070 -1950 8093
rect -2157 8053 -2143 8070
rect -1968 8053 -1950 8070
rect -2157 8030 -1950 8053
rect -2157 8013 -2143 8030
rect -1968 8013 -1950 8030
rect -2157 7990 -1950 8013
rect -2157 7973 -2143 7990
rect -1968 7973 -1950 7990
rect -2157 7950 -1950 7973
rect -2157 7933 -2143 7950
rect -1968 7933 -1950 7950
rect -2157 7910 -1950 7933
rect -2157 7893 -2143 7910
rect -1968 7893 -1950 7910
rect -2157 7870 -1950 7893
rect -2157 7853 -2143 7870
rect -1968 7853 -1950 7870
rect -2157 7830 -1950 7853
rect -2157 7813 -2143 7830
rect -1968 7813 -1950 7830
rect -2157 7790 -1950 7813
rect -2157 7773 -2143 7790
rect -1968 7773 -1950 7790
rect -2157 7750 -1950 7773
rect -2157 7733 -2143 7750
rect -1968 7733 -1950 7750
rect -2157 7710 -1950 7733
rect -2157 7693 -2143 7710
rect -1968 7693 -1950 7710
rect -2157 7670 -1950 7693
rect -2157 7653 -2143 7670
rect -1968 7653 -1950 7670
rect -2157 7630 -1950 7653
rect -2157 7613 -2143 7630
rect -1968 7613 -1950 7630
rect -2157 7590 -1950 7613
rect -2157 7573 -2143 7590
rect -1968 7573 -1950 7590
rect -2157 7550 -1950 7573
rect -2157 7533 -2143 7550
rect -1968 7533 -1950 7550
rect -2157 7510 -1950 7533
rect -2157 7493 -2143 7510
rect -1968 7493 -1950 7510
rect -2157 7470 -1950 7493
rect -2157 7453 -2143 7470
rect -1968 7453 -1950 7470
rect -2157 7430 -1950 7453
rect -2157 7413 -2143 7430
rect -1968 7413 -1950 7430
rect -2157 7390 -1950 7413
rect -2157 7373 -2143 7390
rect -1968 7373 -1950 7390
rect -2157 7350 -1950 7373
rect -2157 7333 -2143 7350
rect -1968 7333 -1950 7350
rect -2157 7310 -1950 7333
rect -2157 7293 -2143 7310
rect -1968 7293 -1950 7310
rect -2157 7270 -1950 7293
rect -2157 7253 -2143 7270
rect -1968 7253 -1950 7270
rect -2157 7230 -1950 7253
rect -2157 7213 -2143 7230
rect -1968 7213 -1950 7230
rect -2157 7190 -1950 7213
rect -2157 7173 -2143 7190
rect -1968 7173 -1950 7190
rect -2157 7150 -1950 7173
rect -2157 7133 -2143 7150
rect -1968 7133 -1950 7150
rect -2157 7110 -1950 7133
rect -2157 7093 -2143 7110
rect -1968 7093 -1950 7110
rect -2157 7070 -1950 7093
rect -2157 7053 -2143 7070
rect -1968 7053 -1950 7070
rect -2157 7030 -1950 7053
rect -2157 7013 -2143 7030
rect -1968 7013 -1950 7030
rect -2157 6990 -1950 7013
rect -2157 6973 -2143 6990
rect -1968 6973 -1950 6990
rect -2157 6950 -1950 6973
rect -2157 6933 -2143 6950
rect -1968 6933 -1950 6950
rect -2157 6910 -1950 6933
rect -2157 6893 -2143 6910
rect -1968 6893 -1950 6910
rect -2157 6870 -1950 6893
rect -2157 6853 -2143 6870
rect -1968 6853 -1950 6870
rect -2157 6830 -1950 6853
rect -2157 6813 -2143 6830
rect -1968 6813 -1950 6830
rect -2157 6790 -1950 6813
rect -2157 6773 -2143 6790
rect -1968 6773 -1950 6790
rect -2157 6750 -1950 6773
rect -2157 6733 -2143 6750
rect -1968 6733 -1950 6750
rect -2157 6710 -1950 6733
rect -2157 6693 -2143 6710
rect -1968 6693 -1950 6710
rect -2157 6670 -1950 6693
rect -2157 6653 -2143 6670
rect -1968 6653 -1950 6670
rect -2157 6630 -1950 6653
rect -2157 6613 -2143 6630
rect -1968 6613 -1950 6630
rect -2157 6590 -1950 6613
rect -2157 6573 -2143 6590
rect -1968 6573 -1950 6590
rect -2157 6550 -1950 6573
rect -2157 6533 -2143 6550
rect -1968 6533 -1950 6550
rect -2157 6510 -1950 6533
rect -2157 6493 -2143 6510
rect -1968 6493 -1950 6510
rect -2157 6470 -1950 6493
rect -2157 6453 -2143 6470
rect -1968 6453 -1950 6470
rect -2157 6430 -1950 6453
rect -2157 6413 -2143 6430
rect -1968 6413 -1950 6430
rect -2157 6390 -1950 6413
rect -2157 6373 -2143 6390
rect -1968 6373 -1950 6390
rect -2157 6350 -1950 6373
rect -2157 6333 -2143 6350
rect -1968 6333 -1950 6350
rect -2157 6310 -1950 6333
rect -2157 6293 -2143 6310
rect -1968 6293 -1950 6310
rect -2157 6270 -1950 6293
rect -2157 6253 -2143 6270
rect -1968 6253 -1950 6270
rect -2157 6230 -1950 6253
rect -2157 6213 -2143 6230
rect -1968 6213 -1950 6230
rect -2157 6190 -1950 6213
rect -2157 6173 -2143 6190
rect -1968 6173 -1950 6190
rect -2157 6150 -1950 6173
rect -2157 6133 -2143 6150
rect -1968 6133 -1950 6150
rect -2157 6110 -1950 6133
rect -2157 6093 -2143 6110
rect -1968 6093 -1950 6110
rect -2157 6070 -1950 6093
rect -2157 6053 -2143 6070
rect -1968 6053 -1950 6070
rect -2157 6030 -1950 6053
rect -2157 6013 -2143 6030
rect -1968 6013 -1950 6030
rect -2157 5990 -1950 6013
rect -2157 5973 -2143 5990
rect -1968 5973 -1950 5990
rect -2157 5950 -1950 5973
rect -2157 5933 -2143 5950
rect -1968 5933 -1950 5950
rect -2157 5910 -1950 5933
rect -2157 5893 -2143 5910
rect -1968 5893 -1950 5910
rect -2157 5870 -1950 5893
rect -2157 5853 -2143 5870
rect -1968 5853 -1950 5870
rect -2157 5830 -1950 5853
rect -2157 5813 -2143 5830
rect -1968 5813 -1950 5830
rect -2157 5790 -1950 5813
rect -2157 5773 -2143 5790
rect -1968 5773 -1950 5790
rect -2157 5750 -1950 5773
rect -2157 5733 -2143 5750
rect -1968 5733 -1950 5750
rect -2157 5710 -1950 5733
rect -2157 5693 -2143 5710
rect -1968 5693 -1950 5710
rect -2157 5670 -1950 5693
rect -2157 5653 -2143 5670
rect -1968 5653 -1950 5670
rect -2157 5630 -1950 5653
rect -2157 5613 -2143 5630
rect -1968 5613 -1950 5630
rect -2157 5590 -1950 5613
rect -2157 5573 -2143 5590
rect -1968 5573 -1950 5590
rect -2157 5550 -1950 5573
rect -2157 5533 -2143 5550
rect -1968 5533 -1950 5550
rect -2157 5510 -1950 5533
rect -2157 5493 -2143 5510
rect -1968 5493 -1950 5510
rect -2157 5470 -1950 5493
rect -2157 5453 -2143 5470
rect -1968 5453 -1950 5470
rect -2157 5430 -1950 5453
rect -2157 5413 -2143 5430
rect -1968 5413 -1950 5430
rect -2157 5390 -1950 5413
rect -2157 5373 -2143 5390
rect -1968 5373 -1950 5390
rect -2157 5350 -1950 5373
rect -2157 5333 -2143 5350
rect -1968 5333 -1950 5350
rect -2157 5310 -1950 5333
rect -2157 5293 -2143 5310
rect -1968 5293 -1950 5310
rect -2157 5270 -1950 5293
rect -2157 5253 -2143 5270
rect -1968 5253 -1950 5270
rect -2157 5230 -1950 5253
rect -2157 5213 -2143 5230
rect -1968 5213 -1950 5230
rect -2157 5190 -1950 5213
rect -2157 5173 -2143 5190
rect -1968 5173 -1950 5190
rect -2157 5150 -1950 5173
rect -2157 5133 -2143 5150
rect -1968 5133 -1950 5150
rect -2157 5110 -1950 5133
rect -2157 5093 -2143 5110
rect -1968 5093 -1950 5110
rect -2157 5070 -1950 5093
rect -2157 5053 -2143 5070
rect -1968 5053 -1950 5070
rect -2157 5030 -1950 5053
rect -2157 5013 -2143 5030
rect -1968 5013 -1950 5030
rect -2157 4990 -1950 5013
rect -2157 4973 -2143 4990
rect -1968 4973 -1950 4990
rect -2157 4950 -1950 4973
rect -2157 4933 -2143 4950
rect -1968 4933 -1950 4950
rect -2157 4910 -1950 4933
rect -2157 4893 -2143 4910
rect -1968 4893 -1950 4910
rect -2157 4870 -1950 4893
rect -2157 4853 -2143 4870
rect -1968 4853 -1950 4870
rect -2157 4830 -1950 4853
rect -2157 4813 -2143 4830
rect -1968 4813 -1950 4830
rect -2157 4790 -1950 4813
rect -2157 4773 -2143 4790
rect -1968 4773 -1950 4790
rect -2157 4750 -1950 4773
rect -2157 4733 -2143 4750
rect -1968 4733 -1950 4750
rect -2157 4710 -1950 4733
rect -2157 4693 -2143 4710
rect -1968 4693 -1950 4710
rect -2157 4670 -1950 4693
rect -2157 4653 -2143 4670
rect -1968 4653 -1950 4670
rect -2157 4630 -1950 4653
rect -2157 4613 -2143 4630
rect -1968 4613 -1950 4630
rect -2157 4590 -1950 4613
rect -2157 4573 -2143 4590
rect -1968 4573 -1950 4590
rect -2157 4550 -1950 4573
rect -2157 4533 -2143 4550
rect -1968 4533 -1950 4550
rect -2157 4510 -1950 4533
rect -2157 4493 -2143 4510
rect -1968 4493 -1950 4510
rect -2157 4470 -1950 4493
rect -2157 4453 -2143 4470
rect -1968 4453 -1950 4470
rect -2157 4430 -1950 4453
rect -2157 4413 -2143 4430
rect -1968 4413 -1950 4430
rect -2157 4390 -1950 4413
rect -2157 4373 -2143 4390
rect -1968 4373 -1950 4390
rect -2157 4350 -1950 4373
rect -2157 4333 -2143 4350
rect -1968 4333 -1950 4350
rect -2157 4310 -1950 4333
rect -2157 4293 -2143 4310
rect -1968 4293 -1950 4310
rect -2157 4270 -1950 4293
rect -2157 4253 -2143 4270
rect -1968 4253 -1950 4270
rect -2157 4230 -1950 4253
rect -2157 4213 -2143 4230
rect -1968 4213 -1950 4230
rect -2157 4190 -1950 4213
rect -2157 4173 -2143 4190
rect -1968 4173 -1950 4190
rect -2157 4150 -1950 4173
rect -2157 4133 -2143 4150
rect -1968 4133 -1950 4150
rect -2157 4110 -1950 4133
rect -2157 4093 -2143 4110
rect -1968 4093 -1950 4110
rect -2157 4070 -1950 4093
rect -2157 4053 -2143 4070
rect -1968 4053 -1950 4070
rect -2157 4030 -1950 4053
rect -2157 4013 -2143 4030
rect -1968 4013 -1950 4030
rect -2157 3990 -1950 4013
rect -2157 3973 -2143 3990
rect -1968 3973 -1950 3990
rect -2157 3950 -1950 3973
rect -2157 3933 -2143 3950
rect -1968 3933 -1950 3950
rect -2157 3910 -1950 3933
rect -2157 3893 -2143 3910
rect -1968 3893 -1950 3910
rect -2157 3870 -1950 3893
rect -2157 3853 -2143 3870
rect -1968 3853 -1950 3870
rect -2157 3830 -1950 3853
rect -2157 3813 -2143 3830
rect -1968 3813 -1950 3830
rect -2157 3790 -1950 3813
rect -2157 3773 -2143 3790
rect -1968 3773 -1950 3790
rect -2157 3750 -1950 3773
rect -2157 3733 -2143 3750
rect -1968 3733 -1950 3750
rect -2157 3710 -1950 3733
rect -2157 3693 -2143 3710
rect -1968 3693 -1950 3710
rect -2157 3670 -1950 3693
rect -2157 3653 -2143 3670
rect -1968 3653 -1950 3670
rect -2157 3630 -1950 3653
rect -2157 3613 -2143 3630
rect -1968 3613 -1950 3630
rect -2157 3590 -1950 3613
rect -2157 3573 -2143 3590
rect -1968 3573 -1950 3590
rect -2157 3550 -1950 3573
rect -2157 3533 -2143 3550
rect -1968 3533 -1950 3550
rect -2157 3510 -1950 3533
rect -2157 3493 -2143 3510
rect -1968 3493 -1950 3510
rect -2157 3470 -1950 3493
rect -2157 3453 -2143 3470
rect -1968 3453 -1950 3470
rect -2157 3430 -1950 3453
rect -2157 3413 -2143 3430
rect -1968 3413 -1950 3430
rect -2157 3390 -1950 3413
rect -2157 3373 -2143 3390
rect -1968 3373 -1950 3390
rect -2157 3350 -1950 3373
rect -2157 3333 -2143 3350
rect -1968 3333 -1950 3350
rect -2157 3310 -1950 3333
rect -2157 3293 -2143 3310
rect -1968 3293 -1950 3310
rect -2157 3270 -1950 3293
rect -2157 3253 -2143 3270
rect -1968 3253 -1950 3270
rect -2157 3230 -1950 3253
rect -2157 3213 -2143 3230
rect -1968 3213 -1950 3230
rect -2157 3190 -1950 3213
rect -2157 3173 -2143 3190
rect -1968 3173 -1950 3190
rect -2157 3150 -1950 3173
rect -2157 3133 -2143 3150
rect -1968 3133 -1950 3150
rect -2157 3110 -1950 3133
rect -2157 3093 -2143 3110
rect -1968 3093 -1950 3110
rect -2157 3070 -1950 3093
rect -2157 3053 -2143 3070
rect -1968 3053 -1950 3070
rect -2157 3030 -1950 3053
rect -2157 3013 -2143 3030
rect -1968 3013 -1950 3030
rect -2157 2990 -1950 3013
rect -2157 2973 -2143 2990
rect -1968 2973 -1950 2990
rect -2157 2950 -1950 2973
rect -2157 2933 -2143 2950
rect -1968 2933 -1950 2950
rect -2157 2910 -1950 2933
rect -2157 2893 -2143 2910
rect -1968 2893 -1950 2910
rect -2157 2870 -1950 2893
rect -2157 2853 -2143 2870
rect -1968 2853 -1950 2870
rect -2157 2830 -1950 2853
rect -2157 2813 -2143 2830
rect -1968 2813 -1950 2830
rect -2157 2790 -1950 2813
rect -2157 2773 -2143 2790
rect -1968 2773 -1950 2790
rect -2157 2750 -1950 2773
rect -2157 2733 -2143 2750
rect -1968 2733 -1950 2750
rect -2157 2710 -1950 2733
rect -2157 2693 -2143 2710
rect -1968 2693 -1950 2710
rect -2157 2670 -1950 2693
rect -2157 2653 -2143 2670
rect -1968 2653 -1950 2670
rect -2157 2630 -1950 2653
rect -2157 2613 -2143 2630
rect -1968 2613 -1950 2630
rect -2157 2590 -1950 2613
rect -2157 2573 -2143 2590
rect -1968 2573 -1950 2590
rect -2157 2550 -1950 2573
rect -2157 2533 -2143 2550
rect -1968 2533 -1950 2550
rect -2157 2510 -1950 2533
rect -2157 2493 -2143 2510
rect -1968 2493 -1950 2510
rect -2157 2470 -1950 2493
rect -2157 2453 -2143 2470
rect -1968 2453 -1950 2470
rect -2157 2430 -1950 2453
rect -2157 2413 -2143 2430
rect -1968 2413 -1950 2430
rect -2157 2390 -1950 2413
rect -2157 2373 -2143 2390
rect -1968 2373 -1950 2390
rect -2157 2350 -1950 2373
rect -2157 2333 -2143 2350
rect -1968 2333 -1950 2350
rect -2157 2310 -1950 2333
rect -2157 2293 -2143 2310
rect -1968 2293 -1950 2310
rect -2157 2270 -1950 2293
rect -2157 2253 -2143 2270
rect -1968 2253 -1950 2270
rect -2157 2230 -1950 2253
rect -2157 2213 -2143 2230
rect -1968 2213 -1950 2230
rect -2157 2190 -1950 2213
rect -2157 2173 -2143 2190
rect -1968 2173 -1950 2190
rect -2157 2150 -1950 2173
rect -2157 2133 -2143 2150
rect -1968 2133 -1950 2150
rect -2157 2110 -1950 2133
rect -2157 2093 -2143 2110
rect -1968 2093 -1950 2110
rect -2157 2070 -1950 2093
rect -2157 2053 -2143 2070
rect -1968 2053 -1950 2070
rect -2157 2030 -1950 2053
rect -2157 2013 -2143 2030
rect -1968 2013 -1950 2030
rect -2157 1990 -1950 2013
rect -2157 1973 -2143 1990
rect -1968 1973 -1950 1990
rect -2157 1950 -1950 1973
rect -2157 1933 -2143 1950
rect -1968 1933 -1950 1950
rect -2157 1910 -1950 1933
rect -2157 1893 -2143 1910
rect -1968 1893 -1950 1910
rect -2157 1870 -1950 1893
rect -2157 1853 -2143 1870
rect -1968 1853 -1950 1870
rect -2157 1830 -1950 1853
rect -2157 1813 -2143 1830
rect -1968 1813 -1950 1830
rect -2157 1790 -1950 1813
rect -2157 1773 -2143 1790
rect -1968 1773 -1950 1790
rect -2157 1750 -1950 1773
rect -2157 1733 -2143 1750
rect -1968 1733 -1950 1750
rect -2157 1710 -1950 1733
rect -2157 1693 -2143 1710
rect -1968 1693 -1950 1710
rect -2157 1670 -1950 1693
rect -2157 1653 -2143 1670
rect -1968 1653 -1950 1670
rect -2157 1630 -1950 1653
rect -2157 1613 -2143 1630
rect -1968 1613 -1950 1630
rect -2157 1590 -1950 1613
rect -2157 1573 -2143 1590
rect -1968 1573 -1950 1590
rect -2157 1550 -1950 1573
rect -2157 1533 -2143 1550
rect -1968 1533 -1950 1550
rect -2157 1510 -1950 1533
rect -2157 1493 -2143 1510
rect -1968 1493 -1950 1510
rect -2157 1470 -1950 1493
rect -2157 1453 -2143 1470
rect -1968 1453 -1950 1470
rect -2157 1430 -1950 1453
rect -2157 1413 -2143 1430
rect -1968 1413 -1950 1430
rect -2157 1390 -1950 1413
rect -2157 1373 -2143 1390
rect -1968 1373 -1950 1390
rect -2157 1350 -1950 1373
rect -2157 1333 -2143 1350
rect -1968 1333 -1950 1350
rect -2157 1310 -1950 1333
rect -2157 1293 -2143 1310
rect -1968 1293 -1950 1310
rect -2157 1270 -1950 1293
rect -2157 1253 -2143 1270
rect -1968 1253 -1950 1270
rect -2157 1230 -1950 1253
rect -2157 1213 -2143 1230
rect -1968 1213 -1950 1230
rect -2157 1190 -1950 1213
rect -2157 1173 -2143 1190
rect -1968 1173 -1950 1190
rect -2157 1150 -1950 1173
rect -2157 1133 -2143 1150
rect -1968 1133 -1950 1150
rect -2157 1110 -1950 1133
rect -2157 1093 -2143 1110
rect -1968 1093 -1950 1110
rect -2157 1070 -1950 1093
rect -2157 1053 -2143 1070
rect -1968 1053 -1950 1070
rect -2157 1030 -1950 1053
rect -2157 1013 -2143 1030
rect -1968 1013 -1950 1030
rect -2157 990 -1950 1013
rect -2157 973 -2143 990
rect -1968 973 -1950 990
rect -2157 950 -1950 973
rect -2157 933 -2143 950
rect -1968 933 -1950 950
rect -2157 910 -1950 933
rect -2157 893 -2143 910
rect -1968 893 -1950 910
rect -2157 870 -1950 893
rect -2157 853 -2143 870
rect -1968 853 -1950 870
rect -2157 830 -1950 853
rect -2157 813 -2143 830
rect -1968 813 -1950 830
rect -2157 790 -1950 813
rect -2157 773 -2143 790
rect -1968 773 -1950 790
rect -2157 750 -1950 773
rect -2157 733 -2143 750
rect -1968 733 -1950 750
rect -2157 710 -1950 733
rect -2157 693 -2143 710
rect -1968 693 -1950 710
rect -2157 670 -1950 693
rect -2157 653 -2143 670
rect -1968 653 -1950 670
rect -2157 630 -1950 653
rect -2157 613 -2143 630
rect -1968 613 -1950 630
rect -2157 590 -1950 613
rect -2157 573 -2143 590
rect -1968 573 -1950 590
rect -2157 550 -1950 573
rect -2157 533 -2143 550
rect -1968 533 -1950 550
rect -2157 510 -1950 533
rect -2157 493 -2143 510
rect -1968 493 -1950 510
rect -2157 470 -1950 493
rect -2157 453 -2143 470
rect -1968 453 -1950 470
rect -2157 430 -1950 453
rect -2157 413 -2143 430
rect -1968 413 -1950 430
rect -2157 390 -1950 413
rect -2157 373 -2143 390
rect -1968 373 -1950 390
rect -2157 350 -1950 373
rect -2157 333 -2143 350
rect -1968 333 -1950 350
rect -2157 310 -1950 333
rect -2157 293 -2143 310
rect -1968 293 -1950 310
rect -2157 270 -1950 293
rect -2157 253 -2143 270
rect -1968 253 -1950 270
rect -2157 230 -1950 253
rect -2157 213 -2143 230
rect -1968 213 -1950 230
rect -2157 190 -1950 213
rect -2157 173 -2143 190
rect -1968 173 -1950 190
rect -2157 150 -1950 173
rect -2157 133 -2143 150
rect -1968 133 -1950 150
rect -2157 110 -1950 133
rect -2157 93 -2143 110
rect -1968 93 -1950 110
rect -2157 70 -1950 93
rect -2157 53 -2143 70
rect -1968 53 -1950 70
rect -2157 30 -1950 53
rect -2157 13 -2143 30
rect -1968 13 -1950 30
rect -2157 -217 -1950 13
rect 17694 9110 17901 9274
rect 17694 9093 17712 9110
rect 17887 9093 17901 9110
rect 17694 9070 17901 9093
rect 17694 9053 17712 9070
rect 17887 9053 17901 9070
rect 17694 9030 17901 9053
rect 17694 9013 17712 9030
rect 17887 9013 17901 9030
rect 17694 8990 17901 9013
rect 17694 8973 17712 8990
rect 17887 8973 17901 8990
rect 17694 8950 17901 8973
rect 17694 8933 17712 8950
rect 17887 8933 17901 8950
rect 17694 8910 17901 8933
rect 17694 8893 17712 8910
rect 17887 8893 17901 8910
rect 17694 8870 17901 8893
rect 17694 8853 17712 8870
rect 17887 8853 17901 8870
rect 17694 8830 17901 8853
rect 17694 8813 17712 8830
rect 17887 8813 17901 8830
rect 17694 8790 17901 8813
rect 17694 8773 17712 8790
rect 17887 8773 17901 8790
rect 17694 8750 17901 8773
rect 17694 8733 17712 8750
rect 17887 8733 17901 8750
rect 17694 8710 17901 8733
rect 17694 8693 17712 8710
rect 17887 8693 17901 8710
rect 17694 8670 17901 8693
rect 17694 8653 17712 8670
rect 17887 8653 17901 8670
rect 17694 8630 17901 8653
rect 17694 8613 17712 8630
rect 17887 8613 17901 8630
rect 17694 8590 17901 8613
rect 17694 8573 17712 8590
rect 17887 8573 17901 8590
rect 17694 8550 17901 8573
rect 17694 8533 17712 8550
rect 17887 8533 17901 8550
rect 17694 8510 17901 8533
rect 17694 8493 17712 8510
rect 17887 8493 17901 8510
rect 17694 8470 17901 8493
rect 17694 8453 17712 8470
rect 17887 8453 17901 8470
rect 17694 8430 17901 8453
rect 17694 8413 17712 8430
rect 17887 8413 17901 8430
rect 17694 8390 17901 8413
rect 17694 8373 17712 8390
rect 17887 8373 17901 8390
rect 17694 8350 17901 8373
rect 17694 8333 17712 8350
rect 17887 8333 17901 8350
rect 17694 8310 17901 8333
rect 17694 8293 17712 8310
rect 17887 8293 17901 8310
rect 17694 8270 17901 8293
rect 17694 8253 17712 8270
rect 17887 8253 17901 8270
rect 17694 8230 17901 8253
rect 17694 8213 17712 8230
rect 17887 8213 17901 8230
rect 17694 8190 17901 8213
rect 17694 8173 17712 8190
rect 17887 8173 17901 8190
rect 17694 8150 17901 8173
rect 17694 8133 17712 8150
rect 17887 8133 17901 8150
rect 17694 8110 17901 8133
rect 17694 8093 17712 8110
rect 17887 8093 17901 8110
rect 17694 8070 17901 8093
rect 17694 8053 17712 8070
rect 17887 8053 17901 8070
rect 17694 8030 17901 8053
rect 17694 8013 17712 8030
rect 17887 8013 17901 8030
rect 17694 7990 17901 8013
rect 17694 7973 17712 7990
rect 17887 7973 17901 7990
rect 17694 7950 17901 7973
rect 17694 7933 17712 7950
rect 17887 7933 17901 7950
rect 17694 7910 17901 7933
rect 17694 7893 17712 7910
rect 17887 7893 17901 7910
rect 17694 7870 17901 7893
rect 17694 7853 17712 7870
rect 17887 7853 17901 7870
rect 17694 7830 17901 7853
rect 17694 7813 17712 7830
rect 17887 7813 17901 7830
rect 17694 7790 17901 7813
rect 17694 7773 17712 7790
rect 17887 7773 17901 7790
rect 17694 7750 17901 7773
rect 17694 7733 17712 7750
rect 17887 7733 17901 7750
rect 17694 7710 17901 7733
rect 17694 7693 17712 7710
rect 17887 7693 17901 7710
rect 17694 7670 17901 7693
rect 17694 7653 17712 7670
rect 17887 7653 17901 7670
rect 17694 7630 17901 7653
rect 17694 7613 17712 7630
rect 17887 7613 17901 7630
rect 17694 7590 17901 7613
rect 17694 7573 17712 7590
rect 17887 7573 17901 7590
rect 17694 7550 17901 7573
rect 17694 7533 17712 7550
rect 17887 7533 17901 7550
rect 17694 7510 17901 7533
rect 17694 7493 17712 7510
rect 17887 7493 17901 7510
rect 17694 7470 17901 7493
rect 17694 7453 17712 7470
rect 17887 7453 17901 7470
rect 17694 7430 17901 7453
rect 17694 7413 17712 7430
rect 17887 7413 17901 7430
rect 17694 7390 17901 7413
rect 17694 7373 17712 7390
rect 17887 7373 17901 7390
rect 17694 7350 17901 7373
rect 17694 7333 17712 7350
rect 17887 7333 17901 7350
rect 17694 7310 17901 7333
rect 17694 7293 17712 7310
rect 17887 7293 17901 7310
rect 17694 7270 17901 7293
rect 17694 7253 17712 7270
rect 17887 7253 17901 7270
rect 17694 7230 17901 7253
rect 17694 7213 17712 7230
rect 17887 7213 17901 7230
rect 17694 7190 17901 7213
rect 17694 7173 17712 7190
rect 17887 7173 17901 7190
rect 17694 7150 17901 7173
rect 17694 7133 17712 7150
rect 17887 7133 17901 7150
rect 17694 7110 17901 7133
rect 17694 7093 17712 7110
rect 17887 7093 17901 7110
rect 17694 7070 17901 7093
rect 17694 7053 17712 7070
rect 17887 7053 17901 7070
rect 17694 7030 17901 7053
rect 17694 7013 17712 7030
rect 17887 7013 17901 7030
rect 17694 6990 17901 7013
rect 17694 6973 17712 6990
rect 17887 6973 17901 6990
rect 17694 6950 17901 6973
rect 17694 6933 17712 6950
rect 17887 6933 17901 6950
rect 17694 6910 17901 6933
rect 17694 6893 17712 6910
rect 17887 6893 17901 6910
rect 17694 6870 17901 6893
rect 17694 6853 17712 6870
rect 17887 6853 17901 6870
rect 17694 6830 17901 6853
rect 17694 6813 17712 6830
rect 17887 6813 17901 6830
rect 17694 6790 17901 6813
rect 17694 6773 17712 6790
rect 17887 6773 17901 6790
rect 17694 6750 17901 6773
rect 17694 6733 17712 6750
rect 17887 6733 17901 6750
rect 17694 6710 17901 6733
rect 17694 6693 17712 6710
rect 17887 6693 17901 6710
rect 17694 6670 17901 6693
rect 17694 6653 17712 6670
rect 17887 6653 17901 6670
rect 17694 6630 17901 6653
rect 17694 6613 17712 6630
rect 17887 6613 17901 6630
rect 17694 6590 17901 6613
rect 17694 6573 17712 6590
rect 17887 6573 17901 6590
rect 17694 6550 17901 6573
rect 17694 6533 17712 6550
rect 17887 6533 17901 6550
rect 17694 6510 17901 6533
rect 17694 6493 17712 6510
rect 17887 6493 17901 6510
rect 17694 6470 17901 6493
rect 17694 6453 17712 6470
rect 17887 6453 17901 6470
rect 17694 6430 17901 6453
rect 17694 6413 17712 6430
rect 17887 6413 17901 6430
rect 17694 6390 17901 6413
rect 17694 6373 17712 6390
rect 17887 6373 17901 6390
rect 17694 6350 17901 6373
rect 17694 6333 17712 6350
rect 17887 6333 17901 6350
rect 17694 6310 17901 6333
rect 17694 6293 17712 6310
rect 17887 6293 17901 6310
rect 17694 6270 17901 6293
rect 17694 6253 17712 6270
rect 17887 6253 17901 6270
rect 17694 6230 17901 6253
rect 17694 6213 17712 6230
rect 17887 6213 17901 6230
rect 17694 6190 17901 6213
rect 17694 6173 17712 6190
rect 17887 6173 17901 6190
rect 17694 6150 17901 6173
rect 17694 6133 17712 6150
rect 17887 6133 17901 6150
rect 17694 6110 17901 6133
rect 17694 6093 17712 6110
rect 17887 6093 17901 6110
rect 17694 6070 17901 6093
rect 17694 6053 17712 6070
rect 17887 6053 17901 6070
rect 17694 6030 17901 6053
rect 17694 6013 17712 6030
rect 17887 6013 17901 6030
rect 17694 5990 17901 6013
rect 17694 5973 17712 5990
rect 17887 5973 17901 5990
rect 17694 5950 17901 5973
rect 17694 5933 17712 5950
rect 17887 5933 17901 5950
rect 17694 5910 17901 5933
rect 17694 5893 17712 5910
rect 17887 5893 17901 5910
rect 17694 5870 17901 5893
rect 17694 5853 17712 5870
rect 17887 5853 17901 5870
rect 17694 5830 17901 5853
rect 17694 5813 17712 5830
rect 17887 5813 17901 5830
rect 17694 5790 17901 5813
rect 17694 5773 17712 5790
rect 17887 5773 17901 5790
rect 17694 5750 17901 5773
rect 17694 5733 17712 5750
rect 17887 5733 17901 5750
rect 17694 5710 17901 5733
rect 17694 5693 17712 5710
rect 17887 5693 17901 5710
rect 17694 5670 17901 5693
rect 17694 5653 17712 5670
rect 17887 5653 17901 5670
rect 17694 5630 17901 5653
rect 17694 5613 17712 5630
rect 17887 5613 17901 5630
rect 17694 5590 17901 5613
rect 17694 5573 17712 5590
rect 17887 5573 17901 5590
rect 17694 5550 17901 5573
rect 17694 5533 17712 5550
rect 17887 5533 17901 5550
rect 17694 5510 17901 5533
rect 17694 5493 17712 5510
rect 17887 5493 17901 5510
rect 17694 5470 17901 5493
rect 17694 5453 17712 5470
rect 17887 5453 17901 5470
rect 17694 5430 17901 5453
rect 17694 5413 17712 5430
rect 17887 5413 17901 5430
rect 17694 5390 17901 5413
rect 17694 5373 17712 5390
rect 17887 5373 17901 5390
rect 17694 5350 17901 5373
rect 17694 5333 17712 5350
rect 17887 5333 17901 5350
rect 17694 5310 17901 5333
rect 17694 5293 17712 5310
rect 17887 5293 17901 5310
rect 17694 5270 17901 5293
rect 17694 5253 17712 5270
rect 17887 5253 17901 5270
rect 17694 5230 17901 5253
rect 17694 5213 17712 5230
rect 17887 5213 17901 5230
rect 17694 5190 17901 5213
rect 17694 5173 17712 5190
rect 17887 5173 17901 5190
rect 17694 5150 17901 5173
rect 17694 5133 17712 5150
rect 17887 5133 17901 5150
rect 17694 5110 17901 5133
rect 17694 5093 17712 5110
rect 17887 5093 17901 5110
rect 17694 5070 17901 5093
rect 17694 5053 17712 5070
rect 17887 5053 17901 5070
rect 17694 5030 17901 5053
rect 17694 5013 17712 5030
rect 17887 5013 17901 5030
rect 17694 4990 17901 5013
rect 17694 4973 17712 4990
rect 17887 4973 17901 4990
rect 17694 4950 17901 4973
rect 17694 4933 17712 4950
rect 17887 4933 17901 4950
rect 17694 4910 17901 4933
rect 17694 4893 17712 4910
rect 17887 4893 17901 4910
rect 17694 4870 17901 4893
rect 17694 4853 17712 4870
rect 17887 4853 17901 4870
rect 17694 4830 17901 4853
rect 17694 4813 17712 4830
rect 17887 4813 17901 4830
rect 17694 4790 17901 4813
rect 17694 4773 17712 4790
rect 17887 4773 17901 4790
rect 17694 4750 17901 4773
rect 17694 4733 17712 4750
rect 17887 4733 17901 4750
rect 17694 4710 17901 4733
rect 17694 4693 17712 4710
rect 17887 4693 17901 4710
rect 17694 4670 17901 4693
rect 17694 4653 17712 4670
rect 17887 4653 17901 4670
rect 17694 4630 17901 4653
rect 17694 4613 17712 4630
rect 17887 4613 17901 4630
rect 17694 4590 17901 4613
rect 17694 4573 17712 4590
rect 17887 4573 17901 4590
rect 17694 4550 17901 4573
rect 17694 4533 17712 4550
rect 17887 4533 17901 4550
rect 17694 4510 17901 4533
rect 17694 4493 17712 4510
rect 17887 4493 17901 4510
rect 17694 4470 17901 4493
rect 17694 4453 17712 4470
rect 17887 4453 17901 4470
rect 17694 4430 17901 4453
rect 17694 4413 17712 4430
rect 17887 4413 17901 4430
rect 17694 4390 17901 4413
rect 17694 4373 17712 4390
rect 17887 4373 17901 4390
rect 17694 4350 17901 4373
rect 17694 4333 17712 4350
rect 17887 4333 17901 4350
rect 17694 4310 17901 4333
rect 17694 4293 17712 4310
rect 17887 4293 17901 4310
rect 17694 4270 17901 4293
rect 17694 4253 17712 4270
rect 17887 4253 17901 4270
rect 17694 4230 17901 4253
rect 17694 4213 17712 4230
rect 17887 4213 17901 4230
rect 17694 4190 17901 4213
rect 17694 4173 17712 4190
rect 17887 4173 17901 4190
rect 17694 4150 17901 4173
rect 17694 4133 17712 4150
rect 17887 4133 17901 4150
rect 17694 4110 17901 4133
rect 17694 4093 17712 4110
rect 17887 4093 17901 4110
rect 17694 4070 17901 4093
rect 17694 4053 17712 4070
rect 17887 4053 17901 4070
rect 17694 4030 17901 4053
rect 17694 4013 17712 4030
rect 17887 4013 17901 4030
rect 17694 3990 17901 4013
rect 17694 3973 17712 3990
rect 17887 3973 17901 3990
rect 17694 3950 17901 3973
rect 17694 3933 17712 3950
rect 17887 3933 17901 3950
rect 17694 3910 17901 3933
rect 17694 3893 17712 3910
rect 17887 3893 17901 3910
rect 17694 3870 17901 3893
rect 17694 3853 17712 3870
rect 17887 3853 17901 3870
rect 17694 3830 17901 3853
rect 17694 3813 17712 3830
rect 17887 3813 17901 3830
rect 17694 3790 17901 3813
rect 17694 3773 17712 3790
rect 17887 3773 17901 3790
rect 17694 3750 17901 3773
rect 17694 3733 17712 3750
rect 17887 3733 17901 3750
rect 17694 3710 17901 3733
rect 17694 3693 17712 3710
rect 17887 3693 17901 3710
rect 17694 3670 17901 3693
rect 17694 3653 17712 3670
rect 17887 3653 17901 3670
rect 17694 3630 17901 3653
rect 17694 3613 17712 3630
rect 17887 3613 17901 3630
rect 17694 3590 17901 3613
rect 17694 3573 17712 3590
rect 17887 3573 17901 3590
rect 17694 3550 17901 3573
rect 17694 3533 17712 3550
rect 17887 3533 17901 3550
rect 17694 3510 17901 3533
rect 17694 3493 17712 3510
rect 17887 3493 17901 3510
rect 17694 3470 17901 3493
rect 17694 3453 17712 3470
rect 17887 3453 17901 3470
rect 17694 3430 17901 3453
rect 17694 3413 17712 3430
rect 17887 3413 17901 3430
rect 17694 3390 17901 3413
rect 17694 3373 17712 3390
rect 17887 3373 17901 3390
rect 17694 3350 17901 3373
rect 17694 3333 17712 3350
rect 17887 3333 17901 3350
rect 17694 3310 17901 3333
rect 17694 3293 17712 3310
rect 17887 3293 17901 3310
rect 17694 3270 17901 3293
rect 17694 3253 17712 3270
rect 17887 3253 17901 3270
rect 17694 3230 17901 3253
rect 17694 3213 17712 3230
rect 17887 3213 17901 3230
rect 17694 3190 17901 3213
rect 17694 3173 17712 3190
rect 17887 3173 17901 3190
rect 17694 3150 17901 3173
rect 17694 3133 17712 3150
rect 17887 3133 17901 3150
rect 17694 3110 17901 3133
rect 17694 3093 17712 3110
rect 17887 3093 17901 3110
rect 17694 3070 17901 3093
rect 17694 3053 17712 3070
rect 17887 3053 17901 3070
rect 17694 3030 17901 3053
rect 17694 3013 17712 3030
rect 17887 3013 17901 3030
rect 17694 2990 17901 3013
rect 17694 2973 17712 2990
rect 17887 2973 17901 2990
rect 17694 2950 17901 2973
rect 17694 2933 17712 2950
rect 17887 2933 17901 2950
rect 17694 2910 17901 2933
rect 17694 2893 17712 2910
rect 17887 2893 17901 2910
rect 17694 2870 17901 2893
rect 17694 2853 17712 2870
rect 17887 2853 17901 2870
rect 17694 2830 17901 2853
rect 17694 2813 17712 2830
rect 17887 2813 17901 2830
rect 17694 2790 17901 2813
rect 17694 2773 17712 2790
rect 17887 2773 17901 2790
rect 17694 2750 17901 2773
rect 17694 2733 17712 2750
rect 17887 2733 17901 2750
rect 17694 2710 17901 2733
rect 17694 2693 17712 2710
rect 17887 2693 17901 2710
rect 17694 2670 17901 2693
rect 17694 2653 17712 2670
rect 17887 2653 17901 2670
rect 17694 2630 17901 2653
rect 17694 2613 17712 2630
rect 17887 2613 17901 2630
rect 17694 2590 17901 2613
rect 17694 2573 17712 2590
rect 17887 2573 17901 2590
rect 17694 2550 17901 2573
rect 17694 2533 17712 2550
rect 17887 2533 17901 2550
rect 17694 2510 17901 2533
rect 17694 2493 17712 2510
rect 17887 2493 17901 2510
rect 17694 2470 17901 2493
rect 17694 2453 17712 2470
rect 17887 2453 17901 2470
rect 17694 2430 17901 2453
rect 17694 2413 17712 2430
rect 17887 2413 17901 2430
rect 17694 2390 17901 2413
rect 17694 2373 17712 2390
rect 17887 2373 17901 2390
rect 17694 2350 17901 2373
rect 17694 2333 17712 2350
rect 17887 2333 17901 2350
rect 17694 2310 17901 2333
rect 17694 2293 17712 2310
rect 17887 2293 17901 2310
rect 17694 2270 17901 2293
rect 17694 2253 17712 2270
rect 17887 2253 17901 2270
rect 17694 2230 17901 2253
rect 17694 2213 17712 2230
rect 17887 2213 17901 2230
rect 17694 2190 17901 2213
rect 17694 2173 17712 2190
rect 17887 2173 17901 2190
rect 17694 2150 17901 2173
rect 17694 2133 17712 2150
rect 17887 2133 17901 2150
rect 17694 2110 17901 2133
rect 17694 2093 17712 2110
rect 17887 2093 17901 2110
rect 17694 2070 17901 2093
rect 17694 2053 17712 2070
rect 17887 2053 17901 2070
rect 17694 2030 17901 2053
rect 17694 2013 17712 2030
rect 17887 2013 17901 2030
rect 17694 1990 17901 2013
rect 17694 1973 17712 1990
rect 17887 1973 17901 1990
rect 17694 1950 17901 1973
rect 17694 1933 17712 1950
rect 17887 1933 17901 1950
rect 17694 1910 17901 1933
rect 17694 1893 17712 1910
rect 17887 1893 17901 1910
rect 17694 1870 17901 1893
rect 17694 1853 17712 1870
rect 17887 1853 17901 1870
rect 17694 1830 17901 1853
rect 17694 1813 17712 1830
rect 17887 1813 17901 1830
rect 17694 1790 17901 1813
rect 17694 1773 17712 1790
rect 17887 1773 17901 1790
rect 17694 1750 17901 1773
rect 17694 1733 17712 1750
rect 17887 1733 17901 1750
rect 17694 1710 17901 1733
rect 17694 1693 17712 1710
rect 17887 1693 17901 1710
rect 17694 1670 17901 1693
rect 17694 1653 17712 1670
rect 17887 1653 17901 1670
rect 17694 1630 17901 1653
rect 17694 1613 17712 1630
rect 17887 1613 17901 1630
rect 17694 1590 17901 1613
rect 17694 1573 17712 1590
rect 17887 1573 17901 1590
rect 17694 1550 17901 1573
rect 17694 1533 17712 1550
rect 17887 1533 17901 1550
rect 17694 1510 17901 1533
rect 17694 1493 17712 1510
rect 17887 1493 17901 1510
rect 17694 1470 17901 1493
rect 17694 1453 17712 1470
rect 17887 1453 17901 1470
rect 17694 1430 17901 1453
rect 17694 1413 17712 1430
rect 17887 1413 17901 1430
rect 17694 1390 17901 1413
rect 17694 1373 17712 1390
rect 17887 1373 17901 1390
rect 17694 1350 17901 1373
rect 17694 1333 17712 1350
rect 17887 1333 17901 1350
rect 17694 1310 17901 1333
rect 17694 1293 17712 1310
rect 17887 1293 17901 1310
rect 17694 1270 17901 1293
rect 17694 1253 17712 1270
rect 17887 1253 17901 1270
rect 17694 1230 17901 1253
rect 17694 1213 17712 1230
rect 17887 1213 17901 1230
rect 17694 1190 17901 1213
rect 17694 1173 17712 1190
rect 17887 1173 17901 1190
rect 17694 1150 17901 1173
rect 17694 1133 17712 1150
rect 17887 1133 17901 1150
rect 17694 1110 17901 1133
rect 17694 1093 17712 1110
rect 17887 1093 17901 1110
rect 17694 1070 17901 1093
rect 17694 1053 17712 1070
rect 17887 1053 17901 1070
rect 17694 1030 17901 1053
rect 17694 1013 17712 1030
rect 17887 1013 17901 1030
rect 17694 990 17901 1013
rect 17694 973 17712 990
rect 17887 973 17901 990
rect 17694 950 17901 973
rect 17694 933 17712 950
rect 17887 933 17901 950
rect 17694 910 17901 933
rect 17694 893 17712 910
rect 17887 893 17901 910
rect 17694 870 17901 893
rect 17694 853 17712 870
rect 17887 853 17901 870
rect 17694 830 17901 853
rect 17694 813 17712 830
rect 17887 813 17901 830
rect 17694 790 17901 813
rect 17694 773 17712 790
rect 17887 773 17901 790
rect 17694 750 17901 773
rect 17694 733 17712 750
rect 17887 733 17901 750
rect 17694 710 17901 733
rect 17694 693 17712 710
rect 17887 693 17901 710
rect 17694 670 17901 693
rect 17694 653 17712 670
rect 17887 653 17901 670
rect 17694 630 17901 653
rect 17694 613 17712 630
rect 17887 613 17901 630
rect 17694 590 17901 613
rect 17694 573 17712 590
rect 17887 573 17901 590
rect 17694 550 17901 573
rect 17694 533 17712 550
rect 17887 533 17901 550
rect 17694 510 17901 533
rect 17694 493 17712 510
rect 17887 493 17901 510
rect 17694 470 17901 493
rect 17694 453 17712 470
rect 17887 453 17901 470
rect 17694 430 17901 453
rect 17694 413 17712 430
rect 17887 413 17901 430
rect 17694 390 17901 413
rect 17694 373 17712 390
rect 17887 373 17901 390
rect 17694 350 17901 373
rect 17694 333 17712 350
rect 17887 333 17901 350
rect 17694 310 17901 333
rect 17694 293 17712 310
rect 17887 293 17901 310
rect 17694 270 17901 293
rect 17694 253 17712 270
rect 17887 253 17901 270
rect 17694 230 17901 253
rect 17694 213 17712 230
rect 17887 213 17901 230
rect 17694 190 17901 213
rect 17694 173 17712 190
rect 17887 173 17901 190
rect 17694 150 17901 173
rect 17694 133 17712 150
rect 17887 133 17901 150
rect 17694 110 17901 133
rect 17694 93 17712 110
rect 17887 93 17901 110
rect 17694 70 17901 93
rect 17694 53 17712 70
rect 17887 53 17901 70
rect 17694 30 17901 53
rect 17694 13 17712 30
rect 17887 13 17901 30
rect 17694 -152 17901 13
<< psubdiffcont >>
rect -2143 9093 -1968 9110
rect -2143 9053 -1968 9070
rect -2143 9013 -1968 9030
rect -2143 8973 -1968 8990
rect -2143 8933 -1968 8950
rect -2143 8893 -1968 8910
rect -2143 8853 -1968 8870
rect -2143 8813 -1968 8830
rect -2143 8773 -1968 8790
rect -2143 8733 -1968 8750
rect -2143 8693 -1968 8710
rect -2143 8653 -1968 8670
rect -2143 8613 -1968 8630
rect -2143 8573 -1968 8590
rect -2143 8533 -1968 8550
rect -2143 8493 -1968 8510
rect -2143 8453 -1968 8470
rect -2143 8413 -1968 8430
rect -2143 8373 -1968 8390
rect -2143 8333 -1968 8350
rect -2143 8293 -1968 8310
rect -2143 8253 -1968 8270
rect -2143 8213 -1968 8230
rect -2143 8173 -1968 8190
rect -2143 8133 -1968 8150
rect -2143 8093 -1968 8110
rect -2143 8053 -1968 8070
rect -2143 8013 -1968 8030
rect -2143 7973 -1968 7990
rect -2143 7933 -1968 7950
rect -2143 7893 -1968 7910
rect -2143 7853 -1968 7870
rect -2143 7813 -1968 7830
rect -2143 7773 -1968 7790
rect -2143 7733 -1968 7750
rect -2143 7693 -1968 7710
rect -2143 7653 -1968 7670
rect -2143 7613 -1968 7630
rect -2143 7573 -1968 7590
rect -2143 7533 -1968 7550
rect -2143 7493 -1968 7510
rect -2143 7453 -1968 7470
rect -2143 7413 -1968 7430
rect -2143 7373 -1968 7390
rect -2143 7333 -1968 7350
rect -2143 7293 -1968 7310
rect -2143 7253 -1968 7270
rect -2143 7213 -1968 7230
rect -2143 7173 -1968 7190
rect -2143 7133 -1968 7150
rect -2143 7093 -1968 7110
rect -2143 7053 -1968 7070
rect -2143 7013 -1968 7030
rect -2143 6973 -1968 6990
rect -2143 6933 -1968 6950
rect -2143 6893 -1968 6910
rect -2143 6853 -1968 6870
rect -2143 6813 -1968 6830
rect -2143 6773 -1968 6790
rect -2143 6733 -1968 6750
rect -2143 6693 -1968 6710
rect -2143 6653 -1968 6670
rect -2143 6613 -1968 6630
rect -2143 6573 -1968 6590
rect -2143 6533 -1968 6550
rect -2143 6493 -1968 6510
rect -2143 6453 -1968 6470
rect -2143 6413 -1968 6430
rect -2143 6373 -1968 6390
rect -2143 6333 -1968 6350
rect -2143 6293 -1968 6310
rect -2143 6253 -1968 6270
rect -2143 6213 -1968 6230
rect -2143 6173 -1968 6190
rect -2143 6133 -1968 6150
rect -2143 6093 -1968 6110
rect -2143 6053 -1968 6070
rect -2143 6013 -1968 6030
rect -2143 5973 -1968 5990
rect -2143 5933 -1968 5950
rect -2143 5893 -1968 5910
rect -2143 5853 -1968 5870
rect -2143 5813 -1968 5830
rect -2143 5773 -1968 5790
rect -2143 5733 -1968 5750
rect -2143 5693 -1968 5710
rect -2143 5653 -1968 5670
rect -2143 5613 -1968 5630
rect -2143 5573 -1968 5590
rect -2143 5533 -1968 5550
rect -2143 5493 -1968 5510
rect -2143 5453 -1968 5470
rect -2143 5413 -1968 5430
rect -2143 5373 -1968 5390
rect -2143 5333 -1968 5350
rect -2143 5293 -1968 5310
rect -2143 5253 -1968 5270
rect -2143 5213 -1968 5230
rect -2143 5173 -1968 5190
rect -2143 5133 -1968 5150
rect -2143 5093 -1968 5110
rect -2143 5053 -1968 5070
rect -2143 5013 -1968 5030
rect -2143 4973 -1968 4990
rect -2143 4933 -1968 4950
rect -2143 4893 -1968 4910
rect -2143 4853 -1968 4870
rect -2143 4813 -1968 4830
rect -2143 4773 -1968 4790
rect -2143 4733 -1968 4750
rect -2143 4693 -1968 4710
rect -2143 4653 -1968 4670
rect -2143 4613 -1968 4630
rect -2143 4573 -1968 4590
rect -2143 4533 -1968 4550
rect -2143 4493 -1968 4510
rect -2143 4453 -1968 4470
rect -2143 4413 -1968 4430
rect -2143 4373 -1968 4390
rect -2143 4333 -1968 4350
rect -2143 4293 -1968 4310
rect -2143 4253 -1968 4270
rect -2143 4213 -1968 4230
rect -2143 4173 -1968 4190
rect -2143 4133 -1968 4150
rect -2143 4093 -1968 4110
rect -2143 4053 -1968 4070
rect -2143 4013 -1968 4030
rect -2143 3973 -1968 3990
rect -2143 3933 -1968 3950
rect -2143 3893 -1968 3910
rect -2143 3853 -1968 3870
rect -2143 3813 -1968 3830
rect -2143 3773 -1968 3790
rect -2143 3733 -1968 3750
rect -2143 3693 -1968 3710
rect -2143 3653 -1968 3670
rect -2143 3613 -1968 3630
rect -2143 3573 -1968 3590
rect -2143 3533 -1968 3550
rect -2143 3493 -1968 3510
rect -2143 3453 -1968 3470
rect -2143 3413 -1968 3430
rect -2143 3373 -1968 3390
rect -2143 3333 -1968 3350
rect -2143 3293 -1968 3310
rect -2143 3253 -1968 3270
rect -2143 3213 -1968 3230
rect -2143 3173 -1968 3190
rect -2143 3133 -1968 3150
rect -2143 3093 -1968 3110
rect -2143 3053 -1968 3070
rect -2143 3013 -1968 3030
rect -2143 2973 -1968 2990
rect -2143 2933 -1968 2950
rect -2143 2893 -1968 2910
rect -2143 2853 -1968 2870
rect -2143 2813 -1968 2830
rect -2143 2773 -1968 2790
rect -2143 2733 -1968 2750
rect -2143 2693 -1968 2710
rect -2143 2653 -1968 2670
rect -2143 2613 -1968 2630
rect -2143 2573 -1968 2590
rect -2143 2533 -1968 2550
rect -2143 2493 -1968 2510
rect -2143 2453 -1968 2470
rect -2143 2413 -1968 2430
rect -2143 2373 -1968 2390
rect -2143 2333 -1968 2350
rect -2143 2293 -1968 2310
rect -2143 2253 -1968 2270
rect -2143 2213 -1968 2230
rect -2143 2173 -1968 2190
rect -2143 2133 -1968 2150
rect -2143 2093 -1968 2110
rect -2143 2053 -1968 2070
rect -2143 2013 -1968 2030
rect -2143 1973 -1968 1990
rect -2143 1933 -1968 1950
rect -2143 1893 -1968 1910
rect -2143 1853 -1968 1870
rect -2143 1813 -1968 1830
rect -2143 1773 -1968 1790
rect -2143 1733 -1968 1750
rect -2143 1693 -1968 1710
rect -2143 1653 -1968 1670
rect -2143 1613 -1968 1630
rect -2143 1573 -1968 1590
rect -2143 1533 -1968 1550
rect -2143 1493 -1968 1510
rect -2143 1453 -1968 1470
rect -2143 1413 -1968 1430
rect -2143 1373 -1968 1390
rect -2143 1333 -1968 1350
rect -2143 1293 -1968 1310
rect -2143 1253 -1968 1270
rect -2143 1213 -1968 1230
rect -2143 1173 -1968 1190
rect -2143 1133 -1968 1150
rect -2143 1093 -1968 1110
rect -2143 1053 -1968 1070
rect -2143 1013 -1968 1030
rect -2143 973 -1968 990
rect -2143 933 -1968 950
rect -2143 893 -1968 910
rect -2143 853 -1968 870
rect -2143 813 -1968 830
rect -2143 773 -1968 790
rect -2143 733 -1968 750
rect -2143 693 -1968 710
rect -2143 653 -1968 670
rect -2143 613 -1968 630
rect -2143 573 -1968 590
rect -2143 533 -1968 550
rect -2143 493 -1968 510
rect -2143 453 -1968 470
rect -2143 413 -1968 430
rect -2143 373 -1968 390
rect -2143 333 -1968 350
rect -2143 293 -1968 310
rect -2143 253 -1968 270
rect -2143 213 -1968 230
rect -2143 173 -1968 190
rect -2143 133 -1968 150
rect -2143 93 -1968 110
rect -2143 53 -1968 70
rect -2143 13 -1968 30
rect 17712 9093 17887 9110
rect 17712 9053 17887 9070
rect 17712 9013 17887 9030
rect 17712 8973 17887 8990
rect 17712 8933 17887 8950
rect 17712 8893 17887 8910
rect 17712 8853 17887 8870
rect 17712 8813 17887 8830
rect 17712 8773 17887 8790
rect 17712 8733 17887 8750
rect 17712 8693 17887 8710
rect 17712 8653 17887 8670
rect 17712 8613 17887 8630
rect 17712 8573 17887 8590
rect 17712 8533 17887 8550
rect 17712 8493 17887 8510
rect 17712 8453 17887 8470
rect 17712 8413 17887 8430
rect 17712 8373 17887 8390
rect 17712 8333 17887 8350
rect 17712 8293 17887 8310
rect 17712 8253 17887 8270
rect 17712 8213 17887 8230
rect 17712 8173 17887 8190
rect 17712 8133 17887 8150
rect 17712 8093 17887 8110
rect 17712 8053 17887 8070
rect 17712 8013 17887 8030
rect 17712 7973 17887 7990
rect 17712 7933 17887 7950
rect 17712 7893 17887 7910
rect 17712 7853 17887 7870
rect 17712 7813 17887 7830
rect 17712 7773 17887 7790
rect 17712 7733 17887 7750
rect 17712 7693 17887 7710
rect 17712 7653 17887 7670
rect 17712 7613 17887 7630
rect 17712 7573 17887 7590
rect 17712 7533 17887 7550
rect 17712 7493 17887 7510
rect 17712 7453 17887 7470
rect 17712 7413 17887 7430
rect 17712 7373 17887 7390
rect 17712 7333 17887 7350
rect 17712 7293 17887 7310
rect 17712 7253 17887 7270
rect 17712 7213 17887 7230
rect 17712 7173 17887 7190
rect 17712 7133 17887 7150
rect 17712 7093 17887 7110
rect 17712 7053 17887 7070
rect 17712 7013 17887 7030
rect 17712 6973 17887 6990
rect 17712 6933 17887 6950
rect 17712 6893 17887 6910
rect 17712 6853 17887 6870
rect 17712 6813 17887 6830
rect 17712 6773 17887 6790
rect 17712 6733 17887 6750
rect 17712 6693 17887 6710
rect 17712 6653 17887 6670
rect 17712 6613 17887 6630
rect 17712 6573 17887 6590
rect 17712 6533 17887 6550
rect 17712 6493 17887 6510
rect 17712 6453 17887 6470
rect 17712 6413 17887 6430
rect 17712 6373 17887 6390
rect 17712 6333 17887 6350
rect 17712 6293 17887 6310
rect 17712 6253 17887 6270
rect 17712 6213 17887 6230
rect 17712 6173 17887 6190
rect 17712 6133 17887 6150
rect 17712 6093 17887 6110
rect 17712 6053 17887 6070
rect 17712 6013 17887 6030
rect 17712 5973 17887 5990
rect 17712 5933 17887 5950
rect 17712 5893 17887 5910
rect 17712 5853 17887 5870
rect 17712 5813 17887 5830
rect 17712 5773 17887 5790
rect 17712 5733 17887 5750
rect 17712 5693 17887 5710
rect 17712 5653 17887 5670
rect 17712 5613 17887 5630
rect 17712 5573 17887 5590
rect 17712 5533 17887 5550
rect 17712 5493 17887 5510
rect 17712 5453 17887 5470
rect 17712 5413 17887 5430
rect 17712 5373 17887 5390
rect 17712 5333 17887 5350
rect 17712 5293 17887 5310
rect 17712 5253 17887 5270
rect 17712 5213 17887 5230
rect 17712 5173 17887 5190
rect 17712 5133 17887 5150
rect 17712 5093 17887 5110
rect 17712 5053 17887 5070
rect 17712 5013 17887 5030
rect 17712 4973 17887 4990
rect 17712 4933 17887 4950
rect 17712 4893 17887 4910
rect 17712 4853 17887 4870
rect 17712 4813 17887 4830
rect 17712 4773 17887 4790
rect 17712 4733 17887 4750
rect 17712 4693 17887 4710
rect 17712 4653 17887 4670
rect 17712 4613 17887 4630
rect 17712 4573 17887 4590
rect 17712 4533 17887 4550
rect 17712 4493 17887 4510
rect 17712 4453 17887 4470
rect 17712 4413 17887 4430
rect 17712 4373 17887 4390
rect 17712 4333 17887 4350
rect 17712 4293 17887 4310
rect 17712 4253 17887 4270
rect 17712 4213 17887 4230
rect 17712 4173 17887 4190
rect 17712 4133 17887 4150
rect 17712 4093 17887 4110
rect 17712 4053 17887 4070
rect 17712 4013 17887 4030
rect 17712 3973 17887 3990
rect 17712 3933 17887 3950
rect 17712 3893 17887 3910
rect 17712 3853 17887 3870
rect 17712 3813 17887 3830
rect 17712 3773 17887 3790
rect 17712 3733 17887 3750
rect 17712 3693 17887 3710
rect 17712 3653 17887 3670
rect 17712 3613 17887 3630
rect 17712 3573 17887 3590
rect 17712 3533 17887 3550
rect 17712 3493 17887 3510
rect 17712 3453 17887 3470
rect 17712 3413 17887 3430
rect 17712 3373 17887 3390
rect 17712 3333 17887 3350
rect 17712 3293 17887 3310
rect 17712 3253 17887 3270
rect 17712 3213 17887 3230
rect 17712 3173 17887 3190
rect 17712 3133 17887 3150
rect 17712 3093 17887 3110
rect 17712 3053 17887 3070
rect 17712 3013 17887 3030
rect 17712 2973 17887 2990
rect 17712 2933 17887 2950
rect 17712 2893 17887 2910
rect 17712 2853 17887 2870
rect 17712 2813 17887 2830
rect 17712 2773 17887 2790
rect 17712 2733 17887 2750
rect 17712 2693 17887 2710
rect 17712 2653 17887 2670
rect 17712 2613 17887 2630
rect 17712 2573 17887 2590
rect 17712 2533 17887 2550
rect 17712 2493 17887 2510
rect 17712 2453 17887 2470
rect 17712 2413 17887 2430
rect 17712 2373 17887 2390
rect 17712 2333 17887 2350
rect 17712 2293 17887 2310
rect 17712 2253 17887 2270
rect 17712 2213 17887 2230
rect 17712 2173 17887 2190
rect 17712 2133 17887 2150
rect 17712 2093 17887 2110
rect 17712 2053 17887 2070
rect 17712 2013 17887 2030
rect 17712 1973 17887 1990
rect 17712 1933 17887 1950
rect 17712 1893 17887 1910
rect 17712 1853 17887 1870
rect 17712 1813 17887 1830
rect 17712 1773 17887 1790
rect 17712 1733 17887 1750
rect 17712 1693 17887 1710
rect 17712 1653 17887 1670
rect 17712 1613 17887 1630
rect 17712 1573 17887 1590
rect 17712 1533 17887 1550
rect 17712 1493 17887 1510
rect 17712 1453 17887 1470
rect 17712 1413 17887 1430
rect 17712 1373 17887 1390
rect 17712 1333 17887 1350
rect 17712 1293 17887 1310
rect 17712 1253 17887 1270
rect 17712 1213 17887 1230
rect 17712 1173 17887 1190
rect 17712 1133 17887 1150
rect 17712 1093 17887 1110
rect 17712 1053 17887 1070
rect 17712 1013 17887 1030
rect 17712 973 17887 990
rect 17712 933 17887 950
rect 17712 893 17887 910
rect 17712 853 17887 870
rect 17712 813 17887 830
rect 17712 773 17887 790
rect 17712 733 17887 750
rect 17712 693 17887 710
rect 17712 653 17887 670
rect 17712 613 17887 630
rect 17712 573 17887 590
rect 17712 533 17887 550
rect 17712 493 17887 510
rect 17712 453 17887 470
rect 17712 413 17887 430
rect 17712 373 17887 390
rect 17712 333 17887 350
rect 17712 293 17887 310
rect 17712 253 17887 270
rect 17712 213 17887 230
rect 17712 173 17887 190
rect 17712 133 17887 150
rect 17712 93 17887 110
rect 17712 53 17887 70
rect 17712 13 17887 30
<< locali >>
rect -2452 -436 -2245 9493
rect -440 9483 -294 9514
rect -440 9455 -430 9483
rect -402 9455 -383 9483
rect -355 9455 -336 9483
rect -308 9455 -294 9483
rect -440 9436 -294 9455
rect -440 9408 -430 9436
rect -402 9408 -383 9436
rect -355 9408 -336 9436
rect -308 9408 -294 9436
rect -440 9389 -294 9408
rect -440 9361 -430 9389
rect -402 9361 -383 9389
rect -355 9361 -336 9389
rect -308 9361 -294 9389
rect -2157 9110 -1950 9274
rect -2157 9093 -2143 9110
rect -1968 9093 -1950 9110
rect -2157 9070 -1950 9093
rect -2157 9053 -2143 9070
rect -1968 9053 -1950 9070
rect -2157 9030 -1950 9053
rect -2157 9013 -2143 9030
rect -1968 9013 -1950 9030
rect -2157 8990 -1950 9013
rect -2157 8973 -2143 8990
rect -1968 8973 -1950 8990
rect -2157 8950 -1950 8973
rect -2157 8933 -2143 8950
rect -1968 8933 -1950 8950
rect -2157 8910 -1950 8933
rect -2157 8893 -2143 8910
rect -1968 8893 -1950 8910
rect -2157 8870 -1950 8893
rect -2157 8853 -2143 8870
rect -1968 8853 -1950 8870
rect -2157 8830 -1950 8853
rect -2157 8813 -2143 8830
rect -1968 8813 -1950 8830
rect -2157 8790 -1950 8813
rect -2157 8773 -2143 8790
rect -1968 8773 -1950 8790
rect -2157 8750 -1950 8773
rect -2157 8733 -2143 8750
rect -1968 8733 -1950 8750
rect -2157 8710 -1950 8733
rect -2157 8693 -2143 8710
rect -1968 8693 -1950 8710
rect -2157 8670 -1950 8693
rect -2157 8653 -2143 8670
rect -1968 8653 -1950 8670
rect -2157 8630 -1950 8653
rect -2157 8613 -2143 8630
rect -1968 8613 -1950 8630
rect -2157 8590 -1950 8613
rect -2157 8573 -2143 8590
rect -1968 8573 -1950 8590
rect -2157 8550 -1950 8573
rect -2157 8533 -2143 8550
rect -1968 8533 -1950 8550
rect -2157 8510 -1950 8533
rect -2157 8493 -2143 8510
rect -1968 8493 -1950 8510
rect -2157 8470 -1950 8493
rect -2157 8453 -2143 8470
rect -1968 8453 -1950 8470
rect -2157 8430 -1950 8453
rect -2157 8413 -2143 8430
rect -1968 8413 -1950 8430
rect -2157 8390 -1950 8413
rect -2157 8373 -2143 8390
rect -1968 8373 -1950 8390
rect -2157 8350 -1950 8373
rect -2157 8333 -2143 8350
rect -1968 8333 -1950 8350
rect -2157 8310 -1950 8333
rect -2157 8293 -2143 8310
rect -1968 8293 -1950 8310
rect -659 8424 -625 9036
rect -659 8407 -651 8424
rect -634 8407 -625 8424
rect -2157 8270 -1950 8293
rect -2157 8253 -2143 8270
rect -1968 8253 -1950 8270
rect -2157 8230 -1950 8253
rect -2157 8213 -2143 8230
rect -1968 8213 -1950 8230
rect -2157 8190 -1950 8213
rect -2157 8173 -2143 8190
rect -1968 8173 -1950 8190
rect -2157 8150 -1950 8173
rect -2157 8133 -2143 8150
rect -1968 8133 -1950 8150
rect -2157 8110 -1950 8133
rect -2157 8093 -2143 8110
rect -1968 8093 -1950 8110
rect -2157 8070 -1950 8093
rect -2157 8053 -2143 8070
rect -1968 8053 -1950 8070
rect -2157 8030 -1950 8053
rect -2157 8013 -2143 8030
rect -1968 8013 -1950 8030
rect -2157 7990 -1950 8013
rect -2157 7973 -2143 7990
rect -1968 7973 -1950 7990
rect -2157 7950 -1950 7973
rect -2157 7933 -2143 7950
rect -1968 7933 -1950 7950
rect -2157 7910 -1950 7933
rect -2157 7893 -2143 7910
rect -1968 7893 -1950 7910
rect -2157 7870 -1950 7893
rect -2157 7853 -2143 7870
rect -1968 7853 -1950 7870
rect -2157 7830 -1950 7853
rect -2157 7813 -2143 7830
rect -1968 7813 -1950 7830
rect -2157 7790 -1950 7813
rect -1374 8302 -1355 8308
rect -1374 8285 -1373 8302
rect -1356 8285 -1355 8302
rect -2157 7773 -2143 7790
rect -1968 7773 -1950 7790
rect -2157 7750 -1950 7773
rect -2157 7733 -2143 7750
rect -1968 7733 -1950 7750
rect -2157 7710 -1950 7733
rect -2157 7693 -2143 7710
rect -1968 7693 -1950 7710
rect -2157 7670 -1950 7693
rect -2157 7653 -2143 7670
rect -1968 7653 -1950 7670
rect -2157 7630 -1950 7653
rect -2157 7613 -2143 7630
rect -1968 7613 -1950 7630
rect -2157 7590 -1950 7613
rect -2157 7573 -2143 7590
rect -1968 7573 -1950 7590
rect -2157 7550 -1950 7573
rect -2157 7533 -2143 7550
rect -1968 7533 -1950 7550
rect -2157 7510 -1950 7533
rect -2157 7493 -2143 7510
rect -1968 7493 -1950 7510
rect -2157 7470 -1950 7493
rect -2157 7453 -2143 7470
rect -1968 7453 -1950 7470
rect -2157 7430 -1950 7453
rect -2157 7413 -2143 7430
rect -1968 7413 -1950 7430
rect -2157 7390 -1950 7413
rect -2157 7373 -2143 7390
rect -1968 7373 -1950 7390
rect -2157 7350 -1950 7373
rect -2157 7333 -2143 7350
rect -1968 7333 -1950 7350
rect -2157 7310 -1950 7333
rect -2157 7293 -2143 7310
rect -1968 7293 -1950 7310
rect -1410 7803 -1391 7809
rect -1410 7786 -1409 7803
rect -1392 7786 -1391 7803
rect -2157 7270 -1950 7293
rect -2157 7253 -2143 7270
rect -1968 7253 -1950 7270
rect -2157 7230 -1950 7253
rect -2157 7213 -2143 7230
rect -1968 7213 -1950 7230
rect -2157 7190 -1950 7213
rect -2157 7173 -2143 7190
rect -1968 7173 -1950 7190
rect -2157 7150 -1950 7173
rect -2157 7133 -2143 7150
rect -1968 7133 -1950 7150
rect -2157 7110 -1950 7133
rect -2157 7093 -2143 7110
rect -1968 7093 -1950 7110
rect -2157 7070 -1950 7093
rect -2157 7053 -2143 7070
rect -1968 7053 -1950 7070
rect -2157 7030 -1950 7053
rect -2157 7013 -2143 7030
rect -1968 7013 -1950 7030
rect -2157 6990 -1950 7013
rect -2157 6973 -2143 6990
rect -1968 6973 -1950 6990
rect -2157 6950 -1950 6973
rect -2157 6933 -2143 6950
rect -1968 6933 -1950 6950
rect -2157 6910 -1950 6933
rect -2157 6893 -2143 6910
rect -1968 6893 -1950 6910
rect -2157 6870 -1950 6893
rect -2157 6853 -2143 6870
rect -1968 6853 -1950 6870
rect -2157 6830 -1950 6853
rect -2157 6813 -2143 6830
rect -1968 6813 -1950 6830
rect -2157 6790 -1950 6813
rect -1446 7300 -1427 7306
rect -1446 7283 -1445 7300
rect -1428 7283 -1427 7300
rect -2157 6773 -2143 6790
rect -1968 6773 -1950 6790
rect -2157 6750 -1950 6773
rect -2157 6733 -2143 6750
rect -1968 6733 -1950 6750
rect -2157 6710 -1950 6733
rect -2157 6693 -2143 6710
rect -1968 6693 -1950 6710
rect -2157 6670 -1950 6693
rect -2157 6653 -2143 6670
rect -1968 6653 -1950 6670
rect -2157 6630 -1950 6653
rect -2157 6613 -2143 6630
rect -1968 6613 -1950 6630
rect -2157 6590 -1950 6613
rect -2157 6573 -2143 6590
rect -1968 6573 -1950 6590
rect -2157 6550 -1950 6573
rect -2157 6533 -2143 6550
rect -1968 6533 -1950 6550
rect -2157 6510 -1950 6533
rect -2157 6493 -2143 6510
rect -1968 6493 -1950 6510
rect -2157 6470 -1950 6493
rect -2157 6453 -2143 6470
rect -1968 6453 -1950 6470
rect -2157 6430 -1950 6453
rect -2157 6413 -2143 6430
rect -1968 6413 -1950 6430
rect -2157 6390 -1950 6413
rect -2157 6373 -2143 6390
rect -1968 6373 -1950 6390
rect -2157 6350 -1950 6373
rect -2157 6333 -2143 6350
rect -1968 6333 -1950 6350
rect -2157 6310 -1950 6333
rect -2157 6293 -2143 6310
rect -1968 6293 -1950 6310
rect -1482 6797 -1463 6803
rect -1482 6780 -1481 6797
rect -1464 6780 -1463 6797
rect -2157 6270 -1950 6293
rect -2157 6253 -2143 6270
rect -1968 6253 -1950 6270
rect -2157 6230 -1950 6253
rect -2157 6213 -2143 6230
rect -1968 6213 -1950 6230
rect -2157 6190 -1950 6213
rect -2157 6173 -2143 6190
rect -1968 6173 -1950 6190
rect -2157 6150 -1950 6173
rect -2157 6133 -2143 6150
rect -1968 6133 -1950 6150
rect -2157 6110 -1950 6133
rect -2157 6093 -2143 6110
rect -1968 6093 -1950 6110
rect -2157 6070 -1950 6093
rect -2157 6053 -2143 6070
rect -1968 6053 -1950 6070
rect -2157 6030 -1950 6053
rect -2157 6013 -2143 6030
rect -1968 6013 -1950 6030
rect -2157 5990 -1950 6013
rect -2157 5973 -2143 5990
rect -1968 5973 -1950 5990
rect -2157 5950 -1950 5973
rect -2157 5933 -2143 5950
rect -1968 5933 -1950 5950
rect -2157 5910 -1950 5933
rect -2157 5893 -2143 5910
rect -1968 5893 -1950 5910
rect -2157 5870 -1950 5893
rect -2157 5853 -2143 5870
rect -1968 5853 -1950 5870
rect -2157 5830 -1950 5853
rect -2157 5813 -2143 5830
rect -1968 5813 -1950 5830
rect -2157 5790 -1950 5813
rect -1518 6297 -1499 6303
rect -1518 6280 -1517 6297
rect -1500 6280 -1499 6297
rect -2157 5773 -2143 5790
rect -1968 5773 -1950 5790
rect -2157 5750 -1950 5773
rect -2157 5733 -2143 5750
rect -1968 5733 -1950 5750
rect -2157 5710 -1950 5733
rect -2157 5693 -2143 5710
rect -1968 5693 -1950 5710
rect -2157 5670 -1950 5693
rect -2157 5653 -2143 5670
rect -1968 5653 -1950 5670
rect -2157 5630 -1950 5653
rect -2157 5613 -2143 5630
rect -1968 5613 -1950 5630
rect -2157 5590 -1950 5613
rect -2157 5573 -2143 5590
rect -1968 5573 -1950 5590
rect -2157 5550 -1950 5573
rect -2157 5533 -2143 5550
rect -1968 5533 -1950 5550
rect -2157 5510 -1950 5533
rect -2157 5493 -2143 5510
rect -1968 5493 -1950 5510
rect -2157 5470 -1950 5493
rect -2157 5453 -2143 5470
rect -1968 5453 -1950 5470
rect -2157 5430 -1950 5453
rect -2157 5413 -2143 5430
rect -1968 5413 -1950 5430
rect -2157 5390 -1950 5413
rect -2157 5373 -2143 5390
rect -1968 5373 -1950 5390
rect -2157 5350 -1950 5373
rect -2157 5333 -2143 5350
rect -1968 5333 -1950 5350
rect -2157 5310 -1950 5333
rect -2157 5293 -2143 5310
rect -1968 5293 -1950 5310
rect -1554 5795 -1535 5801
rect -1554 5778 -1553 5795
rect -1536 5778 -1535 5795
rect -2157 5270 -1950 5293
rect -2157 5253 -2143 5270
rect -1968 5253 -1950 5270
rect -2157 5230 -1950 5253
rect -2157 5213 -2143 5230
rect -1968 5213 -1950 5230
rect -2157 5190 -1950 5213
rect -2157 5173 -2143 5190
rect -1968 5173 -1950 5190
rect -2157 5150 -1950 5173
rect -2157 5133 -2143 5150
rect -1968 5133 -1950 5150
rect -2157 5110 -1950 5133
rect -2157 5093 -2143 5110
rect -1968 5093 -1950 5110
rect -2157 5070 -1950 5093
rect -2157 5053 -2143 5070
rect -1968 5053 -1950 5070
rect -2157 5030 -1950 5053
rect -2157 5013 -2143 5030
rect -1968 5013 -1950 5030
rect -2157 4990 -1950 5013
rect -2157 4973 -2143 4990
rect -1968 4973 -1950 4990
rect -2157 4950 -1950 4973
rect -2157 4933 -2143 4950
rect -1968 4933 -1950 4950
rect -2157 4910 -1950 4933
rect -2157 4893 -2143 4910
rect -1968 4893 -1950 4910
rect -2157 4870 -1950 4893
rect -2157 4853 -2143 4870
rect -1968 4853 -1950 4870
rect -2157 4830 -1950 4853
rect -2157 4813 -2143 4830
rect -1968 4813 -1950 4830
rect -2157 4790 -1950 4813
rect -1590 5293 -1571 5299
rect -1590 5276 -1589 5293
rect -1572 5276 -1571 5293
rect -2157 4773 -2143 4790
rect -1968 4773 -1950 4790
rect -2157 4750 -1950 4773
rect -2157 4733 -2143 4750
rect -1968 4733 -1950 4750
rect -2157 4710 -1950 4733
rect -2157 4693 -2143 4710
rect -1968 4693 -1950 4710
rect -2157 4670 -1950 4693
rect -2157 4653 -2143 4670
rect -1968 4653 -1950 4670
rect -2157 4630 -1950 4653
rect -2157 4613 -2143 4630
rect -1968 4613 -1950 4630
rect -2157 4590 -1950 4613
rect -2157 4573 -2143 4590
rect -1968 4573 -1950 4590
rect -2157 4550 -1950 4573
rect -2157 4533 -2143 4550
rect -1968 4533 -1950 4550
rect -2157 4510 -1950 4533
rect -2157 4493 -2143 4510
rect -1968 4493 -1950 4510
rect -2157 4470 -1950 4493
rect -2157 4453 -2143 4470
rect -1968 4453 -1950 4470
rect -2157 4430 -1950 4453
rect -2157 4413 -2143 4430
rect -1968 4413 -1950 4430
rect -2157 4390 -1950 4413
rect -2157 4373 -2143 4390
rect -1968 4373 -1950 4390
rect -2157 4350 -1950 4373
rect -2157 4333 -2143 4350
rect -1968 4333 -1950 4350
rect -2157 4310 -1950 4333
rect -2157 4293 -2143 4310
rect -1968 4293 -1950 4310
rect -1626 4790 -1607 4796
rect -1626 4773 -1625 4790
rect -1608 4773 -1607 4790
rect -2157 4270 -1950 4293
rect -2157 4253 -2143 4270
rect -1968 4253 -1950 4270
rect -2157 4230 -1950 4253
rect -2157 4213 -2143 4230
rect -1968 4213 -1950 4230
rect -2157 4190 -1950 4213
rect -2157 4173 -2143 4190
rect -1968 4173 -1950 4190
rect -2157 4150 -1950 4173
rect -2157 4133 -2143 4150
rect -1968 4133 -1950 4150
rect -2157 4110 -1950 4133
rect -2157 4093 -2143 4110
rect -1968 4093 -1950 4110
rect -2157 4070 -1950 4093
rect -2157 4053 -2143 4070
rect -1968 4053 -1950 4070
rect -2157 4030 -1950 4053
rect -2157 4013 -2143 4030
rect -1968 4013 -1950 4030
rect -2157 3990 -1950 4013
rect -2157 3973 -2143 3990
rect -1968 3973 -1950 3990
rect -2157 3950 -1950 3973
rect -2157 3933 -2143 3950
rect -1968 3933 -1950 3950
rect -2157 3910 -1950 3933
rect -2157 3893 -2143 3910
rect -1968 3893 -1950 3910
rect -2157 3870 -1950 3893
rect -2157 3853 -2143 3870
rect -1968 3853 -1950 3870
rect -2157 3830 -1950 3853
rect -2157 3813 -2143 3830
rect -1968 3813 -1950 3830
rect -2157 3790 -1950 3813
rect -1662 4289 -1643 4295
rect -1662 4272 -1661 4289
rect -1644 4272 -1643 4289
rect -2157 3773 -2143 3790
rect -1968 3773 -1950 3790
rect -2157 3750 -1950 3773
rect -2157 3733 -2143 3750
rect -1968 3733 -1950 3750
rect -2157 3710 -1950 3733
rect -2157 3693 -2143 3710
rect -1968 3693 -1950 3710
rect -2157 3670 -1950 3693
rect -2157 3653 -2143 3670
rect -1968 3653 -1950 3670
rect -2157 3630 -1950 3653
rect -2157 3613 -2143 3630
rect -1968 3613 -1950 3630
rect -2157 3590 -1950 3613
rect -2157 3573 -2143 3590
rect -1968 3573 -1950 3590
rect -2157 3550 -1950 3573
rect -2157 3533 -2143 3550
rect -1968 3533 -1950 3550
rect -2157 3510 -1950 3533
rect -2157 3493 -2143 3510
rect -1968 3493 -1950 3510
rect -2157 3470 -1950 3493
rect -2157 3453 -2143 3470
rect -1968 3453 -1950 3470
rect -2157 3430 -1950 3453
rect -2157 3413 -2143 3430
rect -1968 3413 -1950 3430
rect -2157 3390 -1950 3413
rect -2157 3373 -2143 3390
rect -1968 3373 -1950 3390
rect -2157 3350 -1950 3373
rect -2157 3333 -2143 3350
rect -1968 3333 -1950 3350
rect -2157 3310 -1950 3333
rect -2157 3293 -2143 3310
rect -1968 3293 -1950 3310
rect -2157 3270 -1950 3293
rect -1698 3787 -1679 3793
rect -1698 3770 -1697 3787
rect -1680 3770 -1679 3787
rect -2157 3253 -2143 3270
rect -1968 3253 -1950 3270
rect -2157 3230 -1950 3253
rect -2157 3213 -2143 3230
rect -1968 3213 -1950 3230
rect -2157 3190 -1950 3213
rect -2157 3173 -2143 3190
rect -1968 3173 -1950 3190
rect -2157 3150 -1950 3173
rect -2157 3133 -2143 3150
rect -1968 3133 -1950 3150
rect -2157 3110 -1950 3133
rect -2157 3093 -2143 3110
rect -1968 3093 -1950 3110
rect -2157 3070 -1950 3093
rect -2157 3053 -2143 3070
rect -1968 3053 -1950 3070
rect -2157 3030 -1950 3053
rect -2157 3013 -2143 3030
rect -1968 3013 -1950 3030
rect -2157 2990 -1950 3013
rect -2157 2973 -2143 2990
rect -1968 2973 -1950 2990
rect -2157 2950 -1950 2973
rect -2157 2933 -2143 2950
rect -1968 2933 -1950 2950
rect -2157 2910 -1950 2933
rect -2157 2893 -2143 2910
rect -1968 2893 -1950 2910
rect -2157 2870 -1950 2893
rect -2157 2853 -2143 2870
rect -1968 2853 -1950 2870
rect -2157 2830 -1950 2853
rect -2157 2813 -2143 2830
rect -1968 2813 -1950 2830
rect -2157 2790 -1950 2813
rect -2157 2773 -2143 2790
rect -1968 2773 -1950 2790
rect -1734 3285 -1715 3291
rect -1734 3268 -1733 3285
rect -1716 3268 -1715 3285
rect -2157 2750 -1950 2773
rect -2157 2733 -2143 2750
rect -1968 2733 -1950 2750
rect -2157 2710 -1950 2733
rect -2157 2693 -2143 2710
rect -1968 2693 -1950 2710
rect -2157 2670 -1950 2693
rect -2157 2653 -2143 2670
rect -1968 2653 -1950 2670
rect -2157 2630 -1950 2653
rect -2157 2613 -2143 2630
rect -1968 2613 -1950 2630
rect -2157 2590 -1950 2613
rect -2157 2573 -2143 2590
rect -1968 2573 -1950 2590
rect -2157 2550 -1950 2573
rect -2157 2533 -2143 2550
rect -1968 2533 -1950 2550
rect -2157 2510 -1950 2533
rect -2157 2493 -2143 2510
rect -1968 2493 -1950 2510
rect -2157 2470 -1950 2493
rect -2157 2453 -2143 2470
rect -1968 2453 -1950 2470
rect -2157 2430 -1950 2453
rect -2157 2413 -2143 2430
rect -1968 2413 -1950 2430
rect -2157 2390 -1950 2413
rect -2157 2373 -2143 2390
rect -1968 2373 -1950 2390
rect -2157 2350 -1950 2373
rect -2157 2333 -2143 2350
rect -1968 2333 -1950 2350
rect -2157 2310 -1950 2333
rect -2157 2293 -2143 2310
rect -1968 2293 -1950 2310
rect -2157 2270 -1950 2293
rect -1770 2783 -1751 2789
rect -1770 2766 -1769 2783
rect -1752 2766 -1751 2783
rect -2157 2253 -2143 2270
rect -1968 2253 -1950 2270
rect -2157 2230 -1950 2253
rect -2157 2213 -2143 2230
rect -1968 2213 -1950 2230
rect -2157 2190 -1950 2213
rect -2157 2173 -2143 2190
rect -1968 2173 -1950 2190
rect -2157 2150 -1950 2173
rect -2157 2133 -2143 2150
rect -1968 2133 -1950 2150
rect -2157 2110 -1950 2133
rect -2157 2093 -2143 2110
rect -1968 2093 -1950 2110
rect -2157 2070 -1950 2093
rect -2157 2053 -2143 2070
rect -1968 2053 -1950 2070
rect -2157 2030 -1950 2053
rect -2157 2013 -2143 2030
rect -1968 2013 -1950 2030
rect -2157 1990 -1950 2013
rect -2157 1973 -2143 1990
rect -1968 1973 -1950 1990
rect -2157 1950 -1950 1973
rect -2157 1933 -2143 1950
rect -1968 1933 -1950 1950
rect -2157 1910 -1950 1933
rect -2157 1893 -2143 1910
rect -1968 1893 -1950 1910
rect -2157 1870 -1950 1893
rect -2157 1853 -2143 1870
rect -1968 1853 -1950 1870
rect -2157 1830 -1950 1853
rect -2157 1813 -2143 1830
rect -1968 1813 -1950 1830
rect -2157 1790 -1950 1813
rect -2157 1773 -2143 1790
rect -1968 1773 -1950 1790
rect -1806 2282 -1787 2288
rect -1806 2265 -1805 2282
rect -1788 2265 -1787 2282
rect -2157 1750 -1950 1773
rect -2157 1733 -2143 1750
rect -1968 1733 -1950 1750
rect -2157 1710 -1950 1733
rect -2157 1693 -2143 1710
rect -1968 1693 -1950 1710
rect -2157 1670 -1950 1693
rect -2157 1653 -2143 1670
rect -1968 1653 -1950 1670
rect -2157 1630 -1950 1653
rect -2157 1613 -2143 1630
rect -1968 1613 -1950 1630
rect -2157 1590 -1950 1613
rect -2157 1573 -2143 1590
rect -1968 1573 -1950 1590
rect -2157 1550 -1950 1573
rect -2157 1533 -2143 1550
rect -1968 1533 -1950 1550
rect -2157 1510 -1950 1533
rect -2157 1493 -2143 1510
rect -1968 1493 -1950 1510
rect -2157 1470 -1950 1493
rect -2157 1453 -2143 1470
rect -1968 1453 -1950 1470
rect -2157 1430 -1950 1453
rect -2157 1413 -2143 1430
rect -1968 1413 -1950 1430
rect -2157 1390 -1950 1413
rect -2157 1373 -2143 1390
rect -1968 1373 -1950 1390
rect -2157 1350 -1950 1373
rect -2157 1333 -2143 1350
rect -1968 1333 -1950 1350
rect -2157 1310 -1950 1333
rect -2157 1293 -2143 1310
rect -1968 1293 -1950 1310
rect -2157 1270 -1950 1293
rect -1842 1779 -1823 1785
rect -1842 1762 -1841 1779
rect -1824 1762 -1823 1779
rect -2157 1253 -2143 1270
rect -1968 1253 -1950 1270
rect -2157 1230 -1950 1253
rect -2157 1213 -2143 1230
rect -1968 1213 -1950 1230
rect -2157 1190 -1950 1213
rect -2157 1173 -2143 1190
rect -1968 1173 -1950 1190
rect -2157 1150 -1950 1173
rect -2157 1133 -2143 1150
rect -1968 1133 -1950 1150
rect -2157 1110 -1950 1133
rect -2157 1093 -2143 1110
rect -1968 1093 -1950 1110
rect -2157 1070 -1950 1093
rect -2157 1053 -2143 1070
rect -1968 1053 -1950 1070
rect -2157 1030 -1950 1053
rect -2157 1013 -2143 1030
rect -1968 1013 -1950 1030
rect -2157 990 -1950 1013
rect -2157 973 -2143 990
rect -1968 973 -1950 990
rect -2157 950 -1950 973
rect -2157 933 -2143 950
rect -1968 933 -1950 950
rect -2157 910 -1950 933
rect -2157 893 -2143 910
rect -1968 893 -1950 910
rect -2157 870 -1950 893
rect -2157 853 -2143 870
rect -1968 853 -1950 870
rect -2157 830 -1950 853
rect -2157 813 -2143 830
rect -1968 813 -1950 830
rect -2157 790 -1950 813
rect -2157 773 -2143 790
rect -1968 773 -1950 790
rect -1878 1276 -1859 1282
rect -1878 1259 -1877 1276
rect -1860 1259 -1859 1276
rect -2157 750 -1950 773
rect -2157 733 -2143 750
rect -1968 733 -1950 750
rect -2157 710 -1950 733
rect -2157 693 -2143 710
rect -1968 693 -1950 710
rect -2157 670 -1950 693
rect -2157 653 -2143 670
rect -1968 653 -1950 670
rect -2157 630 -1950 653
rect -2157 613 -2143 630
rect -1968 613 -1950 630
rect -2157 590 -1950 613
rect -2157 573 -2143 590
rect -1968 573 -1950 590
rect -2157 550 -1950 573
rect -2157 533 -2143 550
rect -1968 533 -1950 550
rect -2157 510 -1950 533
rect -2157 493 -2143 510
rect -1968 493 -1950 510
rect -2157 470 -1950 493
rect -2157 453 -2143 470
rect -1968 453 -1950 470
rect -2157 430 -1950 453
rect -2157 413 -2143 430
rect -1968 413 -1950 430
rect -2157 390 -1950 413
rect -2157 373 -2143 390
rect -1968 373 -1950 390
rect -2157 350 -1950 373
rect -2157 333 -2143 350
rect -1968 333 -1950 350
rect -2157 310 -1950 333
rect -2157 293 -2143 310
rect -1968 293 -1950 310
rect -2157 270 -1950 293
rect -2157 253 -2143 270
rect -1968 253 -1950 270
rect -2157 230 -1950 253
rect -2157 213 -2143 230
rect -1968 213 -1950 230
rect -2157 190 -1950 213
rect -2157 173 -2143 190
rect -1968 173 -1950 190
rect -2157 150 -1950 173
rect -2157 133 -2143 150
rect -1968 133 -1950 150
rect -2157 110 -1950 133
rect -2157 93 -2143 110
rect -1968 93 -1950 110
rect -2157 70 -1950 93
rect -2157 53 -2143 70
rect -1968 53 -1950 70
rect -2157 30 -1950 53
rect -2157 13 -2143 30
rect -1968 13 -1950 30
rect -2157 -217 -1950 13
rect -1914 775 -1895 781
rect -1914 758 -1913 775
rect -1896 758 -1895 775
rect -1914 -457 -1895 758
rect -1878 -457 -1859 1259
rect -1842 -457 -1823 1762
rect -1806 -457 -1787 2265
rect -1770 -457 -1751 2766
rect -1734 -457 -1715 3268
rect -1698 -457 -1679 3770
rect -1662 -457 -1643 4272
rect -1626 -457 -1607 4773
rect -1590 -457 -1571 5276
rect -1554 -457 -1535 5778
rect -1518 -457 -1499 6280
rect -1482 -457 -1463 6780
rect -1446 -457 -1427 7283
rect -1410 -457 -1391 7786
rect -1374 -457 -1355 8285
rect -762 8261 -743 8267
rect -762 8244 -761 8261
rect -744 8244 -743 8261
rect -798 7759 -779 7765
rect -798 7742 -797 7759
rect -780 7742 -779 7759
rect -834 7259 -815 7265
rect -834 7242 -833 7259
rect -816 7242 -815 7259
rect -870 6757 -851 6763
rect -870 6740 -869 6757
rect -852 6740 -851 6757
rect -906 6256 -887 6262
rect -906 6239 -905 6256
rect -888 6239 -887 6256
rect -942 5752 -923 5758
rect -942 5735 -941 5752
rect -924 5735 -923 5752
rect -978 5252 -959 5258
rect -978 5235 -977 5252
rect -960 5235 -959 5252
rect -1014 4749 -995 4755
rect -1014 4732 -1013 4749
rect -996 4732 -995 4749
rect -1050 4250 -1031 4256
rect -1050 4233 -1049 4250
rect -1032 4233 -1031 4250
rect -1086 3747 -1067 3753
rect -1086 3730 -1085 3747
rect -1068 3730 -1067 3747
rect -1122 3245 -1103 3251
rect -1122 3228 -1121 3245
rect -1104 3228 -1103 3245
rect -1158 2744 -1139 2750
rect -1158 2727 -1157 2744
rect -1140 2727 -1139 2744
rect -1194 2239 -1175 2245
rect -1194 2222 -1193 2239
rect -1176 2222 -1175 2239
rect -1230 1736 -1211 1742
rect -1230 1719 -1229 1736
rect -1212 1719 -1211 1736
rect -1266 1233 -1247 1239
rect -1266 1216 -1265 1233
rect -1248 1216 -1247 1233
rect -1302 735 -1283 741
rect -1302 718 -1301 735
rect -1284 718 -1283 735
rect -1302 -457 -1283 718
rect -1266 -457 -1247 1216
rect -1230 -457 -1211 1719
rect -1194 -457 -1175 2222
rect -1158 -457 -1139 2727
rect -1122 -457 -1103 3228
rect -1086 -457 -1067 3730
rect -1050 -457 -1031 4233
rect -1014 -457 -995 4732
rect -978 -457 -959 5235
rect -942 -457 -923 5735
rect -906 -457 -887 6239
rect -870 -457 -851 6740
rect -834 -457 -815 7242
rect -798 -457 -779 7742
rect -762 -457 -743 8244
rect -659 7922 -625 8407
rect -659 7905 -651 7922
rect -634 7905 -625 7922
rect -659 7420 -625 7905
rect -659 7403 -651 7420
rect -634 7403 -625 7420
rect -659 6918 -625 7403
rect -659 6901 -651 6918
rect -634 6901 -625 6918
rect -659 6416 -625 6901
rect -659 6399 -651 6416
rect -634 6399 -625 6416
rect -659 5914 -625 6399
rect -659 5897 -651 5914
rect -634 5897 -625 5914
rect -659 5412 -625 5897
rect -659 5395 -651 5412
rect -634 5395 -625 5412
rect -659 4910 -625 5395
rect -659 4893 -651 4910
rect -634 4893 -625 4910
rect -659 4408 -625 4893
rect -659 4391 -651 4408
rect -634 4391 -625 4408
rect -659 3906 -625 4391
rect -659 3889 -651 3906
rect -634 3889 -625 3906
rect -659 3404 -625 3889
rect -659 3387 -651 3404
rect -634 3387 -625 3404
rect -659 2902 -625 3387
rect -659 2885 -651 2902
rect -634 2885 -625 2902
rect -659 2400 -625 2885
rect -659 2383 -651 2400
rect -634 2383 -625 2400
rect -659 1898 -625 2383
rect -659 1881 -651 1898
rect -634 1881 -625 1898
rect -659 1396 -625 1881
rect -659 1379 -651 1396
rect -634 1379 -625 1396
rect -659 894 -625 1379
rect -659 877 -651 894
rect -634 877 -625 894
rect -659 -457 -625 877
rect -605 8230 -571 9036
rect -605 8213 -597 8230
rect -580 8213 -571 8230
rect -605 7728 -571 8213
rect -605 7711 -597 7728
rect -580 7711 -571 7728
rect -605 7226 -571 7711
rect -605 7209 -597 7226
rect -580 7209 -571 7226
rect -605 6724 -571 7209
rect -605 6707 -597 6724
rect -580 6707 -571 6724
rect -605 6222 -571 6707
rect -605 6205 -597 6222
rect -580 6205 -571 6222
rect -605 5720 -571 6205
rect -605 5703 -597 5720
rect -580 5703 -571 5720
rect -605 5218 -571 5703
rect -605 5201 -597 5218
rect -580 5201 -571 5218
rect -605 4716 -571 5201
rect -605 4699 -597 4716
rect -580 4699 -571 4716
rect -605 4214 -571 4699
rect -605 4197 -597 4214
rect -580 4197 -571 4214
rect -605 3712 -571 4197
rect -605 3695 -597 3712
rect -580 3695 -571 3712
rect -605 3210 -571 3695
rect -605 3193 -597 3210
rect -580 3193 -571 3210
rect -605 2708 -571 3193
rect -605 2691 -597 2708
rect -580 2691 -571 2708
rect -605 2206 -571 2691
rect -605 2189 -597 2206
rect -580 2189 -571 2206
rect -605 1704 -571 2189
rect -605 1687 -597 1704
rect -580 1687 -571 1704
rect -605 1202 -571 1687
rect -605 1185 -597 1202
rect -580 1185 -571 1202
rect -605 700 -571 1185
rect -605 683 -597 700
rect -580 683 -571 700
rect -605 -457 -571 683
rect -551 8661 -483 9036
rect -551 8641 -545 8661
rect -525 8641 -506 8661
rect -486 8641 -483 8661
rect -551 8159 -483 8641
rect -551 8139 -545 8159
rect -525 8139 -506 8159
rect -486 8139 -483 8159
rect -551 7657 -483 8139
rect -551 7637 -545 7657
rect -525 7637 -506 7657
rect -486 7637 -483 7657
rect -551 7155 -483 7637
rect -551 7135 -545 7155
rect -525 7135 -506 7155
rect -486 7135 -483 7155
rect -551 6653 -483 7135
rect -551 6633 -545 6653
rect -525 6633 -506 6653
rect -486 6633 -483 6653
rect -551 6151 -483 6633
rect -551 6131 -545 6151
rect -525 6131 -506 6151
rect -486 6131 -483 6151
rect -551 5649 -483 6131
rect -551 5629 -545 5649
rect -525 5629 -506 5649
rect -486 5629 -483 5649
rect -551 5147 -483 5629
rect -551 5127 -545 5147
rect -525 5127 -506 5147
rect -486 5127 -483 5147
rect -551 4645 -483 5127
rect -551 4625 -545 4645
rect -525 4625 -506 4645
rect -486 4625 -483 4645
rect -551 4143 -483 4625
rect -551 4123 -545 4143
rect -525 4123 -506 4143
rect -486 4123 -483 4143
rect -551 3641 -483 4123
rect -551 3621 -545 3641
rect -525 3621 -506 3641
rect -486 3621 -483 3641
rect -551 3139 -483 3621
rect -551 3119 -545 3139
rect -525 3119 -506 3139
rect -486 3119 -483 3139
rect -551 2637 -483 3119
rect -551 2617 -545 2637
rect -525 2617 -506 2637
rect -486 2617 -483 2637
rect -551 2135 -483 2617
rect -551 2115 -545 2135
rect -525 2115 -506 2135
rect -486 2115 -483 2135
rect -551 1633 -483 2115
rect -551 1613 -545 1633
rect -525 1613 -506 1633
rect -486 1613 -483 1633
rect -551 1131 -483 1613
rect -551 1111 -545 1131
rect -525 1111 -506 1131
rect -486 1111 -483 1131
rect -551 629 -483 1111
rect -551 609 -545 629
rect -525 609 -506 629
rect -486 609 -483 629
rect -551 127 -483 609
rect -551 107 -545 127
rect -525 107 -506 127
rect -486 107 -483 127
rect -551 -457 -483 107
rect -440 8957 -294 9361
rect -440 8937 -434 8957
rect -414 8937 -395 8957
rect -375 8937 -356 8957
rect -336 8937 -317 8957
rect -297 8937 -294 8957
rect -440 8915 -294 8937
rect -440 8895 -434 8915
rect -414 8895 -395 8915
rect -375 8895 -356 8915
rect -336 8895 -317 8915
rect -297 8895 -294 8915
rect -440 8787 -294 8895
rect -440 8767 -434 8787
rect -414 8767 -395 8787
rect -375 8767 -356 8787
rect -336 8767 -317 8787
rect -297 8767 -294 8787
rect -440 8455 -294 8767
rect -440 8435 -434 8455
rect -414 8435 -395 8455
rect -375 8435 -356 8455
rect -336 8435 -317 8455
rect -297 8435 -294 8455
rect -440 7953 -294 8435
rect -440 7933 -434 7953
rect -414 7933 -395 7953
rect -375 7933 -356 7953
rect -336 7933 -317 7953
rect -297 7933 -294 7953
rect -440 7451 -294 7933
rect -440 7431 -434 7451
rect -414 7431 -395 7451
rect -375 7431 -356 7451
rect -336 7431 -317 7451
rect -297 7431 -294 7451
rect -440 6949 -294 7431
rect -440 6929 -434 6949
rect -414 6929 -395 6949
rect -375 6929 -356 6949
rect -336 6929 -317 6949
rect -297 6929 -294 6949
rect -440 6447 -294 6929
rect -440 6427 -434 6447
rect -414 6427 -395 6447
rect -375 6427 -356 6447
rect -336 6427 -317 6447
rect -297 6427 -294 6447
rect -440 5945 -294 6427
rect -440 5925 -434 5945
rect -414 5925 -395 5945
rect -375 5925 -356 5945
rect -336 5925 -317 5945
rect -297 5925 -294 5945
rect -440 5443 -294 5925
rect -440 5423 -434 5443
rect -414 5423 -395 5443
rect -375 5423 -356 5443
rect -336 5423 -317 5443
rect -297 5423 -294 5443
rect -440 4941 -294 5423
rect -440 4921 -434 4941
rect -414 4921 -395 4941
rect -375 4921 -356 4941
rect -336 4921 -317 4941
rect -297 4921 -294 4941
rect -440 4439 -294 4921
rect -440 4419 -434 4439
rect -414 4419 -395 4439
rect -375 4419 -356 4439
rect -336 4419 -317 4439
rect -297 4419 -294 4439
rect -440 3937 -294 4419
rect -440 3917 -434 3937
rect -414 3917 -395 3937
rect -375 3917 -356 3937
rect -336 3917 -317 3937
rect -297 3917 -294 3937
rect -440 3435 -294 3917
rect -440 3415 -434 3435
rect -414 3415 -395 3435
rect -375 3415 -356 3435
rect -336 3415 -317 3435
rect -297 3415 -294 3435
rect -440 2933 -294 3415
rect -440 2913 -434 2933
rect -414 2913 -395 2933
rect -375 2913 -356 2933
rect -336 2913 -317 2933
rect -297 2913 -294 2933
rect -440 2431 -294 2913
rect -440 2411 -434 2431
rect -414 2411 -395 2431
rect -375 2411 -356 2431
rect -336 2411 -317 2431
rect -297 2411 -294 2431
rect -440 1929 -294 2411
rect -440 1909 -434 1929
rect -414 1909 -395 1929
rect -375 1909 -356 1929
rect -336 1909 -317 1929
rect -297 1909 -294 1929
rect -440 1427 -294 1909
rect -440 1407 -434 1427
rect -414 1407 -395 1427
rect -375 1407 -356 1427
rect -336 1407 -317 1427
rect -297 1407 -294 1427
rect -440 925 -294 1407
rect -440 905 -434 925
rect -414 905 -395 925
rect -375 905 -356 925
rect -336 905 -317 925
rect -297 905 -294 925
rect -440 423 -294 905
rect -440 403 -434 423
rect -414 403 -395 423
rect -375 403 -356 423
rect -336 403 -317 423
rect -297 403 -294 423
rect -440 381 -294 403
rect -440 361 -434 381
rect -414 361 -395 381
rect -375 361 -356 381
rect -336 361 -317 381
rect -297 361 -294 381
rect -440 -304 -294 361
rect -440 -332 -430 -304
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -332 -294 -304
rect -440 -351 -294 -332
rect -440 -379 -430 -351
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -294 -351
rect -440 -398 -294 -379
rect -440 -426 -430 -398
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -294 -398
rect -440 -457 -294 -426
rect -251 9264 -105 9514
rect -251 9236 -241 9264
rect -213 9236 -194 9264
rect -166 9236 -147 9264
rect -119 9236 -105 9264
rect -251 9217 -105 9236
rect -251 9189 -241 9217
rect -213 9189 -194 9217
rect -166 9189 -147 9217
rect -119 9189 -105 9217
rect -251 9170 -105 9189
rect -251 9142 -241 9170
rect -213 9142 -194 9170
rect -166 9142 -147 9170
rect -119 9142 -105 9170
rect -251 8731 -105 9142
rect -251 8711 -245 8731
rect -225 8711 -206 8731
rect -186 8711 -167 8731
rect -147 8711 -128 8731
rect -108 8711 -105 8731
rect -251 8626 -105 8711
rect -251 8606 -245 8626
rect -225 8606 -206 8626
rect -186 8606 -167 8626
rect -147 8606 -128 8626
rect -108 8606 -105 8626
rect -251 8124 -105 8606
rect -251 8104 -245 8124
rect -225 8104 -206 8124
rect -186 8104 -167 8124
rect -147 8104 -128 8124
rect -108 8104 -105 8124
rect -251 7622 -105 8104
rect -251 7602 -245 7622
rect -225 7602 -206 7622
rect -186 7602 -167 7622
rect -147 7602 -128 7622
rect -108 7602 -105 7622
rect -251 7120 -105 7602
rect -251 7100 -245 7120
rect -225 7100 -206 7120
rect -186 7100 -167 7120
rect -147 7100 -128 7120
rect -108 7100 -105 7120
rect -251 6618 -105 7100
rect -251 6598 -245 6618
rect -225 6598 -206 6618
rect -186 6598 -167 6618
rect -147 6598 -128 6618
rect -108 6598 -105 6618
rect -251 6116 -105 6598
rect -251 6096 -245 6116
rect -225 6096 -206 6116
rect -186 6096 -167 6116
rect -147 6096 -128 6116
rect -108 6096 -105 6116
rect -251 5614 -105 6096
rect -251 5594 -245 5614
rect -225 5594 -206 5614
rect -186 5594 -167 5614
rect -147 5594 -128 5614
rect -108 5594 -105 5614
rect -251 5112 -105 5594
rect -251 5092 -245 5112
rect -225 5092 -206 5112
rect -186 5092 -167 5112
rect -147 5092 -128 5112
rect -108 5092 -105 5112
rect -251 4610 -105 5092
rect -251 4590 -245 4610
rect -225 4590 -206 4610
rect -186 4590 -167 4610
rect -147 4590 -128 4610
rect -108 4590 -105 4610
rect -251 4108 -105 4590
rect -251 4088 -245 4108
rect -225 4088 -206 4108
rect -186 4088 -167 4108
rect -147 4088 -128 4108
rect -108 4088 -105 4108
rect -251 3606 -105 4088
rect -251 3586 -245 3606
rect -225 3586 -206 3606
rect -186 3586 -167 3606
rect -147 3586 -128 3606
rect -108 3586 -105 3606
rect -251 3104 -105 3586
rect -251 3084 -245 3104
rect -225 3084 -206 3104
rect -186 3084 -167 3104
rect -147 3084 -128 3104
rect -108 3084 -105 3104
rect -251 2602 -105 3084
rect -251 2582 -245 2602
rect -225 2582 -206 2602
rect -186 2582 -167 2602
rect -147 2582 -128 2602
rect -108 2582 -105 2602
rect -251 2100 -105 2582
rect -251 2080 -245 2100
rect -225 2080 -206 2100
rect -186 2080 -167 2100
rect -147 2080 -128 2100
rect -108 2080 -105 2100
rect -251 1598 -105 2080
rect -251 1578 -245 1598
rect -225 1578 -206 1598
rect -186 1578 -167 1598
rect -147 1578 -128 1598
rect -108 1578 -105 1598
rect -251 1096 -105 1578
rect -251 1076 -245 1096
rect -225 1076 -206 1096
rect -186 1076 -167 1096
rect -147 1076 -128 1096
rect -108 1076 -105 1096
rect -251 594 -105 1076
rect -251 574 -245 594
rect -225 574 -206 594
rect -186 574 -167 594
rect -147 574 -128 594
rect -108 574 -105 594
rect -251 253 -105 574
rect -251 233 -245 253
rect -225 233 -206 253
rect -186 233 -167 253
rect -147 233 -128 253
rect -108 233 -105 253
rect -251 197 -105 233
rect -251 177 -245 197
rect -225 177 -206 197
rect -186 177 -167 197
rect -147 177 -128 197
rect -108 177 -105 197
rect -251 92 -105 177
rect -251 72 -245 92
rect -225 72 -206 92
rect -186 72 -167 92
rect -147 72 -128 92
rect -108 72 -105 92
rect -251 -85 -105 72
rect 17167 9259 17313 9509
rect 17167 9231 17181 9259
rect 17209 9231 17228 9259
rect 17256 9231 17275 9259
rect 17303 9231 17313 9259
rect 17167 9212 17313 9231
rect 17167 9184 17181 9212
rect 17209 9184 17228 9212
rect 17256 9184 17275 9212
rect 17303 9184 17313 9212
rect 17167 9165 17313 9184
rect 17167 9137 17181 9165
rect 17209 9137 17228 9165
rect 17256 9137 17275 9165
rect 17303 9137 17313 9165
rect 17167 8626 17313 9137
rect 17167 8606 17170 8626
rect 17190 8606 17209 8626
rect 17229 8606 17248 8626
rect 17268 8606 17287 8626
rect 17307 8606 17313 8626
rect 17167 8124 17313 8606
rect 17167 8104 17170 8124
rect 17190 8104 17209 8124
rect 17229 8104 17248 8124
rect 17268 8104 17287 8124
rect 17307 8104 17313 8124
rect 17167 7622 17313 8104
rect 17167 7602 17170 7622
rect 17190 7602 17209 7622
rect 17229 7602 17248 7622
rect 17268 7602 17287 7622
rect 17307 7602 17313 7622
rect 17167 7120 17313 7602
rect 17167 7100 17170 7120
rect 17190 7100 17209 7120
rect 17229 7100 17248 7120
rect 17268 7100 17287 7120
rect 17307 7100 17313 7120
rect 17167 6618 17313 7100
rect 17167 6598 17170 6618
rect 17190 6598 17209 6618
rect 17229 6598 17248 6618
rect 17268 6598 17287 6618
rect 17307 6598 17313 6618
rect 17167 6116 17313 6598
rect 17167 6096 17170 6116
rect 17190 6096 17209 6116
rect 17229 6096 17248 6116
rect 17268 6096 17287 6116
rect 17307 6096 17313 6116
rect 17167 5614 17313 6096
rect 17167 5594 17170 5614
rect 17190 5594 17209 5614
rect 17229 5594 17248 5614
rect 17268 5594 17287 5614
rect 17307 5594 17313 5614
rect 17167 5112 17313 5594
rect 17167 5092 17170 5112
rect 17190 5092 17209 5112
rect 17229 5092 17248 5112
rect 17268 5092 17287 5112
rect 17307 5092 17313 5112
rect 17167 4610 17313 5092
rect 17167 4590 17170 4610
rect 17190 4590 17209 4610
rect 17229 4590 17248 4610
rect 17268 4590 17287 4610
rect 17307 4590 17313 4610
rect 17167 4108 17313 4590
rect 17167 4088 17170 4108
rect 17190 4088 17209 4108
rect 17229 4088 17248 4108
rect 17268 4088 17287 4108
rect 17307 4088 17313 4108
rect 17167 3606 17313 4088
rect 17167 3586 17170 3606
rect 17190 3586 17209 3606
rect 17229 3586 17248 3606
rect 17268 3586 17287 3606
rect 17307 3586 17313 3606
rect 17167 3104 17313 3586
rect 17167 3084 17170 3104
rect 17190 3084 17209 3104
rect 17229 3084 17248 3104
rect 17268 3084 17287 3104
rect 17307 3084 17313 3104
rect 17167 2602 17313 3084
rect 17167 2582 17170 2602
rect 17190 2582 17209 2602
rect 17229 2582 17248 2602
rect 17268 2582 17287 2602
rect 17307 2582 17313 2602
rect 17167 2100 17313 2582
rect 17167 2080 17170 2100
rect 17190 2080 17209 2100
rect 17229 2080 17248 2100
rect 17268 2080 17287 2100
rect 17307 2080 17313 2100
rect 17167 1598 17313 2080
rect 17167 1578 17170 1598
rect 17190 1578 17209 1598
rect 17229 1578 17248 1598
rect 17268 1578 17287 1598
rect 17307 1578 17313 1598
rect 17167 1096 17313 1578
rect 17167 1076 17170 1096
rect 17190 1076 17209 1096
rect 17229 1076 17248 1096
rect 17268 1076 17287 1096
rect 17307 1076 17313 1096
rect 17167 594 17313 1076
rect 17167 574 17170 594
rect 17190 574 17209 594
rect 17229 574 17248 594
rect 17268 574 17287 594
rect 17307 574 17313 594
rect 17167 92 17313 574
rect 17167 72 17170 92
rect 17190 72 17209 92
rect 17229 72 17248 92
rect 17268 72 17287 92
rect 17307 72 17313 92
rect -251 -113 -241 -85
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -105 -85
rect -251 -132 -105 -113
rect -251 -160 -241 -132
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -105 -132
rect -251 -179 -105 -160
rect -251 -207 -241 -179
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -105 -179
rect -251 -457 -105 -207
rect 427 -292 444 0
rect 422 -295 444 -292
rect 422 -312 425 -295
rect 442 -312 444 -295
rect 422 -316 444 -312
rect 929 -457 946 0
rect 1431 -457 1448 0
rect 1933 -457 1950 0
rect 2435 -457 2452 0
rect 2937 -457 2954 0
rect 3439 -457 3456 0
rect 3941 -457 3958 0
rect 4443 -457 4460 0
rect 4779 -457 4796 0
rect 4945 -457 4962 0
rect 5447 -457 5464 0
rect 5949 -457 5966 0
rect 6451 -457 6468 0
rect 6953 -457 6970 0
rect 7455 -457 7472 0
rect 7957 -457 7974 0
rect 8459 -457 8476 0
rect 8795 -457 8812 0
rect 8961 -457 8978 0
rect 9463 -457 9480 0
rect 9965 -457 9982 0
rect 10467 -457 10484 0
rect 10969 -457 10986 0
rect 11471 -457 11488 0
rect 11973 -457 11990 0
rect 12475 -457 12492 0
rect 12811 -457 12828 0
rect 12977 -457 12994 0
rect 13479 -60 13496 0
rect 13079 -77 13496 -60
rect 13079 -457 13096 -77
rect 13981 -95 13998 0
rect 13181 -112 13998 -95
rect 13181 -457 13198 -112
rect 13283 -136 13300 -135
rect 13283 -457 13300 -153
rect 14483 -136 14500 0
rect 14483 -157 14500 -153
rect 13385 -175 13402 -174
rect 13385 -457 13402 -192
rect 14985 -175 15002 0
rect 14985 -196 15002 -192
rect 13487 -213 13504 -212
rect 13487 -457 13504 -230
rect 15487 -213 15504 0
rect 15487 -234 15504 -230
rect 13589 -251 13606 -250
rect 13589 -457 13606 -268
rect 15989 -251 16006 0
rect 16238 -26 16255 0
rect 15989 -272 16006 -268
rect 16043 -43 16255 -26
rect 13691 -289 13708 -288
rect 13691 -457 13708 -306
rect 16043 -456 16060 -43
rect 16104 -64 16121 -61
rect 16104 -456 16121 -81
rect 16274 -113 16291 0
rect 16348 -64 16365 0
rect 16348 -85 16365 -81
rect 16274 -135 16418 -113
rect 16401 -432 16418 -135
rect 16491 -289 16508 0
rect 16491 -310 16508 -306
rect 16993 -295 17010 0
rect 17167 -20 17313 72
rect 17167 -48 17181 -20
rect 17209 -48 17228 -20
rect 17256 -48 17275 -20
rect 17303 -48 17313 -20
rect 17167 -67 17313 -48
rect 17167 -95 17181 -67
rect 17209 -95 17228 -67
rect 17256 -95 17275 -67
rect 17303 -95 17313 -67
rect 17167 -114 17313 -95
rect 17167 -142 17181 -114
rect 17209 -142 17228 -114
rect 17256 -142 17275 -114
rect 17303 -142 17313 -114
rect 16993 -298 17014 -295
rect 16993 -315 16995 -298
rect 17012 -315 17014 -298
rect 16993 -318 17014 -315
rect 17167 -392 17313 -142
rect 17355 9478 17502 9509
rect 17355 9450 17370 9478
rect 17398 9450 17417 9478
rect 17445 9450 17464 9478
rect 17492 9450 17502 9478
rect 17355 9431 17502 9450
rect 17355 9403 17370 9431
rect 17398 9403 17417 9431
rect 17445 9403 17464 9431
rect 17492 9403 17502 9431
rect 17355 9384 17502 9403
rect 17355 9356 17370 9384
rect 17398 9356 17417 9384
rect 17445 9356 17464 9384
rect 17492 9356 17502 9384
rect 17355 9036 17502 9356
rect 17694 9110 17901 9274
rect 17694 9093 17712 9110
rect 17887 9093 17901 9110
rect 17694 9070 17901 9093
rect 17694 9053 17712 9070
rect 17887 9053 17901 9070
rect 17355 8957 17503 9036
rect 17355 8937 17359 8957
rect 17379 8937 17398 8957
rect 17418 8937 17437 8957
rect 17457 8937 17476 8957
rect 17496 8937 17503 8957
rect 17355 8455 17503 8937
rect 17355 8435 17359 8455
rect 17379 8435 17398 8455
rect 17418 8435 17437 8455
rect 17457 8435 17476 8455
rect 17496 8435 17503 8455
rect 17355 7953 17503 8435
rect 17355 7933 17359 7953
rect 17379 7933 17398 7953
rect 17418 7933 17437 7953
rect 17457 7933 17476 7953
rect 17496 7933 17503 7953
rect 17355 7451 17503 7933
rect 17355 7431 17359 7451
rect 17379 7431 17398 7451
rect 17418 7431 17437 7451
rect 17457 7431 17476 7451
rect 17496 7431 17503 7451
rect 17355 6949 17503 7431
rect 17355 6929 17359 6949
rect 17379 6929 17398 6949
rect 17418 6929 17437 6949
rect 17457 6929 17476 6949
rect 17496 6929 17503 6949
rect 17355 6447 17503 6929
rect 17355 6427 17359 6447
rect 17379 6427 17398 6447
rect 17418 6427 17437 6447
rect 17457 6427 17476 6447
rect 17496 6427 17503 6447
rect 17355 5945 17503 6427
rect 17355 5925 17359 5945
rect 17379 5925 17398 5945
rect 17418 5925 17437 5945
rect 17457 5925 17476 5945
rect 17496 5925 17503 5945
rect 17355 5443 17503 5925
rect 17355 5423 17359 5443
rect 17379 5423 17398 5443
rect 17418 5423 17437 5443
rect 17457 5423 17476 5443
rect 17496 5423 17503 5443
rect 17355 4941 17503 5423
rect 17355 4921 17359 4941
rect 17379 4921 17398 4941
rect 17418 4921 17437 4941
rect 17457 4921 17476 4941
rect 17496 4921 17503 4941
rect 17355 4439 17503 4921
rect 17355 4419 17359 4439
rect 17379 4419 17398 4439
rect 17418 4419 17437 4439
rect 17457 4419 17476 4439
rect 17496 4419 17503 4439
rect 17355 3937 17503 4419
rect 17355 3917 17359 3937
rect 17379 3917 17398 3937
rect 17418 3917 17437 3937
rect 17457 3917 17476 3937
rect 17496 3917 17503 3937
rect 17355 3435 17503 3917
rect 17355 3415 17359 3435
rect 17379 3415 17398 3435
rect 17418 3415 17437 3435
rect 17457 3415 17476 3435
rect 17496 3415 17503 3435
rect 17355 2933 17503 3415
rect 17355 2913 17359 2933
rect 17379 2913 17398 2933
rect 17418 2913 17437 2933
rect 17457 2913 17476 2933
rect 17496 2913 17503 2933
rect 17355 2431 17503 2913
rect 17355 2411 17359 2431
rect 17379 2411 17398 2431
rect 17418 2411 17437 2431
rect 17457 2411 17476 2431
rect 17496 2411 17503 2431
rect 17355 1929 17503 2411
rect 17355 1909 17359 1929
rect 17379 1909 17398 1929
rect 17418 1909 17437 1929
rect 17457 1909 17476 1929
rect 17496 1909 17503 1929
rect 17355 1427 17503 1909
rect 17355 1407 17359 1427
rect 17379 1407 17398 1427
rect 17418 1407 17437 1427
rect 17457 1407 17476 1427
rect 17496 1407 17503 1427
rect 17355 925 17503 1407
rect 17355 905 17359 925
rect 17379 905 17398 925
rect 17418 905 17437 925
rect 17457 905 17476 925
rect 17496 905 17503 925
rect 17355 423 17503 905
rect 17355 403 17359 423
rect 17379 403 17398 423
rect 17418 403 17437 423
rect 17457 403 17476 423
rect 17496 403 17503 423
rect 17355 -238 17503 403
rect 17545 8661 17613 9036
rect 17545 8641 17548 8661
rect 17568 8641 17587 8661
rect 17607 8641 17613 8661
rect 17545 8159 17613 8641
rect 17545 8139 17548 8159
rect 17568 8139 17587 8159
rect 17607 8139 17613 8159
rect 17545 7657 17613 8139
rect 17545 7637 17548 7657
rect 17568 7637 17587 7657
rect 17607 7637 17613 7657
rect 17545 7155 17613 7637
rect 17545 7135 17548 7155
rect 17568 7135 17587 7155
rect 17607 7135 17613 7155
rect 17545 6653 17613 7135
rect 17545 6633 17548 6653
rect 17568 6633 17587 6653
rect 17607 6633 17613 6653
rect 17545 6151 17613 6633
rect 17545 6131 17548 6151
rect 17568 6131 17587 6151
rect 17607 6131 17613 6151
rect 17545 5649 17613 6131
rect 17545 5629 17548 5649
rect 17568 5629 17587 5649
rect 17607 5629 17613 5649
rect 17545 5147 17613 5629
rect 17545 5127 17548 5147
rect 17568 5127 17587 5147
rect 17607 5127 17613 5147
rect 17545 4645 17613 5127
rect 17545 4625 17548 4645
rect 17568 4625 17587 4645
rect 17607 4625 17613 4645
rect 17545 4143 17613 4625
rect 17545 4123 17548 4143
rect 17568 4123 17587 4143
rect 17607 4123 17613 4143
rect 17545 3641 17613 4123
rect 17545 3621 17548 3641
rect 17568 3621 17587 3641
rect 17607 3621 17613 3641
rect 17545 3139 17613 3621
rect 17545 3119 17548 3139
rect 17568 3119 17587 3139
rect 17607 3119 17613 3139
rect 17545 2637 17613 3119
rect 17545 2617 17548 2637
rect 17568 2617 17587 2637
rect 17607 2617 17613 2637
rect 17545 2135 17613 2617
rect 17545 2115 17548 2135
rect 17568 2115 17587 2135
rect 17607 2115 17613 2135
rect 17545 1633 17613 2115
rect 17545 1613 17548 1633
rect 17568 1613 17587 1633
rect 17607 1613 17613 1633
rect 17545 1131 17613 1613
rect 17545 1111 17548 1131
rect 17568 1111 17587 1131
rect 17607 1111 17613 1131
rect 17545 629 17613 1111
rect 17545 609 17548 629
rect 17568 609 17587 629
rect 17607 609 17613 629
rect 17545 127 17613 609
rect 17545 107 17548 127
rect 17568 107 17587 127
rect 17607 107 17613 127
rect 17545 0 17613 107
rect 17694 9030 17901 9053
rect 17694 9013 17712 9030
rect 17887 9013 17901 9030
rect 17694 8990 17901 9013
rect 17694 8973 17712 8990
rect 17887 8973 17901 8990
rect 17694 8950 17901 8973
rect 17694 8933 17712 8950
rect 17887 8933 17901 8950
rect 17694 8910 17901 8933
rect 17694 8893 17712 8910
rect 17887 8893 17901 8910
rect 17694 8870 17901 8893
rect 17694 8853 17712 8870
rect 17887 8853 17901 8870
rect 17694 8830 17901 8853
rect 17694 8813 17712 8830
rect 17887 8813 17901 8830
rect 17694 8790 17901 8813
rect 17694 8773 17712 8790
rect 17887 8773 17901 8790
rect 17694 8750 17901 8773
rect 17694 8733 17712 8750
rect 17887 8733 17901 8750
rect 17694 8710 17901 8733
rect 17694 8693 17712 8710
rect 17887 8693 17901 8710
rect 17694 8670 17901 8693
rect 17694 8653 17712 8670
rect 17887 8653 17901 8670
rect 17694 8630 17901 8653
rect 17694 8613 17712 8630
rect 17887 8613 17901 8630
rect 17694 8590 17901 8613
rect 17694 8573 17712 8590
rect 17887 8573 17901 8590
rect 17694 8550 17901 8573
rect 17694 8533 17712 8550
rect 17887 8533 17901 8550
rect 17694 8510 17901 8533
rect 17694 8493 17712 8510
rect 17887 8493 17901 8510
rect 17694 8470 17901 8493
rect 17694 8453 17712 8470
rect 17887 8453 17901 8470
rect 17694 8430 17901 8453
rect 17694 8413 17712 8430
rect 17887 8413 17901 8430
rect 17694 8390 17901 8413
rect 17694 8373 17712 8390
rect 17887 8373 17901 8390
rect 17694 8350 17901 8373
rect 17694 8333 17712 8350
rect 17887 8333 17901 8350
rect 17694 8310 17901 8333
rect 17694 8293 17712 8310
rect 17887 8293 17901 8310
rect 17694 8270 17901 8293
rect 17694 8253 17712 8270
rect 17887 8253 17901 8270
rect 17694 8230 17901 8253
rect 17694 8213 17712 8230
rect 17887 8213 17901 8230
rect 17694 8190 17901 8213
rect 17694 8173 17712 8190
rect 17887 8173 17901 8190
rect 17694 8150 17901 8173
rect 17694 8133 17712 8150
rect 17887 8133 17901 8150
rect 17694 8110 17901 8133
rect 17694 8093 17712 8110
rect 17887 8093 17901 8110
rect 17694 8070 17901 8093
rect 17694 8053 17712 8070
rect 17887 8053 17901 8070
rect 17694 8030 17901 8053
rect 17694 8013 17712 8030
rect 17887 8013 17901 8030
rect 17694 7990 17901 8013
rect 17694 7973 17712 7990
rect 17887 7973 17901 7990
rect 17694 7950 17901 7973
rect 17694 7933 17712 7950
rect 17887 7933 17901 7950
rect 17694 7910 17901 7933
rect 17694 7893 17712 7910
rect 17887 7893 17901 7910
rect 17694 7870 17901 7893
rect 17694 7853 17712 7870
rect 17887 7853 17901 7870
rect 17694 7830 17901 7853
rect 17694 7813 17712 7830
rect 17887 7813 17901 7830
rect 17694 7790 17901 7813
rect 17694 7773 17712 7790
rect 17887 7773 17901 7790
rect 17694 7750 17901 7773
rect 17694 7733 17712 7750
rect 17887 7733 17901 7750
rect 17694 7710 17901 7733
rect 17694 7693 17712 7710
rect 17887 7693 17901 7710
rect 17694 7670 17901 7693
rect 17694 7653 17712 7670
rect 17887 7653 17901 7670
rect 17694 7630 17901 7653
rect 17694 7613 17712 7630
rect 17887 7613 17901 7630
rect 17694 7590 17901 7613
rect 17694 7573 17712 7590
rect 17887 7573 17901 7590
rect 17694 7550 17901 7573
rect 17694 7533 17712 7550
rect 17887 7533 17901 7550
rect 17694 7510 17901 7533
rect 17694 7493 17712 7510
rect 17887 7493 17901 7510
rect 17694 7470 17901 7493
rect 17694 7453 17712 7470
rect 17887 7453 17901 7470
rect 17694 7430 17901 7453
rect 17694 7413 17712 7430
rect 17887 7413 17901 7430
rect 17694 7390 17901 7413
rect 17694 7373 17712 7390
rect 17887 7373 17901 7390
rect 17694 7350 17901 7373
rect 17694 7333 17712 7350
rect 17887 7333 17901 7350
rect 17694 7310 17901 7333
rect 17694 7293 17712 7310
rect 17887 7293 17901 7310
rect 17694 7270 17901 7293
rect 17694 7253 17712 7270
rect 17887 7253 17901 7270
rect 17694 7230 17901 7253
rect 17694 7213 17712 7230
rect 17887 7213 17901 7230
rect 17694 7190 17901 7213
rect 17694 7173 17712 7190
rect 17887 7173 17901 7190
rect 17694 7150 17901 7173
rect 17694 7133 17712 7150
rect 17887 7133 17901 7150
rect 17694 7110 17901 7133
rect 17694 7093 17712 7110
rect 17887 7093 17901 7110
rect 17694 7070 17901 7093
rect 17694 7053 17712 7070
rect 17887 7053 17901 7070
rect 17694 7030 17901 7053
rect 17694 7013 17712 7030
rect 17887 7013 17901 7030
rect 17694 6990 17901 7013
rect 17694 6973 17712 6990
rect 17887 6973 17901 6990
rect 17694 6950 17901 6973
rect 17694 6933 17712 6950
rect 17887 6933 17901 6950
rect 17694 6910 17901 6933
rect 17694 6893 17712 6910
rect 17887 6893 17901 6910
rect 17694 6870 17901 6893
rect 17694 6853 17712 6870
rect 17887 6853 17901 6870
rect 17694 6830 17901 6853
rect 17694 6813 17712 6830
rect 17887 6813 17901 6830
rect 17694 6790 17901 6813
rect 17694 6773 17712 6790
rect 17887 6773 17901 6790
rect 17694 6750 17901 6773
rect 17694 6733 17712 6750
rect 17887 6733 17901 6750
rect 17694 6710 17901 6733
rect 17694 6693 17712 6710
rect 17887 6693 17901 6710
rect 17694 6670 17901 6693
rect 17694 6653 17712 6670
rect 17887 6653 17901 6670
rect 17694 6630 17901 6653
rect 17694 6613 17712 6630
rect 17887 6613 17901 6630
rect 17694 6590 17901 6613
rect 17694 6573 17712 6590
rect 17887 6573 17901 6590
rect 17694 6550 17901 6573
rect 17694 6533 17712 6550
rect 17887 6533 17901 6550
rect 17694 6510 17901 6533
rect 17694 6493 17712 6510
rect 17887 6493 17901 6510
rect 17694 6470 17901 6493
rect 17694 6453 17712 6470
rect 17887 6453 17901 6470
rect 17694 6430 17901 6453
rect 17694 6413 17712 6430
rect 17887 6413 17901 6430
rect 17694 6390 17901 6413
rect 17694 6373 17712 6390
rect 17887 6373 17901 6390
rect 17694 6350 17901 6373
rect 17694 6333 17712 6350
rect 17887 6333 17901 6350
rect 17694 6310 17901 6333
rect 17694 6293 17712 6310
rect 17887 6293 17901 6310
rect 17694 6270 17901 6293
rect 17694 6253 17712 6270
rect 17887 6253 17901 6270
rect 17694 6230 17901 6253
rect 17694 6213 17712 6230
rect 17887 6213 17901 6230
rect 17694 6190 17901 6213
rect 17694 6173 17712 6190
rect 17887 6173 17901 6190
rect 17694 6150 17901 6173
rect 17694 6133 17712 6150
rect 17887 6133 17901 6150
rect 17694 6110 17901 6133
rect 17694 6093 17712 6110
rect 17887 6093 17901 6110
rect 17694 6070 17901 6093
rect 17694 6053 17712 6070
rect 17887 6053 17901 6070
rect 17694 6030 17901 6053
rect 17694 6013 17712 6030
rect 17887 6013 17901 6030
rect 17694 5990 17901 6013
rect 17694 5973 17712 5990
rect 17887 5973 17901 5990
rect 17694 5950 17901 5973
rect 17694 5933 17712 5950
rect 17887 5933 17901 5950
rect 17694 5910 17901 5933
rect 17694 5893 17712 5910
rect 17887 5893 17901 5910
rect 17694 5870 17901 5893
rect 17694 5853 17712 5870
rect 17887 5853 17901 5870
rect 17694 5830 17901 5853
rect 17694 5813 17712 5830
rect 17887 5813 17901 5830
rect 17694 5790 17901 5813
rect 17694 5773 17712 5790
rect 17887 5773 17901 5790
rect 17694 5750 17901 5773
rect 17694 5733 17712 5750
rect 17887 5733 17901 5750
rect 17694 5710 17901 5733
rect 17694 5693 17712 5710
rect 17887 5693 17901 5710
rect 17694 5670 17901 5693
rect 17694 5653 17712 5670
rect 17887 5653 17901 5670
rect 17694 5630 17901 5653
rect 17694 5613 17712 5630
rect 17887 5613 17901 5630
rect 17694 5590 17901 5613
rect 17694 5573 17712 5590
rect 17887 5573 17901 5590
rect 17694 5550 17901 5573
rect 17694 5533 17712 5550
rect 17887 5533 17901 5550
rect 17694 5510 17901 5533
rect 17694 5493 17712 5510
rect 17887 5493 17901 5510
rect 17694 5470 17901 5493
rect 17694 5453 17712 5470
rect 17887 5453 17901 5470
rect 17694 5430 17901 5453
rect 17694 5413 17712 5430
rect 17887 5413 17901 5430
rect 17694 5390 17901 5413
rect 17694 5373 17712 5390
rect 17887 5373 17901 5390
rect 17694 5350 17901 5373
rect 17694 5333 17712 5350
rect 17887 5333 17901 5350
rect 17694 5310 17901 5333
rect 17694 5293 17712 5310
rect 17887 5293 17901 5310
rect 17694 5270 17901 5293
rect 17694 5253 17712 5270
rect 17887 5253 17901 5270
rect 17694 5230 17901 5253
rect 17694 5213 17712 5230
rect 17887 5213 17901 5230
rect 17694 5190 17901 5213
rect 17694 5173 17712 5190
rect 17887 5173 17901 5190
rect 17694 5150 17901 5173
rect 17694 5133 17712 5150
rect 17887 5133 17901 5150
rect 17694 5110 17901 5133
rect 17694 5093 17712 5110
rect 17887 5093 17901 5110
rect 17694 5070 17901 5093
rect 17694 5053 17712 5070
rect 17887 5053 17901 5070
rect 17694 5030 17901 5053
rect 17694 5013 17712 5030
rect 17887 5013 17901 5030
rect 17694 4990 17901 5013
rect 17694 4973 17712 4990
rect 17887 4973 17901 4990
rect 17694 4950 17901 4973
rect 17694 4933 17712 4950
rect 17887 4933 17901 4950
rect 17694 4910 17901 4933
rect 17694 4893 17712 4910
rect 17887 4893 17901 4910
rect 17694 4870 17901 4893
rect 17694 4853 17712 4870
rect 17887 4853 17901 4870
rect 17694 4830 17901 4853
rect 17694 4813 17712 4830
rect 17887 4813 17901 4830
rect 17694 4790 17901 4813
rect 17694 4773 17712 4790
rect 17887 4773 17901 4790
rect 17694 4750 17901 4773
rect 17694 4733 17712 4750
rect 17887 4733 17901 4750
rect 17694 4710 17901 4733
rect 17694 4693 17712 4710
rect 17887 4693 17901 4710
rect 17694 4670 17901 4693
rect 17694 4653 17712 4670
rect 17887 4653 17901 4670
rect 17694 4630 17901 4653
rect 17694 4613 17712 4630
rect 17887 4613 17901 4630
rect 17694 4590 17901 4613
rect 17694 4573 17712 4590
rect 17887 4573 17901 4590
rect 17694 4550 17901 4573
rect 17694 4533 17712 4550
rect 17887 4533 17901 4550
rect 17694 4510 17901 4533
rect 17694 4493 17712 4510
rect 17887 4493 17901 4510
rect 17694 4470 17901 4493
rect 17694 4453 17712 4470
rect 17887 4453 17901 4470
rect 17694 4430 17901 4453
rect 17694 4413 17712 4430
rect 17887 4413 17901 4430
rect 17694 4390 17901 4413
rect 17694 4373 17712 4390
rect 17887 4373 17901 4390
rect 17694 4350 17901 4373
rect 17694 4333 17712 4350
rect 17887 4333 17901 4350
rect 17694 4310 17901 4333
rect 17694 4293 17712 4310
rect 17887 4293 17901 4310
rect 17694 4270 17901 4293
rect 17694 4253 17712 4270
rect 17887 4253 17901 4270
rect 17694 4230 17901 4253
rect 17694 4213 17712 4230
rect 17887 4213 17901 4230
rect 17694 4190 17901 4213
rect 17694 4173 17712 4190
rect 17887 4173 17901 4190
rect 17694 4150 17901 4173
rect 17694 4133 17712 4150
rect 17887 4133 17901 4150
rect 17694 4110 17901 4133
rect 17694 4093 17712 4110
rect 17887 4093 17901 4110
rect 17694 4070 17901 4093
rect 17694 4053 17712 4070
rect 17887 4053 17901 4070
rect 17694 4030 17901 4053
rect 17694 4013 17712 4030
rect 17887 4013 17901 4030
rect 17694 3990 17901 4013
rect 17694 3973 17712 3990
rect 17887 3973 17901 3990
rect 17694 3950 17901 3973
rect 17694 3933 17712 3950
rect 17887 3933 17901 3950
rect 17694 3910 17901 3933
rect 17694 3893 17712 3910
rect 17887 3893 17901 3910
rect 17694 3870 17901 3893
rect 17694 3853 17712 3870
rect 17887 3853 17901 3870
rect 17694 3830 17901 3853
rect 17694 3813 17712 3830
rect 17887 3813 17901 3830
rect 17694 3790 17901 3813
rect 17694 3773 17712 3790
rect 17887 3773 17901 3790
rect 17694 3750 17901 3773
rect 17694 3733 17712 3750
rect 17887 3733 17901 3750
rect 17694 3710 17901 3733
rect 17694 3693 17712 3710
rect 17887 3693 17901 3710
rect 17694 3670 17901 3693
rect 17694 3653 17712 3670
rect 17887 3653 17901 3670
rect 17694 3630 17901 3653
rect 17694 3613 17712 3630
rect 17887 3613 17901 3630
rect 17694 3590 17901 3613
rect 17694 3573 17712 3590
rect 17887 3573 17901 3590
rect 17694 3550 17901 3573
rect 17694 3533 17712 3550
rect 17887 3533 17901 3550
rect 17694 3510 17901 3533
rect 17694 3493 17712 3510
rect 17887 3493 17901 3510
rect 17694 3470 17901 3493
rect 17694 3453 17712 3470
rect 17887 3453 17901 3470
rect 17694 3430 17901 3453
rect 17694 3413 17712 3430
rect 17887 3413 17901 3430
rect 17694 3390 17901 3413
rect 17694 3373 17712 3390
rect 17887 3373 17901 3390
rect 17694 3350 17901 3373
rect 17694 3333 17712 3350
rect 17887 3333 17901 3350
rect 17694 3310 17901 3333
rect 17694 3293 17712 3310
rect 17887 3293 17901 3310
rect 17694 3270 17901 3293
rect 17694 3253 17712 3270
rect 17887 3253 17901 3270
rect 17694 3230 17901 3253
rect 17694 3213 17712 3230
rect 17887 3213 17901 3230
rect 17694 3190 17901 3213
rect 17694 3173 17712 3190
rect 17887 3173 17901 3190
rect 17694 3150 17901 3173
rect 17694 3133 17712 3150
rect 17887 3133 17901 3150
rect 17694 3110 17901 3133
rect 17694 3093 17712 3110
rect 17887 3093 17901 3110
rect 17694 3070 17901 3093
rect 17694 3053 17712 3070
rect 17887 3053 17901 3070
rect 17694 3030 17901 3053
rect 17694 3013 17712 3030
rect 17887 3013 17901 3030
rect 17694 2990 17901 3013
rect 17694 2973 17712 2990
rect 17887 2973 17901 2990
rect 17694 2950 17901 2973
rect 17694 2933 17712 2950
rect 17887 2933 17901 2950
rect 17694 2910 17901 2933
rect 17694 2893 17712 2910
rect 17887 2893 17901 2910
rect 17694 2870 17901 2893
rect 17694 2853 17712 2870
rect 17887 2853 17901 2870
rect 17694 2830 17901 2853
rect 17694 2813 17712 2830
rect 17887 2813 17901 2830
rect 17694 2790 17901 2813
rect 17694 2773 17712 2790
rect 17887 2773 17901 2790
rect 17694 2750 17901 2773
rect 17694 2733 17712 2750
rect 17887 2733 17901 2750
rect 17694 2710 17901 2733
rect 17694 2693 17712 2710
rect 17887 2693 17901 2710
rect 17694 2670 17901 2693
rect 17694 2653 17712 2670
rect 17887 2653 17901 2670
rect 17694 2630 17901 2653
rect 17694 2613 17712 2630
rect 17887 2613 17901 2630
rect 17694 2590 17901 2613
rect 17694 2573 17712 2590
rect 17887 2573 17901 2590
rect 17694 2550 17901 2573
rect 17694 2533 17712 2550
rect 17887 2533 17901 2550
rect 17694 2510 17901 2533
rect 17694 2493 17712 2510
rect 17887 2493 17901 2510
rect 17694 2470 17901 2493
rect 17694 2453 17712 2470
rect 17887 2453 17901 2470
rect 17694 2430 17901 2453
rect 17694 2413 17712 2430
rect 17887 2413 17901 2430
rect 17694 2390 17901 2413
rect 17694 2373 17712 2390
rect 17887 2373 17901 2390
rect 17694 2350 17901 2373
rect 17694 2333 17712 2350
rect 17887 2333 17901 2350
rect 17694 2310 17901 2333
rect 17694 2293 17712 2310
rect 17887 2293 17901 2310
rect 17694 2270 17901 2293
rect 17694 2253 17712 2270
rect 17887 2253 17901 2270
rect 17694 2230 17901 2253
rect 17694 2213 17712 2230
rect 17887 2213 17901 2230
rect 17694 2190 17901 2213
rect 17694 2173 17712 2190
rect 17887 2173 17901 2190
rect 17694 2150 17901 2173
rect 17694 2133 17712 2150
rect 17887 2133 17901 2150
rect 17694 2110 17901 2133
rect 17694 2093 17712 2110
rect 17887 2093 17901 2110
rect 17694 2070 17901 2093
rect 17694 2053 17712 2070
rect 17887 2053 17901 2070
rect 17694 2030 17901 2053
rect 17694 2013 17712 2030
rect 17887 2013 17901 2030
rect 17694 1990 17901 2013
rect 17694 1973 17712 1990
rect 17887 1973 17901 1990
rect 17694 1950 17901 1973
rect 17694 1933 17712 1950
rect 17887 1933 17901 1950
rect 17694 1910 17901 1933
rect 17694 1893 17712 1910
rect 17887 1893 17901 1910
rect 17694 1870 17901 1893
rect 17694 1853 17712 1870
rect 17887 1853 17901 1870
rect 17694 1830 17901 1853
rect 17694 1813 17712 1830
rect 17887 1813 17901 1830
rect 17694 1790 17901 1813
rect 17694 1773 17712 1790
rect 17887 1773 17901 1790
rect 17694 1750 17901 1773
rect 17694 1733 17712 1750
rect 17887 1733 17901 1750
rect 17694 1710 17901 1733
rect 17694 1693 17712 1710
rect 17887 1693 17901 1710
rect 17694 1670 17901 1693
rect 17694 1653 17712 1670
rect 17887 1653 17901 1670
rect 17694 1630 17901 1653
rect 17694 1613 17712 1630
rect 17887 1613 17901 1630
rect 17694 1590 17901 1613
rect 17694 1573 17712 1590
rect 17887 1573 17901 1590
rect 17694 1550 17901 1573
rect 17694 1533 17712 1550
rect 17887 1533 17901 1550
rect 17694 1510 17901 1533
rect 17694 1493 17712 1510
rect 17887 1493 17901 1510
rect 17694 1470 17901 1493
rect 17694 1453 17712 1470
rect 17887 1453 17901 1470
rect 17694 1430 17901 1453
rect 17694 1413 17712 1430
rect 17887 1413 17901 1430
rect 17694 1390 17901 1413
rect 17694 1373 17712 1390
rect 17887 1373 17901 1390
rect 17694 1350 17901 1373
rect 17694 1333 17712 1350
rect 17887 1333 17901 1350
rect 17694 1310 17901 1333
rect 17694 1293 17712 1310
rect 17887 1293 17901 1310
rect 17694 1270 17901 1293
rect 17694 1253 17712 1270
rect 17887 1253 17901 1270
rect 17694 1230 17901 1253
rect 17694 1213 17712 1230
rect 17887 1213 17901 1230
rect 17694 1190 17901 1213
rect 17694 1173 17712 1190
rect 17887 1173 17901 1190
rect 17694 1150 17901 1173
rect 17694 1133 17712 1150
rect 17887 1133 17901 1150
rect 17694 1110 17901 1133
rect 17694 1093 17712 1110
rect 17887 1093 17901 1110
rect 17694 1070 17901 1093
rect 17694 1053 17712 1070
rect 17887 1053 17901 1070
rect 17694 1030 17901 1053
rect 17694 1013 17712 1030
rect 17887 1013 17901 1030
rect 17694 990 17901 1013
rect 17694 973 17712 990
rect 17887 973 17901 990
rect 17694 950 17901 973
rect 17694 933 17712 950
rect 17887 933 17901 950
rect 17694 910 17901 933
rect 17694 893 17712 910
rect 17887 893 17901 910
rect 17694 870 17901 893
rect 17694 853 17712 870
rect 17887 853 17901 870
rect 17694 830 17901 853
rect 17694 813 17712 830
rect 17887 813 17901 830
rect 17694 790 17901 813
rect 17694 773 17712 790
rect 17887 773 17901 790
rect 17694 750 17901 773
rect 17694 733 17712 750
rect 17887 733 17901 750
rect 17694 710 17901 733
rect 17694 693 17712 710
rect 17887 693 17901 710
rect 17694 670 17901 693
rect 17694 653 17712 670
rect 17887 653 17901 670
rect 17694 630 17901 653
rect 17694 613 17712 630
rect 17887 613 17901 630
rect 17694 590 17901 613
rect 17694 573 17712 590
rect 17887 573 17901 590
rect 17694 550 17901 573
rect 17694 533 17712 550
rect 17887 533 17901 550
rect 17694 510 17901 533
rect 17694 493 17712 510
rect 17887 493 17901 510
rect 17694 470 17901 493
rect 17694 453 17712 470
rect 17887 453 17901 470
rect 17694 430 17901 453
rect 17694 413 17712 430
rect 17887 413 17901 430
rect 17694 390 17901 413
rect 17694 373 17712 390
rect 17887 373 17901 390
rect 17694 350 17901 373
rect 17694 333 17712 350
rect 17887 333 17901 350
rect 17694 310 17901 333
rect 17694 293 17712 310
rect 17887 293 17901 310
rect 17694 270 17901 293
rect 17694 253 17712 270
rect 17887 253 17901 270
rect 17694 230 17901 253
rect 17694 213 17712 230
rect 17887 213 17901 230
rect 17694 190 17901 213
rect 17694 173 17712 190
rect 17887 173 17901 190
rect 17694 150 17901 173
rect 17694 133 17712 150
rect 17887 133 17901 150
rect 17694 110 17901 133
rect 17694 93 17712 110
rect 17887 93 17901 110
rect 17694 70 17901 93
rect 17694 53 17712 70
rect 17887 53 17901 70
rect 17694 30 17901 53
rect 17694 13 17712 30
rect 17887 13 17901 30
rect 17694 -152 17901 13
rect 17355 -266 17370 -238
rect 17398 -266 17417 -238
rect 17445 -266 17464 -238
rect 17492 -266 17503 -238
rect 17355 -285 17503 -266
rect 17355 -313 17370 -285
rect 17398 -313 17417 -285
rect 17445 -313 17464 -285
rect 17492 -313 17503 -285
rect 17355 -332 17503 -313
rect 17355 -360 17370 -332
rect 17398 -360 17417 -332
rect 17445 -360 17464 -332
rect 17492 -360 17503 -332
rect 17355 -392 17503 -360
rect 17989 -371 18196 9493
rect 16437 -432 16454 -429
rect 16395 -449 16401 -432
rect 16418 -449 16437 -432
rect 16454 -449 16460 -432
rect 16401 -456 16418 -449
rect 16437 -453 16454 -449
<< viali >>
rect -430 9455 -402 9483
rect -383 9455 -355 9483
rect -336 9455 -308 9483
rect -430 9408 -402 9436
rect -383 9408 -355 9436
rect -336 9408 -308 9436
rect -430 9361 -402 9389
rect -383 9361 -355 9389
rect -336 9361 -308 9389
rect -2143 8853 -1968 8870
rect -2143 8413 -1968 8430
rect -651 8407 -634 8424
rect -2143 7973 -1968 7990
rect -1373 8285 -1356 8302
rect -2143 7533 -1968 7550
rect -1409 7786 -1392 7803
rect -2143 7093 -1968 7110
rect -1445 7283 -1428 7300
rect -2143 6653 -1968 6670
rect -1481 6780 -1464 6797
rect -2143 6213 -1968 6230
rect -1517 6280 -1500 6297
rect -2143 5773 -1968 5790
rect -2143 5333 -1968 5350
rect -1553 5778 -1536 5795
rect -2143 4893 -1968 4910
rect -1589 5276 -1572 5293
rect -2143 4453 -1968 4470
rect -1625 4773 -1608 4790
rect -2143 4013 -1968 4030
rect -1661 4272 -1644 4289
rect -2143 3573 -1968 3590
rect -1697 3770 -1680 3787
rect -2143 3133 -1968 3150
rect -1733 3268 -1716 3285
rect -2143 2693 -1968 2710
rect -1769 2766 -1752 2783
rect -2143 2253 -1968 2270
rect -2143 1813 -1968 1830
rect -1805 2265 -1788 2282
rect -2143 1373 -1968 1390
rect -1841 1762 -1824 1779
rect -2143 933 -1968 950
rect -1877 1259 -1860 1276
rect -2143 493 -1968 510
rect -2143 53 -1968 70
rect -1913 758 -1896 775
rect -761 8244 -744 8261
rect -797 7742 -780 7759
rect -833 7242 -816 7259
rect -869 6740 -852 6757
rect -905 6239 -888 6256
rect -941 5735 -924 5752
rect -977 5235 -960 5252
rect -1013 4732 -996 4749
rect -1049 4233 -1032 4250
rect -1085 3730 -1068 3747
rect -1121 3228 -1104 3245
rect -1157 2727 -1140 2744
rect -1193 2222 -1176 2239
rect -1229 1719 -1212 1736
rect -1265 1216 -1248 1233
rect -1301 718 -1284 735
rect -651 7905 -634 7922
rect -651 7403 -634 7420
rect -651 6901 -634 6918
rect -651 6399 -634 6416
rect -651 5897 -634 5914
rect -651 5395 -634 5412
rect -651 4893 -634 4910
rect -651 4391 -634 4408
rect -651 3889 -634 3906
rect -651 3387 -634 3404
rect -651 2885 -634 2902
rect -651 2383 -634 2400
rect -651 1881 -634 1898
rect -651 1379 -634 1396
rect -651 877 -634 894
rect -597 8213 -580 8230
rect -597 7711 -580 7728
rect -597 7209 -580 7226
rect -597 6707 -580 6724
rect -597 6205 -580 6222
rect -597 5703 -580 5720
rect -597 5201 -580 5218
rect -597 4699 -580 4716
rect -597 4197 -580 4214
rect -597 3695 -580 3712
rect -597 3193 -580 3210
rect -597 2691 -580 2708
rect -597 2189 -580 2206
rect -597 1687 -580 1704
rect -597 1185 -580 1202
rect -597 683 -580 700
rect -545 8641 -525 8661
rect -506 8641 -486 8661
rect -545 8139 -525 8159
rect -506 8139 -486 8159
rect -545 7637 -525 7657
rect -506 7637 -486 7657
rect -545 7135 -525 7155
rect -506 7135 -486 7155
rect -545 6633 -525 6653
rect -506 6633 -486 6653
rect -545 6131 -525 6151
rect -506 6131 -486 6151
rect -545 5629 -525 5649
rect -506 5629 -486 5649
rect -545 5127 -525 5147
rect -506 5127 -486 5147
rect -545 4625 -525 4645
rect -506 4625 -486 4645
rect -545 4123 -525 4143
rect -506 4123 -486 4143
rect -545 3621 -525 3641
rect -506 3621 -486 3641
rect -545 3119 -525 3139
rect -506 3119 -486 3139
rect -545 2617 -525 2637
rect -506 2617 -486 2637
rect -545 2115 -525 2135
rect -506 2115 -486 2135
rect -545 1613 -525 1633
rect -506 1613 -486 1633
rect -545 1111 -525 1131
rect -506 1111 -486 1131
rect -545 609 -525 629
rect -506 609 -486 629
rect -545 107 -525 127
rect -506 107 -486 127
rect -434 8937 -414 8957
rect -395 8937 -375 8957
rect -356 8937 -336 8957
rect -317 8937 -297 8957
rect -434 8895 -414 8915
rect -395 8895 -375 8915
rect -356 8895 -336 8915
rect -317 8895 -297 8915
rect -434 8767 -414 8787
rect -395 8767 -375 8787
rect -356 8767 -336 8787
rect -317 8767 -297 8787
rect -434 8435 -414 8455
rect -395 8435 -375 8455
rect -356 8435 -336 8455
rect -317 8435 -297 8455
rect -434 7933 -414 7953
rect -395 7933 -375 7953
rect -356 7933 -336 7953
rect -317 7933 -297 7953
rect -434 7431 -414 7451
rect -395 7431 -375 7451
rect -356 7431 -336 7451
rect -317 7431 -297 7451
rect -434 6929 -414 6949
rect -395 6929 -375 6949
rect -356 6929 -336 6949
rect -317 6929 -297 6949
rect -434 6427 -414 6447
rect -395 6427 -375 6447
rect -356 6427 -336 6447
rect -317 6427 -297 6447
rect -434 5925 -414 5945
rect -395 5925 -375 5945
rect -356 5925 -336 5945
rect -317 5925 -297 5945
rect -434 5423 -414 5443
rect -395 5423 -375 5443
rect -356 5423 -336 5443
rect -317 5423 -297 5443
rect -434 4921 -414 4941
rect -395 4921 -375 4941
rect -356 4921 -336 4941
rect -317 4921 -297 4941
rect -434 4419 -414 4439
rect -395 4419 -375 4439
rect -356 4419 -336 4439
rect -317 4419 -297 4439
rect -434 3917 -414 3937
rect -395 3917 -375 3937
rect -356 3917 -336 3937
rect -317 3917 -297 3937
rect -434 3415 -414 3435
rect -395 3415 -375 3435
rect -356 3415 -336 3435
rect -317 3415 -297 3435
rect -434 2913 -414 2933
rect -395 2913 -375 2933
rect -356 2913 -336 2933
rect -317 2913 -297 2933
rect -434 2411 -414 2431
rect -395 2411 -375 2431
rect -356 2411 -336 2431
rect -317 2411 -297 2431
rect -434 1909 -414 1929
rect -395 1909 -375 1929
rect -356 1909 -336 1929
rect -317 1909 -297 1929
rect -434 1407 -414 1427
rect -395 1407 -375 1427
rect -356 1407 -336 1427
rect -317 1407 -297 1427
rect -434 905 -414 925
rect -395 905 -375 925
rect -356 905 -336 925
rect -317 905 -297 925
rect -434 403 -414 423
rect -395 403 -375 423
rect -356 403 -336 423
rect -317 403 -297 423
rect -434 361 -414 381
rect -395 361 -375 381
rect -356 361 -336 381
rect -317 361 -297 381
rect -430 -332 -402 -304
rect -383 -332 -355 -304
rect -336 -332 -308 -304
rect -430 -379 -402 -351
rect -383 -379 -355 -351
rect -336 -379 -308 -351
rect -430 -426 -402 -398
rect -383 -426 -355 -398
rect -336 -426 -308 -398
rect -241 9236 -213 9264
rect -194 9236 -166 9264
rect -147 9236 -119 9264
rect -241 9189 -213 9217
rect -194 9189 -166 9217
rect -147 9189 -119 9217
rect -241 9142 -213 9170
rect -194 9142 -166 9170
rect -147 9142 -119 9170
rect -245 8711 -225 8731
rect -206 8711 -186 8731
rect -167 8711 -147 8731
rect -128 8711 -108 8731
rect -245 8606 -225 8626
rect -206 8606 -186 8626
rect -167 8606 -147 8626
rect -128 8606 -108 8626
rect -245 8104 -225 8124
rect -206 8104 -186 8124
rect -167 8104 -147 8124
rect -128 8104 -108 8124
rect -245 7602 -225 7622
rect -206 7602 -186 7622
rect -167 7602 -147 7622
rect -128 7602 -108 7622
rect -245 7100 -225 7120
rect -206 7100 -186 7120
rect -167 7100 -147 7120
rect -128 7100 -108 7120
rect -245 6598 -225 6618
rect -206 6598 -186 6618
rect -167 6598 -147 6618
rect -128 6598 -108 6618
rect -245 6096 -225 6116
rect -206 6096 -186 6116
rect -167 6096 -147 6116
rect -128 6096 -108 6116
rect -245 5594 -225 5614
rect -206 5594 -186 5614
rect -167 5594 -147 5614
rect -128 5594 -108 5614
rect -245 5092 -225 5112
rect -206 5092 -186 5112
rect -167 5092 -147 5112
rect -128 5092 -108 5112
rect -245 4590 -225 4610
rect -206 4590 -186 4610
rect -167 4590 -147 4610
rect -128 4590 -108 4610
rect -245 4088 -225 4108
rect -206 4088 -186 4108
rect -167 4088 -147 4108
rect -128 4088 -108 4108
rect -245 3586 -225 3606
rect -206 3586 -186 3606
rect -167 3586 -147 3606
rect -128 3586 -108 3606
rect -245 3084 -225 3104
rect -206 3084 -186 3104
rect -167 3084 -147 3104
rect -128 3084 -108 3104
rect -245 2582 -225 2602
rect -206 2582 -186 2602
rect -167 2582 -147 2602
rect -128 2582 -108 2602
rect -245 2080 -225 2100
rect -206 2080 -186 2100
rect -167 2080 -147 2100
rect -128 2080 -108 2100
rect -245 1578 -225 1598
rect -206 1578 -186 1598
rect -167 1578 -147 1598
rect -128 1578 -108 1598
rect -245 1076 -225 1096
rect -206 1076 -186 1096
rect -167 1076 -147 1096
rect -128 1076 -108 1096
rect -245 574 -225 594
rect -206 574 -186 594
rect -167 574 -147 594
rect -128 574 -108 594
rect -245 233 -225 253
rect -206 233 -186 253
rect -167 233 -147 253
rect -128 233 -108 253
rect -245 177 -225 197
rect -206 177 -186 197
rect -167 177 -147 197
rect -128 177 -108 197
rect -245 72 -225 92
rect -206 72 -186 92
rect -167 72 -147 92
rect -128 72 -108 92
rect 17181 9231 17209 9259
rect 17228 9231 17256 9259
rect 17275 9231 17303 9259
rect 17181 9184 17209 9212
rect 17228 9184 17256 9212
rect 17275 9184 17303 9212
rect 17181 9137 17209 9165
rect 17228 9137 17256 9165
rect 17275 9137 17303 9165
rect 17170 8606 17190 8626
rect 17209 8606 17229 8626
rect 17248 8606 17268 8626
rect 17287 8606 17307 8626
rect 17170 8104 17190 8124
rect 17209 8104 17229 8124
rect 17248 8104 17268 8124
rect 17287 8104 17307 8124
rect 17170 7602 17190 7622
rect 17209 7602 17229 7622
rect 17248 7602 17268 7622
rect 17287 7602 17307 7622
rect 17170 7100 17190 7120
rect 17209 7100 17229 7120
rect 17248 7100 17268 7120
rect 17287 7100 17307 7120
rect 17170 6598 17190 6618
rect 17209 6598 17229 6618
rect 17248 6598 17268 6618
rect 17287 6598 17307 6618
rect 17170 6096 17190 6116
rect 17209 6096 17229 6116
rect 17248 6096 17268 6116
rect 17287 6096 17307 6116
rect 17170 5594 17190 5614
rect 17209 5594 17229 5614
rect 17248 5594 17268 5614
rect 17287 5594 17307 5614
rect 17170 5092 17190 5112
rect 17209 5092 17229 5112
rect 17248 5092 17268 5112
rect 17287 5092 17307 5112
rect 17170 4590 17190 4610
rect 17209 4590 17229 4610
rect 17248 4590 17268 4610
rect 17287 4590 17307 4610
rect 17170 4088 17190 4108
rect 17209 4088 17229 4108
rect 17248 4088 17268 4108
rect 17287 4088 17307 4108
rect 17170 3586 17190 3606
rect 17209 3586 17229 3606
rect 17248 3586 17268 3606
rect 17287 3586 17307 3606
rect 17170 3084 17190 3104
rect 17209 3084 17229 3104
rect 17248 3084 17268 3104
rect 17287 3084 17307 3104
rect 17170 2582 17190 2602
rect 17209 2582 17229 2602
rect 17248 2582 17268 2602
rect 17287 2582 17307 2602
rect 17170 2080 17190 2100
rect 17209 2080 17229 2100
rect 17248 2080 17268 2100
rect 17287 2080 17307 2100
rect 17170 1578 17190 1598
rect 17209 1578 17229 1598
rect 17248 1578 17268 1598
rect 17287 1578 17307 1598
rect 17170 1076 17190 1096
rect 17209 1076 17229 1096
rect 17248 1076 17268 1096
rect 17287 1076 17307 1096
rect 17170 574 17190 594
rect 17209 574 17229 594
rect 17248 574 17268 594
rect 17287 574 17307 594
rect 17170 72 17190 92
rect 17209 72 17229 92
rect 17248 72 17268 92
rect 17287 72 17307 92
rect -241 -113 -213 -85
rect -194 -113 -166 -85
rect -147 -113 -119 -85
rect -241 -160 -213 -132
rect -194 -160 -166 -132
rect -147 -160 -119 -132
rect -241 -207 -213 -179
rect -194 -207 -166 -179
rect -147 -207 -119 -179
rect 425 -312 442 -295
rect 13283 -153 13300 -136
rect 14483 -153 14500 -136
rect 13385 -192 13402 -175
rect 14985 -192 15002 -175
rect 13487 -230 13504 -213
rect 15487 -230 15504 -213
rect 13589 -268 13606 -251
rect 15989 -268 16006 -251
rect 13691 -306 13708 -289
rect 16104 -81 16121 -64
rect 16348 -81 16365 -64
rect 16491 -306 16508 -289
rect 17181 -48 17209 -20
rect 17228 -48 17256 -20
rect 17275 -48 17303 -20
rect 17181 -95 17209 -67
rect 17228 -95 17256 -67
rect 17275 -95 17303 -67
rect 17181 -142 17209 -114
rect 17228 -142 17256 -114
rect 17275 -142 17303 -114
rect 16995 -315 17012 -298
rect 17370 9450 17398 9478
rect 17417 9450 17445 9478
rect 17464 9450 17492 9478
rect 17370 9403 17398 9431
rect 17417 9403 17445 9431
rect 17464 9403 17492 9431
rect 17370 9356 17398 9384
rect 17417 9356 17445 9384
rect 17464 9356 17492 9384
rect 17359 8937 17379 8957
rect 17398 8937 17418 8957
rect 17437 8937 17457 8957
rect 17476 8937 17496 8957
rect 17359 8435 17379 8455
rect 17398 8435 17418 8455
rect 17437 8435 17457 8455
rect 17476 8435 17496 8455
rect 17359 7933 17379 7953
rect 17398 7933 17418 7953
rect 17437 7933 17457 7953
rect 17476 7933 17496 7953
rect 17359 7431 17379 7451
rect 17398 7431 17418 7451
rect 17437 7431 17457 7451
rect 17476 7431 17496 7451
rect 17359 6929 17379 6949
rect 17398 6929 17418 6949
rect 17437 6929 17457 6949
rect 17476 6929 17496 6949
rect 17359 6427 17379 6447
rect 17398 6427 17418 6447
rect 17437 6427 17457 6447
rect 17476 6427 17496 6447
rect 17359 5925 17379 5945
rect 17398 5925 17418 5945
rect 17437 5925 17457 5945
rect 17476 5925 17496 5945
rect 17359 5423 17379 5443
rect 17398 5423 17418 5443
rect 17437 5423 17457 5443
rect 17476 5423 17496 5443
rect 17359 4921 17379 4941
rect 17398 4921 17418 4941
rect 17437 4921 17457 4941
rect 17476 4921 17496 4941
rect 17359 4419 17379 4439
rect 17398 4419 17418 4439
rect 17437 4419 17457 4439
rect 17476 4419 17496 4439
rect 17359 3917 17379 3937
rect 17398 3917 17418 3937
rect 17437 3917 17457 3937
rect 17476 3917 17496 3937
rect 17359 3415 17379 3435
rect 17398 3415 17418 3435
rect 17437 3415 17457 3435
rect 17476 3415 17496 3435
rect 17359 2913 17379 2933
rect 17398 2913 17418 2933
rect 17437 2913 17457 2933
rect 17476 2913 17496 2933
rect 17359 2411 17379 2431
rect 17398 2411 17418 2431
rect 17437 2411 17457 2431
rect 17476 2411 17496 2431
rect 17359 1909 17379 1929
rect 17398 1909 17418 1929
rect 17437 1909 17457 1929
rect 17476 1909 17496 1929
rect 17359 1407 17379 1427
rect 17398 1407 17418 1427
rect 17437 1407 17457 1427
rect 17476 1407 17496 1427
rect 17359 905 17379 925
rect 17398 905 17418 925
rect 17437 905 17457 925
rect 17476 905 17496 925
rect 17359 403 17379 423
rect 17398 403 17418 423
rect 17437 403 17457 423
rect 17476 403 17496 423
rect 17548 8641 17568 8661
rect 17587 8641 17607 8661
rect 17548 8139 17568 8159
rect 17587 8139 17607 8159
rect 17548 7637 17568 7657
rect 17587 7637 17607 7657
rect 17548 7135 17568 7155
rect 17587 7135 17607 7155
rect 17548 6633 17568 6653
rect 17587 6633 17607 6653
rect 17548 6131 17568 6151
rect 17587 6131 17607 6151
rect 17548 5629 17568 5649
rect 17587 5629 17607 5649
rect 17548 5127 17568 5147
rect 17587 5127 17607 5147
rect 17548 4625 17568 4645
rect 17587 4625 17607 4645
rect 17548 4123 17568 4143
rect 17587 4123 17607 4143
rect 17548 3621 17568 3641
rect 17587 3621 17607 3641
rect 17548 3119 17568 3139
rect 17587 3119 17607 3139
rect 17548 2617 17568 2637
rect 17587 2617 17607 2637
rect 17548 2115 17568 2135
rect 17587 2115 17607 2135
rect 17548 1613 17568 1633
rect 17587 1613 17607 1633
rect 17548 1111 17568 1131
rect 17587 1111 17607 1131
rect 17548 609 17568 629
rect 17587 609 17607 629
rect 17548 107 17568 127
rect 17587 107 17607 127
rect 17712 8853 17887 8870
rect 17712 8413 17887 8430
rect 17712 7973 17887 7990
rect 17712 7533 17887 7550
rect 17712 7093 17887 7110
rect 17712 6653 17887 6670
rect 17712 6213 17887 6230
rect 17712 5773 17887 5790
rect 17712 5333 17887 5350
rect 17712 4893 17887 4910
rect 17712 4453 17887 4470
rect 17712 4013 17887 4030
rect 17712 3573 17887 3590
rect 17712 3133 17887 3150
rect 17712 2693 17887 2710
rect 17712 2253 17887 2270
rect 17712 1813 17887 1830
rect 17712 1373 17887 1390
rect 17712 933 17887 950
rect 17712 493 17887 510
rect 17712 53 17887 70
rect 17370 -266 17398 -238
rect 17417 -266 17445 -238
rect 17464 -266 17492 -238
rect 17370 -313 17398 -285
rect 17417 -313 17445 -285
rect 17464 -313 17492 -285
rect 17370 -360 17398 -332
rect 17417 -360 17445 -332
rect 17464 -360 17492 -332
rect 16401 -449 16418 -432
rect 16437 -449 16454 -432
<< metal1 >>
rect -2452 9489 18196 9493
rect -2452 9457 -2437 9489
rect -2405 9457 -2393 9489
rect -2361 9457 -2349 9489
rect -2317 9457 -2305 9489
rect -2273 9483 18017 9489
rect -2273 9457 -430 9483
rect -2452 9455 -430 9457
rect -402 9455 -383 9483
rect -355 9455 -336 9483
rect -308 9478 18017 9483
rect -308 9455 17370 9478
rect -2452 9450 17370 9455
rect 17398 9450 17417 9478
rect 17445 9450 17464 9478
rect 17492 9457 18017 9478
rect 18049 9457 18061 9489
rect 18093 9457 18105 9489
rect 18137 9457 18149 9489
rect 18181 9457 18196 9489
rect 17492 9450 18196 9457
rect -2452 9444 18196 9450
rect -2452 9412 -2437 9444
rect -2405 9412 -2393 9444
rect -2361 9412 -2349 9444
rect -2317 9412 -2305 9444
rect -2273 9436 18017 9444
rect -2273 9412 -430 9436
rect -2452 9408 -430 9412
rect -402 9408 -383 9436
rect -355 9408 -336 9436
rect -308 9431 18017 9436
rect -308 9408 17370 9431
rect -2452 9403 17370 9408
rect 17398 9403 17417 9431
rect 17445 9403 17464 9431
rect 17492 9412 18017 9431
rect 18049 9412 18061 9444
rect 18093 9412 18105 9444
rect 18137 9412 18149 9444
rect 18181 9412 18196 9444
rect 17492 9403 18196 9412
rect -2452 9399 18196 9403
rect -2452 9367 -2437 9399
rect -2405 9367 -2393 9399
rect -2361 9367 -2349 9399
rect -2317 9367 -2305 9399
rect -2273 9389 18017 9399
rect -2273 9367 -430 9389
rect -2452 9361 -430 9367
rect -402 9361 -383 9389
rect -355 9361 -336 9389
rect -308 9384 18017 9389
rect -308 9361 17370 9384
rect -2452 9356 17370 9361
rect 17398 9356 17417 9384
rect 17445 9356 17464 9384
rect 17492 9367 18017 9384
rect 18049 9367 18061 9399
rect 18093 9367 18105 9399
rect 18137 9367 18149 9399
rect 18181 9367 18196 9399
rect 17492 9356 18196 9367
rect -2452 9353 18196 9356
rect 17166 9348 17502 9353
rect -2157 9270 17901 9274
rect -2157 9238 -2142 9270
rect -2110 9238 -2098 9270
rect -2066 9238 -2054 9270
rect -2022 9238 -2010 9270
rect -1978 9264 17722 9270
rect -1978 9238 -241 9264
rect -2157 9236 -241 9238
rect -213 9236 -194 9264
rect -166 9236 -147 9264
rect -119 9259 17722 9264
rect -119 9236 17181 9259
rect -2157 9231 17181 9236
rect 17209 9231 17228 9259
rect 17256 9231 17275 9259
rect 17303 9238 17722 9259
rect 17754 9238 17766 9270
rect 17798 9238 17810 9270
rect 17842 9238 17854 9270
rect 17886 9238 17901 9270
rect 17303 9231 17901 9238
rect -2157 9225 17901 9231
rect -2157 9193 -2142 9225
rect -2110 9193 -2098 9225
rect -2066 9193 -2054 9225
rect -2022 9193 -2010 9225
rect -1978 9217 17722 9225
rect -1978 9193 -241 9217
rect -2157 9189 -241 9193
rect -213 9189 -194 9217
rect -166 9189 -147 9217
rect -119 9212 17722 9217
rect -119 9189 17181 9212
rect -2157 9184 17181 9189
rect 17209 9184 17228 9212
rect 17256 9184 17275 9212
rect 17303 9193 17722 9212
rect 17754 9193 17766 9225
rect 17798 9193 17810 9225
rect 17842 9193 17854 9225
rect 17886 9193 17901 9225
rect 17303 9184 17901 9193
rect -2157 9180 17901 9184
rect -2157 9148 -2142 9180
rect -2110 9148 -2098 9180
rect -2066 9148 -2054 9180
rect -2022 9148 -2010 9180
rect -1978 9170 17722 9180
rect -1978 9148 -241 9170
rect -2157 9142 -241 9148
rect -213 9142 -194 9170
rect -166 9142 -147 9170
rect -119 9165 17722 9170
rect -119 9142 17181 9165
rect -2157 9137 17181 9142
rect 17209 9137 17228 9165
rect 17256 9137 17275 9165
rect 17303 9148 17722 9165
rect 17754 9148 17766 9180
rect 17798 9148 17810 9180
rect 17842 9148 17854 9180
rect 17886 9148 17901 9180
rect 17303 9137 17901 9148
rect -2157 9135 17901 9137
rect -2156 9134 17900 9135
rect 17166 9129 17502 9134
rect -440 8957 0 8961
rect -440 8937 -434 8957
rect -414 8937 -395 8957
rect -375 8937 -356 8957
rect -336 8937 -317 8957
rect -297 8937 0 8957
rect -440 8933 0 8937
rect 17068 8957 17503 8961
rect 17068 8937 17359 8957
rect 17379 8937 17398 8957
rect 17418 8937 17437 8957
rect 17457 8937 17476 8957
rect 17496 8937 17503 8957
rect 17068 8933 17503 8937
rect -440 8915 0 8919
rect -440 8895 -434 8915
rect -414 8895 -395 8915
rect -375 8895 -356 8915
rect -336 8895 -317 8915
rect -297 8905 0 8915
rect -297 8895 -291 8905
rect -440 8891 -291 8895
rect -2149 8848 -2143 8874
rect -1968 8848 -1962 8874
rect 17706 8848 17712 8874
rect 17887 8848 17893 8874
rect -440 8790 0 8804
rect -440 8787 -291 8790
rect -440 8767 -434 8787
rect -414 8767 -395 8787
rect -375 8767 -356 8787
rect -336 8767 -317 8787
rect -297 8767 -291 8787
rect -440 8763 -291 8767
rect -440 8749 0 8763
rect -251 8731 0 8735
rect -251 8711 -245 8731
rect -225 8711 -206 8731
rect -186 8711 -167 8731
rect -147 8711 -128 8731
rect -108 8721 0 8731
rect -108 8711 -102 8721
rect -251 8707 -102 8711
rect -551 8661 -465 8664
rect -551 8641 -545 8661
rect -525 8641 -506 8661
rect -486 8658 -465 8661
rect 17527 8661 17613 8664
rect 17527 8658 17548 8661
rect -486 8644 0 8658
rect 17068 8644 17548 8658
rect -486 8641 -465 8644
rect -551 8638 -465 8641
rect 17527 8641 17548 8644
rect 17568 8641 17587 8661
rect 17607 8641 17613 8661
rect 17527 8638 17613 8641
rect -251 8626 0 8630
rect -251 8606 -245 8626
rect -225 8606 -206 8626
rect -186 8606 -167 8626
rect -147 8606 -128 8626
rect -108 8606 0 8626
rect -251 8602 0 8606
rect 17068 8626 17313 8630
rect 17068 8606 17170 8626
rect 17190 8606 17209 8626
rect 17229 8606 17248 8626
rect 17268 8606 17287 8626
rect 17307 8606 17313 8626
rect 17068 8602 17313 8606
rect -440 8455 0 8459
rect -440 8435 -434 8455
rect -414 8435 -395 8455
rect -375 8435 -356 8455
rect -336 8435 -317 8455
rect -297 8435 0 8455
rect -2149 8408 -2143 8434
rect -1968 8408 -1962 8434
rect -440 8431 0 8435
rect 17068 8455 17503 8459
rect 17068 8435 17359 8455
rect 17379 8435 17398 8455
rect 17418 8435 17437 8455
rect 17457 8435 17476 8455
rect 17496 8435 17503 8455
rect 17068 8431 17503 8435
rect -659 8424 -625 8427
rect -659 8407 -651 8424
rect -634 8417 -625 8424
rect -634 8407 0 8417
rect 17706 8408 17712 8434
rect 17887 8408 17893 8434
rect -659 8403 0 8407
rect -1376 8302 -1353 8308
rect -1376 8285 -1373 8302
rect -1356 8288 0 8302
rect -1356 8285 -1353 8288
rect -1376 8279 -1353 8285
rect -764 8261 -741 8267
rect -764 8244 -761 8261
rect -744 8247 0 8261
rect -744 8244 -741 8247
rect -764 8238 -741 8244
rect -605 8230 0 8233
rect -605 8213 -597 8230
rect -580 8219 0 8230
rect -580 8213 -571 8219
rect -605 8209 -571 8213
rect -551 8159 -465 8162
rect -551 8139 -545 8159
rect -525 8139 -506 8159
rect -486 8156 -465 8159
rect 17527 8159 17613 8162
rect 17527 8156 17548 8159
rect -486 8142 0 8156
rect 17068 8142 17548 8156
rect -486 8139 -465 8142
rect -551 8136 -465 8139
rect 17527 8139 17548 8142
rect 17568 8139 17587 8159
rect 17607 8139 17613 8159
rect 17527 8136 17613 8139
rect -251 8124 0 8128
rect -251 8104 -245 8124
rect -225 8104 -206 8124
rect -186 8104 -167 8124
rect -147 8104 -128 8124
rect -108 8104 0 8124
rect -251 8100 0 8104
rect 17068 8124 17313 8128
rect 17068 8104 17170 8124
rect 17190 8104 17209 8124
rect 17229 8104 17248 8124
rect 17268 8104 17287 8124
rect 17307 8104 17313 8124
rect 17068 8100 17313 8104
rect -2149 7968 -2143 7994
rect -1968 7968 -1962 7994
rect 17706 7968 17712 7994
rect 17887 7968 17893 7994
rect -440 7953 0 7957
rect -440 7933 -434 7953
rect -414 7933 -395 7953
rect -375 7933 -356 7953
rect -336 7933 -317 7953
rect -297 7933 0 7953
rect -440 7929 0 7933
rect 17068 7953 17503 7957
rect 17068 7933 17359 7953
rect 17379 7933 17398 7953
rect 17418 7933 17437 7953
rect 17457 7933 17476 7953
rect 17496 7933 17503 7953
rect 17068 7929 17503 7933
rect -659 7922 -625 7925
rect -659 7905 -651 7922
rect -634 7915 -625 7922
rect -634 7905 0 7915
rect -659 7901 0 7905
rect -1412 7803 -1389 7809
rect -1412 7786 -1409 7803
rect -1392 7800 -1389 7803
rect -1392 7786 0 7800
rect -1412 7780 -1389 7786
rect -800 7759 -777 7765
rect -800 7742 -797 7759
rect -780 7745 0 7759
rect -780 7742 -777 7745
rect -800 7736 -777 7742
rect -605 7728 0 7731
rect -605 7711 -597 7728
rect -580 7717 0 7728
rect -580 7711 -571 7717
rect -605 7707 -571 7711
rect -551 7657 -465 7660
rect -551 7637 -545 7657
rect -525 7637 -506 7657
rect -486 7654 -465 7657
rect 17527 7657 17613 7660
rect 17527 7654 17548 7657
rect -486 7640 0 7654
rect 17068 7640 17548 7654
rect -486 7637 -465 7640
rect -551 7634 -465 7637
rect 17527 7637 17548 7640
rect 17568 7637 17587 7657
rect 17607 7637 17613 7657
rect 17527 7634 17613 7637
rect -251 7622 0 7626
rect -251 7602 -245 7622
rect -225 7602 -206 7622
rect -186 7602 -167 7622
rect -147 7602 -128 7622
rect -108 7602 0 7622
rect -251 7598 0 7602
rect 17068 7622 17313 7626
rect 17068 7602 17170 7622
rect 17190 7602 17209 7622
rect 17229 7602 17248 7622
rect 17268 7602 17287 7622
rect 17307 7602 17313 7622
rect 17068 7598 17313 7602
rect -2149 7528 -2143 7554
rect -1968 7528 -1962 7554
rect 17706 7528 17712 7554
rect 17887 7528 17893 7554
rect -440 7451 0 7455
rect -440 7431 -434 7451
rect -414 7431 -395 7451
rect -375 7431 -356 7451
rect -336 7431 -317 7451
rect -297 7431 0 7451
rect -440 7427 0 7431
rect 17068 7451 17503 7455
rect 17068 7431 17359 7451
rect 17379 7431 17398 7451
rect 17418 7431 17437 7451
rect 17457 7431 17476 7451
rect 17496 7431 17503 7451
rect 17068 7427 17503 7431
rect -659 7420 -625 7423
rect -659 7403 -651 7420
rect -634 7413 -625 7420
rect -634 7403 0 7413
rect -659 7399 0 7403
rect -1448 7300 -1425 7306
rect -1448 7283 -1445 7300
rect -1428 7298 -1425 7300
rect -1428 7284 0 7298
rect -1428 7283 -1425 7284
rect -1448 7277 -1425 7283
rect -836 7259 -813 7265
rect -836 7242 -833 7259
rect -816 7257 -813 7259
rect -816 7243 0 7257
rect -816 7242 -813 7243
rect -836 7236 -813 7242
rect -605 7226 0 7229
rect -605 7209 -597 7226
rect -580 7215 0 7226
rect -580 7209 -571 7215
rect -605 7205 -571 7209
rect -551 7155 -465 7158
rect -551 7135 -545 7155
rect -525 7135 -506 7155
rect -486 7152 -465 7155
rect 17527 7155 17613 7158
rect 17527 7152 17548 7155
rect -486 7138 0 7152
rect 17068 7138 17548 7152
rect -486 7135 -465 7138
rect -551 7132 -465 7135
rect 17527 7135 17548 7138
rect 17568 7135 17587 7155
rect 17607 7135 17613 7155
rect 17527 7132 17613 7135
rect -251 7120 0 7124
rect -2149 7088 -2143 7114
rect -1968 7088 -1962 7114
rect -251 7100 -245 7120
rect -225 7100 -206 7120
rect -186 7100 -167 7120
rect -147 7100 -128 7120
rect -108 7100 0 7120
rect -251 7096 0 7100
rect 17068 7120 17313 7124
rect 17068 7100 17170 7120
rect 17190 7100 17209 7120
rect 17229 7100 17248 7120
rect 17268 7100 17287 7120
rect 17307 7100 17313 7120
rect 17068 7096 17313 7100
rect 17706 7088 17712 7114
rect 17887 7088 17893 7114
rect -440 6949 0 6953
rect -440 6929 -434 6949
rect -414 6929 -395 6949
rect -375 6929 -356 6949
rect -336 6929 -317 6949
rect -297 6929 0 6949
rect -440 6925 0 6929
rect 17068 6949 17503 6953
rect 17068 6929 17359 6949
rect 17379 6929 17398 6949
rect 17418 6929 17437 6949
rect 17457 6929 17476 6949
rect 17496 6929 17503 6949
rect 17068 6925 17503 6929
rect -659 6918 -625 6921
rect -659 6901 -651 6918
rect -634 6911 -625 6918
rect -634 6901 0 6911
rect -659 6897 0 6901
rect -1484 6797 -1461 6803
rect -1484 6780 -1481 6797
rect -1464 6796 -1461 6797
rect -1464 6782 0 6796
rect -1464 6780 -1461 6782
rect -1484 6774 -1461 6780
rect -872 6757 -849 6763
rect -872 6740 -869 6757
rect -852 6755 -849 6757
rect -852 6741 0 6755
rect -852 6740 -849 6741
rect -872 6734 -849 6740
rect -605 6724 0 6727
rect -605 6707 -597 6724
rect -580 6713 0 6724
rect -580 6707 -571 6713
rect -605 6703 -571 6707
rect -2149 6648 -2143 6674
rect -1968 6648 -1962 6674
rect -551 6653 -465 6656
rect -551 6633 -545 6653
rect -525 6633 -506 6653
rect -486 6650 -465 6653
rect 17527 6653 17613 6656
rect 17527 6650 17548 6653
rect -486 6636 0 6650
rect 17068 6636 17548 6650
rect -486 6633 -465 6636
rect -551 6630 -465 6633
rect 17527 6633 17548 6636
rect 17568 6633 17587 6653
rect 17607 6633 17613 6653
rect 17706 6648 17712 6674
rect 17887 6648 17893 6674
rect 17527 6630 17613 6633
rect -251 6618 0 6622
rect -251 6598 -245 6618
rect -225 6598 -206 6618
rect -186 6598 -167 6618
rect -147 6598 -128 6618
rect -108 6598 0 6618
rect -251 6594 0 6598
rect 17068 6618 17313 6622
rect 17068 6598 17170 6618
rect 17190 6598 17209 6618
rect 17229 6598 17248 6618
rect 17268 6598 17287 6618
rect 17307 6598 17313 6618
rect 17068 6594 17313 6598
rect -440 6447 0 6451
rect -440 6427 -434 6447
rect -414 6427 -395 6447
rect -375 6427 -356 6447
rect -336 6427 -317 6447
rect -297 6427 0 6447
rect -440 6423 0 6427
rect 17068 6447 17503 6451
rect 17068 6427 17359 6447
rect 17379 6427 17398 6447
rect 17418 6427 17437 6447
rect 17457 6427 17476 6447
rect 17496 6427 17503 6447
rect 17068 6423 17503 6427
rect -659 6416 -625 6419
rect -659 6399 -651 6416
rect -634 6409 -625 6416
rect -634 6399 0 6409
rect -659 6395 0 6399
rect -1520 6297 -1497 6303
rect -1520 6280 -1517 6297
rect -1500 6294 -1497 6297
rect -1500 6280 0 6294
rect -1520 6274 -1497 6280
rect -908 6256 -885 6262
rect -908 6239 -905 6256
rect -888 6253 -885 6256
rect -888 6239 0 6253
rect -2149 6208 -2143 6234
rect -1968 6208 -1962 6234
rect -908 6233 -885 6239
rect -605 6222 0 6225
rect -605 6205 -597 6222
rect -580 6211 0 6222
rect -580 6205 -571 6211
rect 17706 6208 17712 6234
rect 17887 6208 17893 6234
rect -605 6201 -571 6205
rect -551 6151 -465 6154
rect -551 6131 -545 6151
rect -525 6131 -506 6151
rect -486 6148 -465 6151
rect 17527 6151 17613 6154
rect 17527 6148 17548 6151
rect -486 6134 0 6148
rect 17068 6134 17548 6148
rect -486 6131 -465 6134
rect -551 6128 -465 6131
rect 17527 6131 17548 6134
rect 17568 6131 17587 6151
rect 17607 6131 17613 6151
rect 17527 6128 17613 6131
rect -251 6116 0 6120
rect -251 6096 -245 6116
rect -225 6096 -206 6116
rect -186 6096 -167 6116
rect -147 6096 -128 6116
rect -108 6096 0 6116
rect -251 6092 0 6096
rect 17068 6116 17313 6120
rect 17068 6096 17170 6116
rect 17190 6096 17209 6116
rect 17229 6096 17248 6116
rect 17268 6096 17287 6116
rect 17307 6096 17313 6116
rect 17068 6092 17313 6096
rect -440 5945 0 5949
rect -440 5925 -434 5945
rect -414 5925 -395 5945
rect -375 5925 -356 5945
rect -336 5925 -317 5945
rect -297 5925 0 5945
rect -440 5921 0 5925
rect 17068 5945 17503 5949
rect 17068 5925 17359 5945
rect 17379 5925 17398 5945
rect 17418 5925 17437 5945
rect 17457 5925 17476 5945
rect 17496 5925 17503 5945
rect 17068 5921 17503 5925
rect -659 5914 -625 5917
rect -659 5897 -651 5914
rect -634 5907 -625 5914
rect -634 5897 0 5907
rect -659 5893 0 5897
rect -1556 5795 -1533 5801
rect -2149 5768 -2143 5794
rect -1968 5768 -1962 5794
rect -1556 5778 -1553 5795
rect -1536 5792 -1533 5795
rect -1536 5778 0 5792
rect -1556 5772 -1533 5778
rect 17706 5768 17712 5794
rect 17887 5768 17893 5794
rect -944 5752 -921 5758
rect -944 5735 -941 5752
rect -924 5751 -921 5752
rect -924 5737 0 5751
rect -924 5735 -921 5737
rect -944 5729 -921 5735
rect -605 5720 0 5723
rect -605 5703 -597 5720
rect -580 5709 0 5720
rect -580 5703 -571 5709
rect -605 5699 -571 5703
rect -551 5649 -465 5652
rect -551 5629 -545 5649
rect -525 5629 -506 5649
rect -486 5646 -465 5649
rect 17527 5649 17613 5652
rect 17527 5646 17548 5649
rect -486 5632 0 5646
rect 17068 5632 17548 5646
rect -486 5629 -465 5632
rect -551 5626 -465 5629
rect 17527 5629 17548 5632
rect 17568 5629 17587 5649
rect 17607 5629 17613 5649
rect 17527 5626 17613 5629
rect -251 5614 0 5618
rect -251 5594 -245 5614
rect -225 5594 -206 5614
rect -186 5594 -167 5614
rect -147 5594 -128 5614
rect -108 5594 0 5614
rect -251 5590 0 5594
rect 17068 5614 17313 5618
rect 17068 5594 17170 5614
rect 17190 5594 17209 5614
rect 17229 5594 17248 5614
rect 17268 5594 17287 5614
rect 17307 5594 17313 5614
rect 17068 5590 17313 5594
rect -440 5443 0 5447
rect -440 5423 -434 5443
rect -414 5423 -395 5443
rect -375 5423 -356 5443
rect -336 5423 -317 5443
rect -297 5423 0 5443
rect -440 5419 0 5423
rect 17068 5443 17503 5447
rect 17068 5423 17359 5443
rect 17379 5423 17398 5443
rect 17418 5423 17437 5443
rect 17457 5423 17476 5443
rect 17496 5423 17503 5443
rect 17068 5419 17503 5423
rect -659 5412 -625 5415
rect -659 5395 -651 5412
rect -634 5405 -625 5412
rect -634 5395 0 5405
rect -659 5391 0 5395
rect -2149 5328 -2143 5354
rect -1968 5328 -1962 5354
rect 17706 5328 17712 5354
rect 17887 5328 17893 5354
rect -1592 5293 -1569 5299
rect -1592 5276 -1589 5293
rect -1572 5290 -1569 5293
rect -1572 5276 0 5290
rect -1592 5270 -1569 5276
rect -980 5252 -957 5258
rect -980 5235 -977 5252
rect -960 5249 -957 5252
rect -960 5235 0 5249
rect -980 5229 -957 5235
rect -605 5218 0 5221
rect -605 5201 -597 5218
rect -580 5207 0 5218
rect -580 5201 -571 5207
rect -605 5197 -571 5201
rect -551 5147 -465 5150
rect -551 5127 -545 5147
rect -525 5127 -506 5147
rect -486 5144 -465 5147
rect 17527 5147 17613 5150
rect 17527 5144 17548 5147
rect -486 5130 0 5144
rect 17068 5130 17548 5144
rect -486 5127 -465 5130
rect -551 5124 -465 5127
rect 17527 5127 17548 5130
rect 17568 5127 17587 5147
rect 17607 5127 17613 5147
rect 17527 5124 17613 5127
rect -251 5112 0 5116
rect -251 5092 -245 5112
rect -225 5092 -206 5112
rect -186 5092 -167 5112
rect -147 5092 -128 5112
rect -108 5092 0 5112
rect -251 5088 0 5092
rect 17068 5112 17313 5116
rect 17068 5092 17170 5112
rect 17190 5092 17209 5112
rect 17229 5092 17248 5112
rect 17268 5092 17287 5112
rect 17307 5092 17313 5112
rect 17068 5088 17313 5092
rect -440 4941 0 4945
rect -440 4921 -434 4941
rect -414 4921 -395 4941
rect -375 4921 -356 4941
rect -336 4921 -317 4941
rect -297 4921 0 4941
rect -440 4917 0 4921
rect 17068 4941 17503 4945
rect 17068 4921 17359 4941
rect 17379 4921 17398 4941
rect 17418 4921 17437 4941
rect 17457 4921 17476 4941
rect 17496 4921 17503 4941
rect 17068 4917 17503 4921
rect -2149 4888 -2143 4914
rect -1968 4888 -1962 4914
rect -659 4910 -625 4913
rect -659 4893 -651 4910
rect -634 4903 -625 4910
rect -634 4893 0 4903
rect -659 4889 0 4893
rect 17706 4888 17712 4914
rect 17887 4888 17893 4914
rect -1628 4790 -1605 4796
rect -1628 4773 -1625 4790
rect -1608 4788 -1605 4790
rect -1608 4774 0 4788
rect -1608 4773 -1605 4774
rect -1628 4767 -1605 4773
rect -1016 4749 -993 4755
rect -1016 4732 -1013 4749
rect -996 4747 -993 4749
rect -996 4733 0 4747
rect -996 4732 -993 4733
rect -1016 4726 -993 4732
rect -605 4716 0 4719
rect -605 4699 -597 4716
rect -580 4705 0 4716
rect -580 4699 -571 4705
rect -605 4695 -571 4699
rect -551 4645 -465 4648
rect -551 4625 -545 4645
rect -525 4625 -506 4645
rect -486 4642 -465 4645
rect 17527 4645 17613 4648
rect 17527 4642 17548 4645
rect -486 4628 0 4642
rect 17068 4628 17548 4642
rect -486 4625 -465 4628
rect -551 4622 -465 4625
rect 17527 4625 17548 4628
rect 17568 4625 17587 4645
rect 17607 4625 17613 4645
rect 17527 4622 17613 4625
rect -251 4610 0 4614
rect -251 4590 -245 4610
rect -225 4590 -206 4610
rect -186 4590 -167 4610
rect -147 4590 -128 4610
rect -108 4590 0 4610
rect -251 4586 0 4590
rect 17068 4610 17313 4614
rect 17068 4590 17170 4610
rect 17190 4590 17209 4610
rect 17229 4590 17248 4610
rect 17268 4590 17287 4610
rect 17307 4590 17313 4610
rect 17068 4586 17313 4590
rect -2149 4448 -2143 4474
rect -1968 4448 -1962 4474
rect 17706 4448 17712 4474
rect 17887 4448 17893 4474
rect -440 4439 0 4443
rect -440 4419 -434 4439
rect -414 4419 -395 4439
rect -375 4419 -356 4439
rect -336 4419 -317 4439
rect -297 4419 0 4439
rect -440 4415 0 4419
rect 17068 4439 17503 4443
rect 17068 4419 17359 4439
rect 17379 4419 17398 4439
rect 17418 4419 17437 4439
rect 17457 4419 17476 4439
rect 17496 4419 17503 4439
rect 17068 4415 17503 4419
rect -659 4408 -625 4411
rect -659 4391 -651 4408
rect -634 4401 -625 4408
rect -634 4391 0 4401
rect -659 4387 0 4391
rect -1664 4289 -1641 4295
rect -1664 4272 -1661 4289
rect -1644 4286 -1641 4289
rect -1644 4272 0 4286
rect -1664 4266 -1641 4272
rect -1052 4250 -1029 4256
rect -1052 4233 -1049 4250
rect -1032 4245 -1029 4250
rect -1032 4233 0 4245
rect -1052 4231 0 4233
rect -1052 4227 -1029 4231
rect -605 4214 0 4217
rect -605 4197 -597 4214
rect -580 4203 0 4214
rect -580 4197 -571 4203
rect -605 4193 -571 4197
rect -551 4143 -465 4146
rect -551 4123 -545 4143
rect -525 4123 -506 4143
rect -486 4140 -465 4143
rect 17527 4143 17613 4146
rect 17527 4140 17548 4143
rect -486 4126 0 4140
rect 17068 4126 17548 4140
rect -486 4123 -465 4126
rect -551 4120 -465 4123
rect 17527 4123 17548 4126
rect 17568 4123 17587 4143
rect 17607 4123 17613 4143
rect 17527 4120 17613 4123
rect -251 4108 0 4112
rect -251 4088 -245 4108
rect -225 4088 -206 4108
rect -186 4088 -167 4108
rect -147 4088 -128 4108
rect -108 4088 0 4108
rect -251 4084 0 4088
rect 17068 4108 17313 4112
rect 17068 4088 17170 4108
rect 17190 4088 17209 4108
rect 17229 4088 17248 4108
rect 17268 4088 17287 4108
rect 17307 4088 17313 4108
rect 17068 4084 17313 4088
rect -2149 4008 -2143 4034
rect -1968 4008 -1962 4034
rect 17706 4008 17712 4034
rect 17887 4008 17893 4034
rect -440 3937 0 3941
rect -440 3917 -434 3937
rect -414 3917 -395 3937
rect -375 3917 -356 3937
rect -336 3917 -317 3937
rect -297 3917 0 3937
rect -440 3913 0 3917
rect 17068 3937 17503 3941
rect 17068 3917 17359 3937
rect 17379 3917 17398 3937
rect 17418 3917 17437 3937
rect 17457 3917 17476 3937
rect 17496 3917 17503 3937
rect 17068 3913 17503 3917
rect -659 3906 -625 3909
rect -659 3889 -651 3906
rect -634 3899 -625 3906
rect -634 3889 0 3899
rect -659 3885 0 3889
rect -1700 3787 -1677 3793
rect -1700 3770 -1697 3787
rect -1680 3784 -1677 3787
rect -1680 3770 0 3784
rect -1700 3764 -1677 3770
rect -1088 3747 -1065 3753
rect -1088 3730 -1085 3747
rect -1068 3743 -1065 3747
rect -1068 3730 0 3743
rect -1088 3729 0 3730
rect -1088 3724 -1065 3729
rect -605 3712 0 3715
rect -605 3695 -597 3712
rect -580 3701 0 3712
rect -580 3695 -571 3701
rect -605 3691 -571 3695
rect -551 3641 -465 3644
rect -551 3621 -545 3641
rect -525 3621 -506 3641
rect -486 3638 -465 3641
rect 17527 3641 17613 3644
rect 17527 3638 17548 3641
rect -486 3624 0 3638
rect 17068 3624 17548 3638
rect -486 3621 -465 3624
rect -551 3618 -465 3621
rect 17527 3621 17548 3624
rect 17568 3621 17587 3641
rect 17607 3621 17613 3641
rect 17527 3618 17613 3621
rect -251 3606 0 3610
rect -2149 3568 -2143 3594
rect -1968 3568 -1962 3594
rect -251 3586 -245 3606
rect -225 3586 -206 3606
rect -186 3586 -167 3606
rect -147 3586 -128 3606
rect -108 3586 0 3606
rect -251 3582 0 3586
rect 17068 3606 17313 3610
rect 17068 3586 17170 3606
rect 17190 3586 17209 3606
rect 17229 3586 17248 3606
rect 17268 3586 17287 3606
rect 17307 3586 17313 3606
rect 17068 3582 17313 3586
rect 17706 3568 17712 3594
rect 17887 3568 17893 3594
rect -440 3435 0 3439
rect -440 3415 -434 3435
rect -414 3415 -395 3435
rect -375 3415 -356 3435
rect -336 3415 -317 3435
rect -297 3415 0 3435
rect -440 3411 0 3415
rect 17068 3435 17503 3439
rect 17068 3415 17359 3435
rect 17379 3415 17398 3435
rect 17418 3415 17437 3435
rect 17457 3415 17476 3435
rect 17496 3415 17503 3435
rect 17068 3411 17503 3415
rect -659 3404 -625 3407
rect -659 3387 -651 3404
rect -634 3397 -625 3404
rect -634 3387 0 3397
rect -659 3383 0 3387
rect -1736 3285 -1713 3291
rect -1736 3268 -1733 3285
rect -1716 3282 -1713 3285
rect -1716 3268 0 3282
rect -1736 3262 -1713 3268
rect -1124 3245 -1101 3251
rect -1124 3228 -1121 3245
rect -1104 3241 -1101 3245
rect -1104 3228 0 3241
rect -1124 3227 0 3228
rect -1124 3222 -1101 3227
rect -605 3210 0 3213
rect -605 3193 -597 3210
rect -580 3199 0 3210
rect -580 3193 -571 3199
rect -605 3189 -571 3193
rect -2149 3128 -2143 3154
rect -1968 3128 -1962 3154
rect -551 3139 -465 3142
rect -551 3119 -545 3139
rect -525 3119 -506 3139
rect -486 3136 -465 3139
rect 17527 3139 17613 3142
rect 17527 3136 17548 3139
rect -486 3122 0 3136
rect 17068 3122 17548 3136
rect -486 3119 -465 3122
rect -551 3116 -465 3119
rect 17527 3119 17548 3122
rect 17568 3119 17587 3139
rect 17607 3119 17613 3139
rect 17706 3128 17712 3154
rect 17887 3128 17893 3154
rect 17527 3116 17613 3119
rect -251 3104 0 3108
rect -251 3084 -245 3104
rect -225 3084 -206 3104
rect -186 3084 -167 3104
rect -147 3084 -128 3104
rect -108 3084 0 3104
rect -251 3080 0 3084
rect 17068 3104 17313 3108
rect 17068 3084 17170 3104
rect 17190 3084 17209 3104
rect 17229 3084 17248 3104
rect 17268 3084 17287 3104
rect 17307 3084 17313 3104
rect 17068 3080 17313 3084
rect -440 2933 0 2937
rect -440 2913 -434 2933
rect -414 2913 -395 2933
rect -375 2913 -356 2933
rect -336 2913 -317 2933
rect -297 2913 0 2933
rect -440 2909 0 2913
rect 17068 2933 17503 2937
rect 17068 2913 17359 2933
rect 17379 2913 17398 2933
rect 17418 2913 17437 2933
rect 17457 2913 17476 2933
rect 17496 2913 17503 2933
rect 17068 2909 17503 2913
rect -659 2902 -625 2905
rect -659 2885 -651 2902
rect -634 2895 -625 2902
rect -634 2885 0 2895
rect -659 2881 0 2885
rect -1772 2783 -1749 2789
rect -1772 2766 -1769 2783
rect -1752 2780 -1749 2783
rect -1752 2766 0 2780
rect -1772 2760 -1749 2766
rect -1160 2744 -1137 2750
rect -1160 2727 -1157 2744
rect -1140 2739 -1137 2744
rect -1140 2727 0 2739
rect -1160 2725 0 2727
rect -1160 2721 -1137 2725
rect -2149 2688 -2143 2714
rect -1968 2688 -1962 2714
rect -605 2708 0 2711
rect -605 2691 -597 2708
rect -580 2697 0 2708
rect -580 2691 -571 2697
rect -605 2687 -571 2691
rect 17706 2688 17712 2714
rect 17887 2688 17893 2714
rect -551 2637 -465 2640
rect -551 2617 -545 2637
rect -525 2617 -506 2637
rect -486 2634 -465 2637
rect 17527 2637 17613 2640
rect 17527 2634 17548 2637
rect -486 2620 0 2634
rect 17068 2620 17548 2634
rect -486 2617 -465 2620
rect -551 2614 -465 2617
rect 17527 2617 17548 2620
rect 17568 2617 17587 2637
rect 17607 2617 17613 2637
rect 17527 2614 17613 2617
rect -251 2602 0 2606
rect -251 2582 -245 2602
rect -225 2582 -206 2602
rect -186 2582 -167 2602
rect -147 2582 -128 2602
rect -108 2582 0 2602
rect -251 2578 0 2582
rect 17068 2602 17313 2606
rect 17068 2582 17170 2602
rect 17190 2582 17209 2602
rect 17229 2582 17248 2602
rect 17268 2582 17287 2602
rect 17307 2582 17313 2602
rect 17068 2578 17313 2582
rect -440 2431 0 2435
rect -440 2411 -434 2431
rect -414 2411 -395 2431
rect -375 2411 -356 2431
rect -336 2411 -317 2431
rect -297 2411 0 2431
rect -440 2407 0 2411
rect 17068 2431 17503 2435
rect 17068 2411 17359 2431
rect 17379 2411 17398 2431
rect 17418 2411 17437 2431
rect 17457 2411 17476 2431
rect 17496 2411 17503 2431
rect 17068 2407 17503 2411
rect -659 2400 -625 2403
rect -659 2383 -651 2400
rect -634 2393 -625 2400
rect -634 2383 0 2393
rect -659 2379 0 2383
rect -1808 2282 -1785 2288
rect -2149 2248 -2143 2274
rect -1968 2248 -1962 2274
rect -1808 2265 -1805 2282
rect -1788 2278 -1785 2282
rect -1788 2265 0 2278
rect -1808 2264 0 2265
rect -1808 2259 -1785 2264
rect 17706 2248 17712 2274
rect 17887 2248 17893 2274
rect -1196 2239 -1173 2245
rect -1196 2222 -1193 2239
rect -1176 2237 -1173 2239
rect -1176 2223 0 2237
rect -1176 2222 -1173 2223
rect -1196 2216 -1173 2222
rect -605 2206 0 2209
rect -605 2189 -597 2206
rect -580 2195 0 2206
rect -580 2189 -571 2195
rect -605 2185 -571 2189
rect -551 2135 -465 2138
rect -551 2115 -545 2135
rect -525 2115 -506 2135
rect -486 2132 -465 2135
rect 17527 2135 17613 2138
rect 17527 2132 17548 2135
rect -486 2118 0 2132
rect 17068 2118 17548 2132
rect -486 2115 -465 2118
rect -551 2112 -465 2115
rect 17527 2115 17548 2118
rect 17568 2115 17587 2135
rect 17607 2115 17613 2135
rect 17527 2112 17613 2115
rect -251 2100 0 2104
rect -251 2080 -245 2100
rect -225 2080 -206 2100
rect -186 2080 -167 2100
rect -147 2080 -128 2100
rect -108 2080 0 2100
rect -251 2076 0 2080
rect 17068 2100 17313 2104
rect 17068 2080 17170 2100
rect 17190 2080 17209 2100
rect 17229 2080 17248 2100
rect 17268 2080 17287 2100
rect 17307 2080 17313 2100
rect 17068 2076 17313 2080
rect -440 1929 0 1933
rect -440 1909 -434 1929
rect -414 1909 -395 1929
rect -375 1909 -356 1929
rect -336 1909 -317 1929
rect -297 1909 0 1929
rect -440 1905 0 1909
rect 17068 1929 17503 1933
rect 17068 1909 17359 1929
rect 17379 1909 17398 1929
rect 17418 1909 17437 1929
rect 17457 1909 17476 1929
rect 17496 1909 17503 1929
rect 17068 1905 17503 1909
rect -659 1898 -625 1901
rect -659 1881 -651 1898
rect -634 1891 -625 1898
rect -634 1881 0 1891
rect -659 1877 0 1881
rect -2149 1808 -2143 1834
rect -1968 1808 -1962 1834
rect 17706 1808 17712 1834
rect 17887 1808 17893 1834
rect -1844 1779 -1821 1785
rect -1844 1762 -1841 1779
rect -1824 1776 -1821 1779
rect -1824 1762 0 1776
rect -1844 1756 -1821 1762
rect -1232 1736 -1209 1742
rect -1232 1719 -1229 1736
rect -1212 1735 -1209 1736
rect -1212 1721 0 1735
rect -1212 1719 -1209 1721
rect -1232 1713 -1209 1719
rect -605 1704 0 1707
rect -605 1687 -597 1704
rect -580 1693 0 1704
rect -580 1687 -571 1693
rect -605 1683 -571 1687
rect -551 1633 -465 1636
rect -551 1613 -545 1633
rect -525 1613 -506 1633
rect -486 1630 -465 1633
rect 17527 1633 17613 1636
rect 17527 1630 17548 1633
rect -486 1616 0 1630
rect 17068 1616 17548 1630
rect -486 1613 -465 1616
rect -551 1610 -465 1613
rect 17527 1613 17548 1616
rect 17568 1613 17587 1633
rect 17607 1613 17613 1633
rect 17527 1610 17613 1613
rect -251 1598 0 1602
rect -251 1578 -245 1598
rect -225 1578 -206 1598
rect -186 1578 -167 1598
rect -147 1578 -128 1598
rect -108 1578 0 1598
rect -251 1574 0 1578
rect 17068 1598 17313 1602
rect 17068 1578 17170 1598
rect 17190 1578 17209 1598
rect 17229 1578 17248 1598
rect 17268 1578 17287 1598
rect 17307 1578 17313 1598
rect 17068 1574 17313 1578
rect -440 1427 0 1431
rect -440 1407 -434 1427
rect -414 1407 -395 1427
rect -375 1407 -356 1427
rect -336 1407 -317 1427
rect -297 1407 0 1427
rect -440 1403 0 1407
rect 17068 1427 17503 1431
rect 17068 1407 17359 1427
rect 17379 1407 17398 1427
rect 17418 1407 17437 1427
rect 17457 1407 17476 1427
rect 17496 1407 17503 1427
rect 17068 1403 17503 1407
rect -659 1396 -625 1399
rect -2149 1368 -2143 1394
rect -1968 1368 -1962 1394
rect -659 1379 -651 1396
rect -634 1389 -625 1396
rect -634 1379 0 1389
rect -659 1375 0 1379
rect 17706 1368 17712 1394
rect 17887 1368 17893 1394
rect -1880 1276 -1857 1282
rect -1880 1259 -1877 1276
rect -1860 1274 -1857 1276
rect -1860 1260 0 1274
rect -1860 1259 -1857 1260
rect -1880 1253 -1857 1259
rect -1268 1233 -1245 1239
rect -1268 1216 -1265 1233
rect -1248 1219 0 1233
rect -1248 1216 -1245 1219
rect -1268 1210 -1245 1216
rect -605 1202 0 1205
rect -605 1185 -597 1202
rect -580 1191 0 1202
rect -580 1185 -571 1191
rect -605 1181 -571 1185
rect -551 1131 -465 1134
rect -551 1111 -545 1131
rect -525 1111 -506 1131
rect -486 1128 -465 1131
rect 17527 1131 17613 1134
rect 17527 1128 17548 1131
rect -486 1114 0 1128
rect 17068 1114 17548 1128
rect -486 1111 -465 1114
rect -551 1108 -465 1111
rect 17527 1111 17548 1114
rect 17568 1111 17587 1131
rect 17607 1111 17613 1131
rect 17527 1108 17613 1111
rect -251 1096 0 1100
rect -251 1076 -245 1096
rect -225 1076 -206 1096
rect -186 1076 -167 1096
rect -147 1076 -128 1096
rect -108 1076 0 1096
rect -251 1072 0 1076
rect 17068 1096 17313 1100
rect 17068 1076 17170 1096
rect 17190 1076 17209 1096
rect 17229 1076 17248 1096
rect 17268 1076 17287 1096
rect 17307 1076 17313 1096
rect 17068 1072 17313 1076
rect -2149 928 -2143 954
rect -1968 928 -1962 954
rect -440 925 0 929
rect -440 905 -434 925
rect -414 905 -395 925
rect -375 905 -356 925
rect -336 905 -317 925
rect -297 905 0 925
rect -440 901 0 905
rect 17068 925 17503 929
rect 17706 928 17712 954
rect 17887 928 17893 954
rect 17068 905 17359 925
rect 17379 905 17398 925
rect 17418 905 17437 925
rect 17457 905 17476 925
rect 17496 905 17503 925
rect 17068 901 17503 905
rect -659 894 -625 897
rect -659 877 -651 894
rect -634 887 -625 894
rect -634 877 0 887
rect -659 873 0 877
rect -1916 775 -1893 781
rect -1916 758 -1913 775
rect -1896 772 -1893 775
rect -1896 758 0 772
rect -1916 752 -1893 758
rect -1304 735 -1281 741
rect -1304 718 -1301 735
rect -1284 731 -1281 735
rect -1284 718 0 731
rect -1304 717 0 718
rect -1304 712 -1281 717
rect -605 700 0 703
rect -605 683 -597 700
rect -580 689 0 700
rect -580 683 -571 689
rect -605 679 -571 683
rect -551 629 -465 632
rect -551 609 -545 629
rect -525 609 -506 629
rect -486 626 -465 629
rect 17527 629 17613 632
rect 17527 626 17548 629
rect -486 612 0 626
rect 17068 612 17548 626
rect -486 609 -465 612
rect -551 606 -465 609
rect 17527 609 17548 612
rect 17568 609 17587 629
rect 17607 609 17613 629
rect 17527 606 17613 609
rect -251 594 0 598
rect -251 574 -245 594
rect -225 574 -206 594
rect -186 574 -167 594
rect -147 574 -128 594
rect -108 574 0 594
rect -251 570 0 574
rect 17068 594 17313 598
rect 17068 574 17170 594
rect 17190 574 17209 594
rect 17229 574 17248 594
rect 17268 574 17287 594
rect 17307 574 17313 594
rect 17068 570 17313 574
rect -2149 488 -2143 514
rect -1968 488 -1962 514
rect 17706 488 17712 514
rect 17887 488 17893 514
rect -440 423 0 427
rect -440 403 -434 423
rect -414 403 -395 423
rect -375 403 -356 423
rect -336 403 -317 423
rect -297 403 0 423
rect -440 399 0 403
rect 17068 423 17503 427
rect 17068 403 17359 423
rect 17379 403 17398 423
rect 17418 403 17437 423
rect 17457 403 17476 423
rect 17496 403 17503 423
rect 17068 399 17503 403
rect -440 381 0 385
rect -440 361 -434 381
rect -414 361 -395 381
rect -375 361 -356 381
rect -336 361 -317 381
rect -297 371 0 381
rect -297 361 -291 371
rect -440 357 -291 361
rect -251 256 0 270
rect -251 253 -102 256
rect -251 233 -245 253
rect -225 233 -206 253
rect -186 233 -167 253
rect -147 233 -128 253
rect -108 233 -102 253
rect -251 229 -102 233
rect -251 215 0 229
rect -251 197 0 201
rect -251 177 -245 197
rect -225 177 -206 197
rect -186 177 -167 197
rect -147 177 -128 197
rect -108 187 0 197
rect -108 177 -102 187
rect -251 173 -102 177
rect -551 127 -465 130
rect -551 107 -545 127
rect -525 107 -506 127
rect -486 124 -465 127
rect 17527 127 17613 130
rect 17527 124 17548 127
rect -486 110 0 124
rect 17068 110 17548 124
rect -486 107 -465 110
rect -551 104 -465 107
rect 17527 107 17548 110
rect 17568 107 17587 127
rect 17607 107 17613 127
rect 17527 104 17613 107
rect -251 92 0 96
rect -2149 48 -2143 74
rect -1968 48 -1962 74
rect -251 72 -245 92
rect -225 72 -206 92
rect -186 72 -167 92
rect -147 72 -128 92
rect -108 72 0 92
rect -251 68 0 72
rect 17068 92 17313 96
rect 17068 72 17170 92
rect 17190 72 17209 92
rect 17229 72 17248 92
rect 17268 72 17287 92
rect 17307 72 17313 92
rect 17068 68 17313 72
rect 17706 48 17712 74
rect 17887 48 17893 74
rect 17146 -13 17900 -12
rect 17146 -20 17901 -13
rect 17146 -48 17181 -20
rect 17209 -48 17228 -20
rect 17256 -48 17275 -20
rect 17303 -26 17901 -20
rect 17303 -48 17722 -26
rect 17146 -58 17722 -48
rect 17754 -58 17766 -26
rect 17798 -58 17810 -26
rect 17842 -58 17854 -26
rect 17886 -58 17901 -26
rect 16098 -64 16371 -61
rect -2156 -78 -1950 -77
rect -2157 -91 -1950 -78
rect -2157 -123 -2142 -91
rect -2110 -123 -2098 -91
rect -2066 -123 -2054 -91
rect -2022 -123 -2010 -91
rect -1978 -123 -1950 -91
rect -2157 -136 -1950 -123
rect -2157 -168 -2142 -136
rect -2110 -168 -2098 -136
rect -2066 -168 -2054 -136
rect -2022 -168 -2010 -136
rect -1978 -168 -1950 -136
rect -2157 -181 -1950 -168
rect -2157 -213 -2142 -181
rect -2110 -213 -2098 -181
rect -2066 -213 -2054 -181
rect -2022 -213 -2010 -181
rect -1978 -213 -1950 -181
rect -2157 -217 -1950 -213
rect -273 -85 -91 -77
rect 16098 -81 16104 -64
rect 16121 -81 16348 -64
rect 16365 -81 16371 -64
rect 16098 -85 16371 -81
rect 17146 -67 17901 -58
rect -273 -113 -241 -85
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -91 -85
rect -273 -132 -91 -113
rect -273 -160 -241 -132
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -91 -132
rect 17146 -95 17181 -67
rect 17209 -95 17228 -67
rect 17256 -95 17275 -67
rect 17303 -71 17901 -67
rect 17303 -95 17722 -71
rect 17146 -103 17722 -95
rect 17754 -103 17766 -71
rect 17798 -103 17810 -71
rect 17842 -103 17854 -71
rect 17886 -103 17901 -71
rect 17146 -114 17901 -103
rect 13277 -136 14506 -133
rect 13277 -153 13283 -136
rect 13300 -153 14483 -136
rect 14500 -153 14506 -136
rect 17146 -142 17181 -114
rect 17209 -142 17228 -114
rect 17256 -142 17275 -114
rect 17303 -116 17901 -114
rect 17303 -142 17722 -116
rect 17146 -148 17722 -142
rect 17754 -148 17766 -116
rect 17798 -148 17810 -116
rect 17842 -148 17854 -116
rect 17886 -148 17901 -116
rect 17146 -152 17901 -148
rect 13277 -157 14506 -153
rect -273 -179 -91 -160
rect -273 -207 -241 -179
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -91 -179
rect 13379 -175 15008 -172
rect 13379 -192 13385 -175
rect 13402 -192 14985 -175
rect 15002 -192 15008 -175
rect 13379 -196 15008 -192
rect -273 -217 -91 -207
rect 13481 -213 15510 -210
rect 13481 -230 13487 -213
rect 13504 -230 15487 -213
rect 15504 -230 15510 -213
rect 13481 -234 15510 -230
rect 17146 -231 17503 -230
rect 17146 -238 18196 -231
rect 13583 -251 16012 -248
rect 13583 -268 13589 -251
rect 13606 -268 15989 -251
rect 16006 -268 16012 -251
rect 13583 -272 16012 -268
rect 17146 -266 17370 -238
rect 17398 -266 17417 -238
rect 17445 -266 17464 -238
rect 17492 -245 18196 -238
rect 17492 -266 18017 -245
rect 17146 -277 18017 -266
rect 18049 -277 18061 -245
rect 18093 -277 18105 -245
rect 18137 -277 18149 -245
rect 18181 -277 18196 -245
rect 17146 -285 18196 -277
rect 13685 -289 16514 -286
rect 422 -295 448 -292
rect -385 -296 425 -295
rect -2452 -310 -2245 -296
rect -2452 -342 -2437 -310
rect -2405 -342 -2393 -310
rect -2361 -342 -2349 -310
rect -2317 -342 -2305 -310
rect -2273 -342 -2245 -310
rect -2452 -355 -2245 -342
rect -2452 -387 -2437 -355
rect -2405 -387 -2393 -355
rect -2361 -387 -2349 -355
rect -2317 -387 -2305 -355
rect -2273 -387 -2245 -355
rect -2452 -400 -2245 -387
rect -2452 -432 -2437 -400
rect -2405 -432 -2393 -400
rect -2361 -432 -2349 -400
rect -2317 -432 -2305 -400
rect -2273 -432 -2245 -400
rect -2452 -436 -2245 -432
rect -462 -304 425 -296
rect -462 -332 -430 -304
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -312 425 -304
rect 442 -312 448 -295
rect 13685 -306 13691 -289
rect 13708 -306 16491 -289
rect 16508 -306 16514 -289
rect 17146 -295 17370 -285
rect 13685 -310 16514 -306
rect 16989 -298 17370 -295
rect -308 -316 448 -312
rect 16989 -315 16995 -298
rect 17012 -313 17370 -298
rect 17398 -313 17417 -285
rect 17445 -313 17464 -285
rect 17492 -290 18196 -285
rect 17492 -313 18017 -290
rect 17012 -315 18017 -313
rect -308 -332 -91 -316
rect 16989 -319 18017 -315
rect -462 -351 -91 -332
rect -462 -379 -430 -351
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -91 -351
rect 17146 -322 18017 -319
rect 18049 -322 18061 -290
rect 18093 -322 18105 -290
rect 18137 -322 18149 -290
rect 18181 -322 18196 -290
rect 17146 -332 18196 -322
rect 17146 -360 17370 -332
rect 17398 -360 17417 -332
rect 17445 -360 17464 -332
rect 17492 -335 18196 -332
rect 17492 -360 18017 -335
rect 17146 -367 18017 -360
rect 18049 -367 18061 -335
rect 18093 -367 18105 -335
rect 18137 -367 18149 -335
rect 18181 -367 18196 -335
rect 17146 -370 18196 -367
rect 17694 -371 18196 -370
rect -462 -398 -91 -379
rect -462 -426 -430 -398
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -91 -398
rect -462 -435 -91 -426
rect 16395 -432 18196 -429
rect -462 -436 -280 -435
rect 16395 -449 16401 -432
rect 16418 -449 16437 -432
rect 16454 -449 18196 -432
rect 16395 -453 18196 -449
<< via1 >>
rect -2437 9457 -2405 9489
rect -2393 9457 -2361 9489
rect -2349 9457 -2317 9489
rect -2305 9457 -2273 9489
rect 18017 9457 18049 9489
rect 18061 9457 18093 9489
rect 18105 9457 18137 9489
rect 18149 9457 18181 9489
rect -2437 9412 -2405 9444
rect -2393 9412 -2361 9444
rect -2349 9412 -2317 9444
rect -2305 9412 -2273 9444
rect 18017 9412 18049 9444
rect 18061 9412 18093 9444
rect 18105 9412 18137 9444
rect 18149 9412 18181 9444
rect -2437 9367 -2405 9399
rect -2393 9367 -2361 9399
rect -2349 9367 -2317 9399
rect -2305 9367 -2273 9399
rect 18017 9367 18049 9399
rect 18061 9367 18093 9399
rect 18105 9367 18137 9399
rect 18149 9367 18181 9399
rect -2142 9238 -2110 9270
rect -2098 9238 -2066 9270
rect -2054 9238 -2022 9270
rect -2010 9238 -1978 9270
rect 17722 9238 17754 9270
rect 17766 9238 17798 9270
rect 17810 9238 17842 9270
rect 17854 9238 17886 9270
rect -2142 9193 -2110 9225
rect -2098 9193 -2066 9225
rect -2054 9193 -2022 9225
rect -2010 9193 -1978 9225
rect 17722 9193 17754 9225
rect 17766 9193 17798 9225
rect 17810 9193 17842 9225
rect 17854 9193 17886 9225
rect -2142 9148 -2110 9180
rect -2098 9148 -2066 9180
rect -2054 9148 -2022 9180
rect -2010 9148 -1978 9180
rect 17722 9148 17754 9180
rect 17766 9148 17798 9180
rect 17810 9148 17842 9180
rect 17854 9148 17886 9180
rect -2143 8870 -1968 8874
rect -2143 8853 -1968 8870
rect -2143 8848 -1968 8853
rect 17712 8870 17887 8874
rect 17712 8853 17887 8870
rect 17712 8848 17887 8853
rect -2143 8430 -1968 8434
rect -2143 8413 -1968 8430
rect -2143 8408 -1968 8413
rect 17712 8430 17887 8434
rect 17712 8413 17887 8430
rect 17712 8408 17887 8413
rect -2143 7990 -1968 7994
rect -2143 7973 -1968 7990
rect -2143 7968 -1968 7973
rect 17712 7990 17887 7994
rect 17712 7973 17887 7990
rect 17712 7968 17887 7973
rect -2143 7550 -1968 7554
rect -2143 7533 -1968 7550
rect -2143 7528 -1968 7533
rect 17712 7550 17887 7554
rect 17712 7533 17887 7550
rect 17712 7528 17887 7533
rect -2143 7110 -1968 7114
rect -2143 7093 -1968 7110
rect -2143 7088 -1968 7093
rect 17712 7110 17887 7114
rect 17712 7093 17887 7110
rect 17712 7088 17887 7093
rect -2143 6670 -1968 6674
rect -2143 6653 -1968 6670
rect -2143 6648 -1968 6653
rect 17712 6670 17887 6674
rect 17712 6653 17887 6670
rect 17712 6648 17887 6653
rect -2143 6230 -1968 6234
rect -2143 6213 -1968 6230
rect -2143 6208 -1968 6213
rect 17712 6230 17887 6234
rect 17712 6213 17887 6230
rect 17712 6208 17887 6213
rect -2143 5790 -1968 5794
rect -2143 5773 -1968 5790
rect -2143 5768 -1968 5773
rect 17712 5790 17887 5794
rect 17712 5773 17887 5790
rect 17712 5768 17887 5773
rect -2143 5350 -1968 5354
rect -2143 5333 -1968 5350
rect -2143 5328 -1968 5333
rect 17712 5350 17887 5354
rect 17712 5333 17887 5350
rect 17712 5328 17887 5333
rect -2143 4910 -1968 4914
rect -2143 4893 -1968 4910
rect -2143 4888 -1968 4893
rect 17712 4910 17887 4914
rect 17712 4893 17887 4910
rect 17712 4888 17887 4893
rect -2143 4470 -1968 4474
rect -2143 4453 -1968 4470
rect -2143 4448 -1968 4453
rect 17712 4470 17887 4474
rect 17712 4453 17887 4470
rect 17712 4448 17887 4453
rect -2143 4030 -1968 4034
rect -2143 4013 -1968 4030
rect -2143 4008 -1968 4013
rect 17712 4030 17887 4034
rect 17712 4013 17887 4030
rect 17712 4008 17887 4013
rect -2143 3590 -1968 3594
rect -2143 3573 -1968 3590
rect -2143 3568 -1968 3573
rect 17712 3590 17887 3594
rect 17712 3573 17887 3590
rect 17712 3568 17887 3573
rect -2143 3150 -1968 3154
rect -2143 3133 -1968 3150
rect -2143 3128 -1968 3133
rect 17712 3150 17887 3154
rect 17712 3133 17887 3150
rect 17712 3128 17887 3133
rect -2143 2710 -1968 2714
rect -2143 2693 -1968 2710
rect -2143 2688 -1968 2693
rect 17712 2710 17887 2714
rect 17712 2693 17887 2710
rect 17712 2688 17887 2693
rect -2143 2270 -1968 2274
rect -2143 2253 -1968 2270
rect -2143 2248 -1968 2253
rect 17712 2270 17887 2274
rect 17712 2253 17887 2270
rect 17712 2248 17887 2253
rect -2143 1830 -1968 1834
rect -2143 1813 -1968 1830
rect -2143 1808 -1968 1813
rect 17712 1830 17887 1834
rect 17712 1813 17887 1830
rect 17712 1808 17887 1813
rect -2143 1390 -1968 1394
rect -2143 1373 -1968 1390
rect -2143 1368 -1968 1373
rect 17712 1390 17887 1394
rect 17712 1373 17887 1390
rect 17712 1368 17887 1373
rect -2143 950 -1968 954
rect -2143 933 -1968 950
rect -2143 928 -1968 933
rect 17712 950 17887 954
rect 17712 933 17887 950
rect 17712 928 17887 933
rect -2143 510 -1968 514
rect -2143 493 -1968 510
rect -2143 488 -1968 493
rect 17712 510 17887 514
rect 17712 493 17887 510
rect 17712 488 17887 493
rect -2143 70 -1968 74
rect -2143 53 -1968 70
rect -2143 48 -1968 53
rect 17712 70 17887 74
rect 17712 53 17887 70
rect 17712 48 17887 53
rect 17722 -58 17754 -26
rect 17766 -58 17798 -26
rect 17810 -58 17842 -26
rect 17854 -58 17886 -26
rect -2142 -123 -2110 -91
rect -2098 -123 -2066 -91
rect -2054 -123 -2022 -91
rect -2010 -123 -1978 -91
rect -2142 -168 -2110 -136
rect -2098 -168 -2066 -136
rect -2054 -168 -2022 -136
rect -2010 -168 -1978 -136
rect -2142 -213 -2110 -181
rect -2098 -213 -2066 -181
rect -2054 -213 -2022 -181
rect -2010 -213 -1978 -181
rect -241 -113 -213 -85
rect -194 -113 -166 -85
rect -147 -113 -119 -85
rect -241 -160 -213 -132
rect -194 -160 -166 -132
rect -147 -160 -119 -132
rect 17722 -103 17754 -71
rect 17766 -103 17798 -71
rect 17810 -103 17842 -71
rect 17854 -103 17886 -71
rect 17722 -148 17754 -116
rect 17766 -148 17798 -116
rect 17810 -148 17842 -116
rect 17854 -148 17886 -116
rect -241 -207 -213 -179
rect -194 -207 -166 -179
rect -147 -207 -119 -179
rect 18017 -277 18049 -245
rect 18061 -277 18093 -245
rect 18105 -277 18137 -245
rect 18149 -277 18181 -245
rect -2437 -342 -2405 -310
rect -2393 -342 -2361 -310
rect -2349 -342 -2317 -310
rect -2305 -342 -2273 -310
rect -2437 -387 -2405 -355
rect -2393 -387 -2361 -355
rect -2349 -387 -2317 -355
rect -2305 -387 -2273 -355
rect -2437 -432 -2405 -400
rect -2393 -432 -2361 -400
rect -2349 -432 -2317 -400
rect -2305 -432 -2273 -400
rect -430 -332 -402 -304
rect -383 -332 -355 -304
rect -336 -332 -308 -304
rect -430 -379 -402 -351
rect -383 -379 -355 -351
rect -336 -379 -308 -351
rect 18017 -322 18049 -290
rect 18061 -322 18093 -290
rect 18105 -322 18137 -290
rect 18149 -322 18181 -290
rect 18017 -367 18049 -335
rect 18061 -367 18093 -335
rect 18105 -367 18137 -335
rect 18149 -367 18181 -335
rect -430 -426 -402 -398
rect -383 -426 -355 -398
rect -336 -426 -308 -398
<< metal2 >>
rect -2452 9489 -2245 9493
rect -2452 9457 -2437 9489
rect -2405 9457 -2393 9489
rect -2361 9457 -2349 9489
rect -2317 9457 -2305 9489
rect -2273 9457 -2245 9489
rect -2452 9444 -2245 9457
rect -2452 9412 -2437 9444
rect -2405 9412 -2393 9444
rect -2361 9412 -2349 9444
rect -2317 9412 -2305 9444
rect -2273 9412 -2245 9444
rect -2452 9399 -2245 9412
rect -2452 9367 -2437 9399
rect -2405 9367 -2393 9399
rect -2361 9367 -2349 9399
rect -2317 9367 -2305 9399
rect -2273 9367 -2245 9399
rect -2452 9353 -2245 9367
rect 17989 9489 18196 9493
rect 17989 9457 18017 9489
rect 18049 9457 18061 9489
rect 18093 9457 18105 9489
rect 18137 9457 18149 9489
rect 18181 9457 18196 9489
rect 17989 9444 18196 9457
rect 17989 9412 18017 9444
rect 18049 9412 18061 9444
rect 18093 9412 18105 9444
rect 18137 9412 18149 9444
rect 18181 9412 18196 9444
rect 17989 9399 18196 9412
rect 17989 9367 18017 9399
rect 18049 9367 18061 9399
rect 18093 9367 18105 9399
rect 18137 9367 18149 9399
rect 18181 9367 18196 9399
rect 17989 9353 18196 9367
rect -2157 9270 -1950 9274
rect -2157 9238 -2142 9270
rect -2110 9238 -2098 9270
rect -2066 9238 -2054 9270
rect -2022 9238 -2010 9270
rect -1978 9238 -1950 9270
rect -2157 9225 -1950 9238
rect -2157 9193 -2142 9225
rect -2110 9193 -2098 9225
rect -2066 9193 -2054 9225
rect -2022 9193 -2010 9225
rect -1978 9193 -1950 9225
rect -2157 9180 -1950 9193
rect -2157 9148 -2142 9180
rect -2110 9148 -2098 9180
rect -2066 9148 -2054 9180
rect -2022 9148 -2010 9180
rect -1978 9148 -1950 9180
rect -2157 9134 -1950 9148
rect 17694 9270 17901 9274
rect 17694 9238 17722 9270
rect 17754 9238 17766 9270
rect 17798 9238 17810 9270
rect 17842 9238 17854 9270
rect 17886 9238 17901 9270
rect 17694 9225 17901 9238
rect 17694 9193 17722 9225
rect 17754 9193 17766 9225
rect 17798 9193 17810 9225
rect 17842 9193 17854 9225
rect 17886 9193 17901 9225
rect 17694 9180 17901 9193
rect 17694 9148 17722 9180
rect 17754 9148 17766 9180
rect 17798 9148 17810 9180
rect 17842 9148 17854 9180
rect 17886 9148 17901 9180
rect 17694 9134 17901 9148
rect -2149 8847 -2143 8875
rect -1968 8847 -1962 8875
rect 17706 8847 17712 8875
rect 17887 8847 17893 8875
rect -2149 8407 -2143 8435
rect -1968 8407 -1962 8435
rect 17706 8407 17712 8435
rect 17887 8407 17893 8435
rect -2149 7967 -2143 7995
rect -1968 7967 -1962 7995
rect 17706 7967 17712 7995
rect 17887 7967 17893 7995
rect -2149 7527 -2143 7555
rect -1968 7527 -1962 7555
rect 17706 7527 17712 7555
rect 17887 7527 17893 7555
rect -2149 7087 -2143 7115
rect -1968 7087 -1962 7115
rect 17706 7087 17712 7115
rect 17887 7087 17893 7115
rect -2149 6647 -2143 6675
rect -1968 6647 -1962 6675
rect 17706 6647 17712 6675
rect 17887 6647 17893 6675
rect -2149 6207 -2143 6235
rect -1968 6207 -1962 6235
rect 17706 6207 17712 6235
rect 17887 6207 17893 6235
rect -2149 5767 -2143 5795
rect -1968 5767 -1962 5795
rect 17706 5767 17712 5795
rect 17887 5767 17893 5795
rect -2149 5327 -2143 5355
rect -1968 5327 -1962 5355
rect 17706 5327 17712 5355
rect 17887 5327 17893 5355
rect -2149 4887 -2143 4915
rect -1968 4887 -1962 4915
rect 17706 4887 17712 4915
rect 17887 4887 17893 4915
rect -2149 4447 -2143 4475
rect -1968 4447 -1962 4475
rect 17706 4447 17712 4475
rect 17887 4447 17893 4475
rect -2149 4007 -2143 4035
rect -1968 4007 -1962 4035
rect 17706 4007 17712 4035
rect 17887 4007 17893 4035
rect -2149 3567 -2143 3595
rect -1968 3567 -1962 3595
rect 17706 3567 17712 3595
rect 17887 3567 17893 3595
rect -2149 3127 -2143 3155
rect -1968 3127 -1962 3155
rect 17706 3127 17712 3155
rect 17887 3127 17893 3155
rect -2149 2687 -2143 2715
rect -1968 2687 -1962 2715
rect 17706 2687 17712 2715
rect 17887 2687 17893 2715
rect -2149 2247 -2143 2275
rect -1968 2247 -1962 2275
rect 17706 2247 17712 2275
rect 17887 2247 17893 2275
rect -2149 1807 -2143 1835
rect -1968 1807 -1962 1835
rect 17706 1807 17712 1835
rect 17887 1807 17893 1835
rect -2149 1367 -2143 1395
rect -1968 1367 -1962 1395
rect 17706 1367 17712 1395
rect 17887 1367 17893 1395
rect -2149 927 -2143 955
rect -1968 927 -1962 955
rect 17706 927 17712 955
rect 17887 927 17893 955
rect -2149 487 -2143 515
rect -1968 487 -1962 515
rect 17706 487 17712 515
rect 17887 487 17893 515
rect -2149 47 -2143 75
rect -1968 47 -1962 75
rect 17706 47 17712 75
rect 17887 47 17893 75
rect 17694 -26 17901 -12
rect 17694 -58 17722 -26
rect 17754 -58 17766 -26
rect 17798 -58 17810 -26
rect 17842 -58 17854 -26
rect 17886 -58 17901 -26
rect 17694 -71 17901 -58
rect -2157 -91 -1950 -77
rect -2157 -123 -2142 -91
rect -2110 -123 -2098 -91
rect -2066 -123 -2054 -91
rect -2022 -123 -2010 -91
rect -1978 -123 -1950 -91
rect -2157 -136 -1950 -123
rect -2157 -168 -2142 -136
rect -2110 -168 -2098 -136
rect -2066 -168 -2054 -136
rect -2022 -168 -2010 -136
rect -1978 -168 -1950 -136
rect -2157 -181 -1950 -168
rect -2157 -213 -2142 -181
rect -2110 -213 -2098 -181
rect -2066 -213 -2054 -181
rect -2022 -213 -2010 -181
rect -1978 -213 -1950 -181
rect -2157 -217 -1950 -213
rect -273 -85 -91 -76
rect -273 -113 -241 -85
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -91 -85
rect -273 -132 -91 -113
rect -273 -160 -241 -132
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -91 -132
rect 17694 -103 17722 -71
rect 17754 -103 17766 -71
rect 17798 -103 17810 -71
rect 17842 -103 17854 -71
rect 17886 -103 17901 -71
rect 17694 -116 17901 -103
rect 17694 -148 17722 -116
rect 17754 -148 17766 -116
rect 17798 -148 17810 -116
rect 17842 -148 17854 -116
rect 17886 -148 17901 -116
rect 17694 -152 17901 -148
rect -273 -179 -91 -160
rect -273 -207 -241 -179
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -91 -179
rect -273 -217 -91 -207
rect 17989 -245 18196 -231
rect 17989 -277 18017 -245
rect 18049 -277 18061 -245
rect 18093 -277 18105 -245
rect 18137 -277 18149 -245
rect 18181 -277 18196 -245
rect 17989 -290 18196 -277
rect -2452 -310 -2245 -296
rect -2452 -342 -2437 -310
rect -2405 -342 -2393 -310
rect -2361 -342 -2349 -310
rect -2317 -342 -2305 -310
rect -2273 -342 -2245 -310
rect -2452 -355 -2245 -342
rect -2452 -387 -2437 -355
rect -2405 -387 -2393 -355
rect -2361 -387 -2349 -355
rect -2317 -387 -2305 -355
rect -2273 -387 -2245 -355
rect -2452 -400 -2245 -387
rect -2452 -432 -2437 -400
rect -2405 -432 -2393 -400
rect -2361 -432 -2349 -400
rect -2317 -432 -2305 -400
rect -2273 -432 -2245 -400
rect -2452 -436 -2245 -432
rect -462 -304 -280 -295
rect -462 -332 -430 -304
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -332 -280 -304
rect -462 -351 -280 -332
rect -462 -379 -430 -351
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -280 -351
rect 17989 -322 18017 -290
rect 18049 -322 18061 -290
rect 18093 -322 18105 -290
rect 18137 -322 18149 -290
rect 18181 -322 18196 -290
rect 17989 -335 18196 -322
rect 17989 -367 18017 -335
rect 18049 -367 18061 -335
rect 18093 -367 18105 -335
rect 18137 -367 18149 -335
rect 18181 -367 18196 -335
rect 17989 -371 18196 -367
rect -462 -398 -280 -379
rect -462 -426 -430 -398
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -280 -398
rect -462 -436 -280 -426
<< via2 >>
rect -2437 9457 -2405 9489
rect -2393 9457 -2361 9489
rect -2349 9457 -2317 9489
rect -2305 9457 -2273 9489
rect -2437 9412 -2405 9444
rect -2393 9412 -2361 9444
rect -2349 9412 -2317 9444
rect -2305 9412 -2273 9444
rect -2437 9367 -2405 9399
rect -2393 9367 -2361 9399
rect -2349 9367 -2317 9399
rect -2305 9367 -2273 9399
rect 18017 9457 18049 9489
rect 18061 9457 18093 9489
rect 18105 9457 18137 9489
rect 18149 9457 18181 9489
rect 18017 9412 18049 9444
rect 18061 9412 18093 9444
rect 18105 9412 18137 9444
rect 18149 9412 18181 9444
rect 18017 9367 18049 9399
rect 18061 9367 18093 9399
rect 18105 9367 18137 9399
rect 18149 9367 18181 9399
rect -2142 9238 -2110 9270
rect -2098 9238 -2066 9270
rect -2054 9238 -2022 9270
rect -2010 9238 -1978 9270
rect -2142 9193 -2110 9225
rect -2098 9193 -2066 9225
rect -2054 9193 -2022 9225
rect -2010 9193 -1978 9225
rect -2142 9148 -2110 9180
rect -2098 9148 -2066 9180
rect -2054 9148 -2022 9180
rect -2010 9148 -1978 9180
rect 17722 9238 17754 9270
rect 17766 9238 17798 9270
rect 17810 9238 17842 9270
rect 17854 9238 17886 9270
rect 17722 9193 17754 9225
rect 17766 9193 17798 9225
rect 17810 9193 17842 9225
rect 17854 9193 17886 9225
rect 17722 9148 17754 9180
rect 17766 9148 17798 9180
rect 17810 9148 17842 9180
rect 17854 9148 17886 9180
rect -2143 8874 -1968 8875
rect -2143 8848 -1968 8874
rect -2143 8847 -1968 8848
rect 17712 8874 17887 8875
rect 17712 8848 17887 8874
rect 17712 8847 17887 8848
rect -2143 8434 -1968 8435
rect -2143 8408 -1968 8434
rect -2143 8407 -1968 8408
rect 17712 8434 17887 8435
rect 17712 8408 17887 8434
rect 17712 8407 17887 8408
rect -2143 7994 -1968 7995
rect -2143 7968 -1968 7994
rect -2143 7967 -1968 7968
rect 17712 7994 17887 7995
rect 17712 7968 17887 7994
rect 17712 7967 17887 7968
rect -2143 7554 -1968 7555
rect -2143 7528 -1968 7554
rect -2143 7527 -1968 7528
rect 17712 7554 17887 7555
rect 17712 7528 17887 7554
rect 17712 7527 17887 7528
rect -2143 7114 -1968 7115
rect -2143 7088 -1968 7114
rect -2143 7087 -1968 7088
rect 17712 7114 17887 7115
rect 17712 7088 17887 7114
rect 17712 7087 17887 7088
rect -2143 6674 -1968 6675
rect -2143 6648 -1968 6674
rect -2143 6647 -1968 6648
rect 17712 6674 17887 6675
rect 17712 6648 17887 6674
rect 17712 6647 17887 6648
rect -2143 6234 -1968 6235
rect -2143 6208 -1968 6234
rect -2143 6207 -1968 6208
rect 17712 6234 17887 6235
rect 17712 6208 17887 6234
rect 17712 6207 17887 6208
rect -2143 5794 -1968 5795
rect -2143 5768 -1968 5794
rect -2143 5767 -1968 5768
rect 17712 5794 17887 5795
rect 17712 5768 17887 5794
rect 17712 5767 17887 5768
rect -2143 5354 -1968 5355
rect -2143 5328 -1968 5354
rect -2143 5327 -1968 5328
rect 17712 5354 17887 5355
rect 17712 5328 17887 5354
rect 17712 5327 17887 5328
rect -2143 4914 -1968 4915
rect -2143 4888 -1968 4914
rect -2143 4887 -1968 4888
rect 17712 4914 17887 4915
rect 17712 4888 17887 4914
rect 17712 4887 17887 4888
rect -2143 4474 -1968 4475
rect -2143 4448 -1968 4474
rect -2143 4447 -1968 4448
rect 17712 4474 17887 4475
rect 17712 4448 17887 4474
rect 17712 4447 17887 4448
rect -2143 4034 -1968 4035
rect -2143 4008 -1968 4034
rect -2143 4007 -1968 4008
rect 17712 4034 17887 4035
rect 17712 4008 17887 4034
rect 17712 4007 17887 4008
rect -2143 3594 -1968 3595
rect -2143 3568 -1968 3594
rect -2143 3567 -1968 3568
rect 17712 3594 17887 3595
rect 17712 3568 17887 3594
rect 17712 3567 17887 3568
rect -2143 3154 -1968 3155
rect -2143 3128 -1968 3154
rect -2143 3127 -1968 3128
rect 17712 3154 17887 3155
rect 17712 3128 17887 3154
rect 17712 3127 17887 3128
rect -2143 2714 -1968 2715
rect -2143 2688 -1968 2714
rect -2143 2687 -1968 2688
rect 17712 2714 17887 2715
rect 17712 2688 17887 2714
rect 17712 2687 17887 2688
rect -2143 2274 -1968 2275
rect -2143 2248 -1968 2274
rect -2143 2247 -1968 2248
rect 17712 2274 17887 2275
rect 17712 2248 17887 2274
rect 17712 2247 17887 2248
rect -2143 1834 -1968 1835
rect -2143 1808 -1968 1834
rect -2143 1807 -1968 1808
rect 17712 1834 17887 1835
rect 17712 1808 17887 1834
rect 17712 1807 17887 1808
rect -2143 1394 -1968 1395
rect -2143 1368 -1968 1394
rect -2143 1367 -1968 1368
rect 17712 1394 17887 1395
rect 17712 1368 17887 1394
rect 17712 1367 17887 1368
rect -2143 954 -1968 955
rect -2143 928 -1968 954
rect -2143 927 -1968 928
rect 17712 954 17887 955
rect 17712 928 17887 954
rect 17712 927 17887 928
rect -2143 514 -1968 515
rect -2143 488 -1968 514
rect -2143 487 -1968 488
rect 17712 514 17887 515
rect 17712 488 17887 514
rect 17712 487 17887 488
rect -2143 74 -1968 75
rect -2143 48 -1968 74
rect -2143 47 -1968 48
rect 17712 74 17887 75
rect 17712 48 17887 74
rect 17712 47 17887 48
rect 17722 -58 17754 -26
rect 17766 -58 17798 -26
rect 17810 -58 17842 -26
rect 17854 -58 17886 -26
rect -2142 -123 -2110 -91
rect -2098 -123 -2066 -91
rect -2054 -123 -2022 -91
rect -2010 -123 -1978 -91
rect -2142 -168 -2110 -136
rect -2098 -168 -2066 -136
rect -2054 -168 -2022 -136
rect -2010 -168 -1978 -136
rect -2142 -213 -2110 -181
rect -2098 -213 -2066 -181
rect -2054 -213 -2022 -181
rect -2010 -213 -1978 -181
rect -241 -113 -213 -85
rect -194 -113 -166 -85
rect -147 -113 -119 -85
rect -241 -160 -213 -132
rect -194 -160 -166 -132
rect -147 -160 -119 -132
rect 17722 -103 17754 -71
rect 17766 -103 17798 -71
rect 17810 -103 17842 -71
rect 17854 -103 17886 -71
rect 17722 -148 17754 -116
rect 17766 -148 17798 -116
rect 17810 -148 17842 -116
rect 17854 -148 17886 -116
rect -241 -207 -213 -179
rect -194 -207 -166 -179
rect -147 -207 -119 -179
rect 18017 -277 18049 -245
rect 18061 -277 18093 -245
rect 18105 -277 18137 -245
rect 18149 -277 18181 -245
rect -2437 -342 -2405 -310
rect -2393 -342 -2361 -310
rect -2349 -342 -2317 -310
rect -2305 -342 -2273 -310
rect -2437 -387 -2405 -355
rect -2393 -387 -2361 -355
rect -2349 -387 -2317 -355
rect -2305 -387 -2273 -355
rect -2437 -432 -2405 -400
rect -2393 -432 -2361 -400
rect -2349 -432 -2317 -400
rect -2305 -432 -2273 -400
rect -430 -332 -402 -304
rect -383 -332 -355 -304
rect -336 -332 -308 -304
rect -430 -379 -402 -351
rect -383 -379 -355 -351
rect -336 -379 -308 -351
rect 18017 -322 18049 -290
rect 18061 -322 18093 -290
rect 18105 -322 18137 -290
rect 18149 -322 18181 -290
rect 18017 -367 18049 -335
rect 18061 -367 18093 -335
rect 18105 -367 18137 -335
rect 18149 -367 18181 -335
rect -430 -426 -402 -398
rect -383 -426 -355 -398
rect -336 -426 -308 -398
<< metal3 >>
rect -2452 9489 -2245 9493
rect -2452 9457 -2437 9489
rect -2405 9457 -2393 9489
rect -2361 9457 -2349 9489
rect -2317 9457 -2305 9489
rect -2273 9457 -2245 9489
rect -2452 9444 -2245 9457
rect -2452 9412 -2437 9444
rect -2405 9412 -2393 9444
rect -2361 9412 -2349 9444
rect -2317 9412 -2305 9444
rect -2273 9412 -2245 9444
rect -2452 9399 -2245 9412
rect -2452 9367 -2437 9399
rect -2405 9367 -2393 9399
rect -2361 9367 -2349 9399
rect -2317 9367 -2305 9399
rect -2273 9367 -2245 9399
rect -2452 9353 -2245 9367
rect 17989 9489 18196 9493
rect 17989 9457 18017 9489
rect 18049 9457 18061 9489
rect 18093 9457 18105 9489
rect 18137 9457 18149 9489
rect 18181 9457 18196 9489
rect 17989 9444 18196 9457
rect 17989 9412 18017 9444
rect 18049 9412 18061 9444
rect 18093 9412 18105 9444
rect 18137 9412 18149 9444
rect 18181 9412 18196 9444
rect 17989 9399 18196 9412
rect 17989 9367 18017 9399
rect 18049 9367 18061 9399
rect 18093 9367 18105 9399
rect 18137 9367 18149 9399
rect 18181 9367 18196 9399
rect 17989 9353 18196 9367
rect -2157 9270 -1950 9274
rect -2157 9238 -2142 9270
rect -2110 9238 -2098 9270
rect -2066 9238 -2054 9270
rect -2022 9238 -2010 9270
rect -1978 9238 -1950 9270
rect -2157 9225 -1950 9238
rect -2157 9193 -2142 9225
rect -2110 9193 -2098 9225
rect -2066 9193 -2054 9225
rect -2022 9193 -2010 9225
rect -1978 9193 -1950 9225
rect -2157 9180 -1950 9193
rect -2157 9148 -2142 9180
rect -2110 9148 -2098 9180
rect -2066 9148 -2054 9180
rect -2022 9148 -2010 9180
rect -1978 9148 -1950 9180
rect -2157 9134 -1950 9148
rect 17694 9270 17901 9274
rect 17694 9238 17722 9270
rect 17754 9238 17766 9270
rect 17798 9238 17810 9270
rect 17842 9238 17854 9270
rect 17886 9238 17901 9270
rect 17694 9225 17901 9238
rect 17694 9193 17722 9225
rect 17754 9193 17766 9225
rect 17798 9193 17810 9225
rect 17842 9193 17854 9225
rect 17886 9193 17901 9225
rect 17694 9180 17901 9193
rect 17694 9148 17722 9180
rect 17754 9148 17766 9180
rect 17798 9148 17810 9180
rect 17842 9148 17854 9180
rect 17886 9148 17901 9180
rect 17694 9134 17901 9148
rect -2149 8877 -1962 8878
rect -2149 8845 -2143 8877
rect -1968 8845 -1962 8877
rect -2149 8844 -1962 8845
rect 17706 8877 17893 8878
rect 17706 8845 17712 8877
rect 17887 8845 17893 8877
rect 17706 8844 17893 8845
rect -2149 8437 -1962 8438
rect -2149 8405 -2143 8437
rect -1968 8405 -1962 8437
rect -2149 8404 -1962 8405
rect 17706 8437 17893 8438
rect 17706 8405 17712 8437
rect 17887 8405 17893 8437
rect 17706 8404 17893 8405
rect -2149 7997 -1962 7998
rect -2149 7965 -2143 7997
rect -1968 7965 -1962 7997
rect -2149 7964 -1962 7965
rect 17706 7997 17893 7998
rect 17706 7965 17712 7997
rect 17887 7965 17893 7997
rect 17706 7964 17893 7965
rect -2149 7557 -1962 7558
rect -2149 7525 -2143 7557
rect -1968 7525 -1962 7557
rect -2149 7524 -1962 7525
rect 17706 7557 17893 7558
rect 17706 7525 17712 7557
rect 17887 7525 17893 7557
rect 17706 7524 17893 7525
rect -2149 7117 -1962 7118
rect -2149 7085 -2143 7117
rect -1968 7085 -1962 7117
rect -2149 7084 -1962 7085
rect 17706 7117 17893 7118
rect 17706 7085 17712 7117
rect 17887 7085 17893 7117
rect 17706 7084 17893 7085
rect -2149 6677 -1962 6678
rect -2149 6645 -2143 6677
rect -1968 6645 -1962 6677
rect -2149 6644 -1962 6645
rect 17706 6677 17893 6678
rect 17706 6645 17712 6677
rect 17887 6645 17893 6677
rect 17706 6644 17893 6645
rect -2149 6237 -1962 6238
rect -2149 6205 -2143 6237
rect -1968 6205 -1962 6237
rect -2149 6204 -1962 6205
rect 17706 6237 17893 6238
rect 17706 6205 17712 6237
rect 17887 6205 17893 6237
rect 17706 6204 17893 6205
rect -2149 5797 -1962 5798
rect -2149 5765 -2143 5797
rect -1968 5765 -1962 5797
rect -2149 5764 -1962 5765
rect 17706 5797 17893 5798
rect 17706 5765 17712 5797
rect 17887 5765 17893 5797
rect 17706 5764 17893 5765
rect -2149 5357 -1962 5358
rect -2149 5325 -2143 5357
rect -1968 5325 -1962 5357
rect -2149 5324 -1962 5325
rect 17706 5357 17893 5358
rect 17706 5325 17712 5357
rect 17887 5325 17893 5357
rect 17706 5324 17893 5325
rect -2149 4917 -1962 4918
rect -2149 4885 -2143 4917
rect -1968 4885 -1962 4917
rect -2149 4884 -1962 4885
rect 17706 4917 17893 4918
rect 17706 4885 17712 4917
rect 17887 4885 17893 4917
rect 17706 4884 17893 4885
rect -2149 4477 -1962 4478
rect -2149 4445 -2143 4477
rect -1968 4445 -1962 4477
rect -2149 4444 -1962 4445
rect 17706 4477 17893 4478
rect 17706 4445 17712 4477
rect 17887 4445 17893 4477
rect 17706 4444 17893 4445
rect -2149 4037 -1962 4038
rect -2149 4005 -2143 4037
rect -1968 4005 -1962 4037
rect -2149 4004 -1962 4005
rect 17706 4037 17893 4038
rect 17706 4005 17712 4037
rect 17887 4005 17893 4037
rect 17706 4004 17893 4005
rect -2149 3597 -1962 3598
rect -2149 3565 -2143 3597
rect -1968 3565 -1962 3597
rect -2149 3564 -1962 3565
rect 17706 3597 17893 3598
rect 17706 3565 17712 3597
rect 17887 3565 17893 3597
rect 17706 3564 17893 3565
rect -2149 3157 -1962 3158
rect -2149 3125 -2143 3157
rect -1968 3125 -1962 3157
rect -2149 3124 -1962 3125
rect 17706 3157 17893 3158
rect 17706 3125 17712 3157
rect 17887 3125 17893 3157
rect 17706 3124 17893 3125
rect -2149 2717 -1962 2718
rect -2149 2685 -2143 2717
rect -1968 2685 -1962 2717
rect -2149 2684 -1962 2685
rect 17706 2717 17893 2718
rect 17706 2685 17712 2717
rect 17887 2685 17893 2717
rect 17706 2684 17893 2685
rect -2149 2277 -1962 2278
rect -2149 2245 -2143 2277
rect -1968 2245 -1962 2277
rect -2149 2244 -1962 2245
rect 17706 2277 17893 2278
rect 17706 2245 17712 2277
rect 17887 2245 17893 2277
rect 17706 2244 17893 2245
rect -2149 1837 -1962 1838
rect -2149 1805 -2143 1837
rect -1968 1805 -1962 1837
rect -2149 1804 -1962 1805
rect 17706 1837 17893 1838
rect 17706 1805 17712 1837
rect 17887 1805 17893 1837
rect 17706 1804 17893 1805
rect -2149 1397 -1962 1398
rect -2149 1365 -2143 1397
rect -1968 1365 -1962 1397
rect -2149 1364 -1962 1365
rect 17706 1397 17893 1398
rect 17706 1365 17712 1397
rect 17887 1365 17893 1397
rect 17706 1364 17893 1365
rect -2149 957 -1962 958
rect -2149 925 -2143 957
rect -1968 925 -1962 957
rect -2149 924 -1962 925
rect 17706 957 17893 958
rect 17706 925 17712 957
rect 17887 925 17893 957
rect 17706 924 17893 925
rect -2149 517 -1962 518
rect -2149 485 -2143 517
rect -1968 485 -1962 517
rect -2149 484 -1962 485
rect 17706 517 17893 518
rect 17706 485 17712 517
rect 17887 485 17893 517
rect 17706 484 17893 485
rect -2149 77 -1962 78
rect -2149 45 -2143 77
rect -1968 45 -1962 77
rect -2149 44 -1962 45
rect 17706 77 17893 78
rect 17706 45 17712 77
rect 17887 45 17893 77
rect 17706 44 17893 45
rect 17694 -26 17901 -12
rect 17694 -58 17722 -26
rect 17754 -58 17766 -26
rect 17798 -58 17810 -26
rect 17842 -58 17854 -26
rect 17886 -58 17901 -26
rect 17694 -71 17901 -58
rect -2158 -85 -91 -76
rect -2158 -91 -241 -85
rect -2158 -123 -2142 -91
rect -2110 -123 -2098 -91
rect -2066 -123 -2054 -91
rect -2022 -123 -2010 -91
rect -1978 -113 -241 -91
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -91 -85
rect -1978 -123 -91 -113
rect -2158 -132 -91 -123
rect -2158 -136 -241 -132
rect -2158 -168 -2142 -136
rect -2110 -168 -2098 -136
rect -2066 -168 -2054 -136
rect -2022 -168 -2010 -136
rect -1978 -160 -241 -136
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -91 -132
rect 17694 -103 17722 -71
rect 17754 -103 17766 -71
rect 17798 -103 17810 -71
rect 17842 -103 17854 -71
rect 17886 -103 17901 -71
rect 17694 -116 17901 -103
rect 17694 -148 17722 -116
rect 17754 -148 17766 -116
rect 17798 -148 17810 -116
rect 17842 -148 17854 -116
rect 17886 -148 17901 -116
rect 17694 -152 17901 -148
rect -1978 -168 -91 -160
rect -2158 -179 -91 -168
rect -2158 -181 -241 -179
rect -2158 -213 -2142 -181
rect -2110 -213 -2098 -181
rect -2066 -213 -2054 -181
rect -2022 -213 -2010 -181
rect -1978 -207 -241 -181
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -91 -179
rect -1978 -213 -91 -207
rect -2158 -217 -91 -213
rect 17989 -245 18196 -231
rect 17989 -277 18017 -245
rect 18049 -277 18061 -245
rect 18093 -277 18105 -245
rect 18137 -277 18149 -245
rect 18181 -277 18196 -245
rect 17989 -290 18196 -277
rect -2245 -296 -280 -295
rect -2452 -304 -280 -296
rect -2452 -310 -430 -304
rect -2452 -342 -2437 -310
rect -2405 -342 -2393 -310
rect -2361 -342 -2349 -310
rect -2317 -342 -2305 -310
rect -2273 -332 -430 -310
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -332 -280 -304
rect -2273 -342 -280 -332
rect -2452 -351 -280 -342
rect -2452 -355 -430 -351
rect -2452 -387 -2437 -355
rect -2405 -387 -2393 -355
rect -2361 -387 -2349 -355
rect -2317 -387 -2305 -355
rect -2273 -379 -430 -355
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -280 -351
rect 17989 -322 18017 -290
rect 18049 -322 18061 -290
rect 18093 -322 18105 -290
rect 18137 -322 18149 -290
rect 18181 -322 18196 -290
rect 17989 -335 18196 -322
rect 17989 -367 18017 -335
rect 18049 -367 18061 -335
rect 18093 -367 18105 -335
rect 18137 -367 18149 -335
rect 18181 -367 18196 -335
rect 17989 -371 18196 -367
rect -2273 -387 -280 -379
rect -2452 -398 -280 -387
rect -2452 -400 -430 -398
rect -2452 -432 -2437 -400
rect -2405 -432 -2393 -400
rect -2361 -432 -2349 -400
rect -2317 -432 -2305 -400
rect -2273 -426 -430 -400
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -280 -398
rect -2273 -432 -280 -426
rect -2452 -436 -280 -432
<< via3 >>
rect -2437 9457 -2405 9489
rect -2393 9457 -2361 9489
rect -2349 9457 -2317 9489
rect -2305 9457 -2273 9489
rect -2437 9412 -2405 9444
rect -2393 9412 -2361 9444
rect -2349 9412 -2317 9444
rect -2305 9412 -2273 9444
rect -2437 9367 -2405 9399
rect -2393 9367 -2361 9399
rect -2349 9367 -2317 9399
rect -2305 9367 -2273 9399
rect 18017 9457 18049 9489
rect 18061 9457 18093 9489
rect 18105 9457 18137 9489
rect 18149 9457 18181 9489
rect 18017 9412 18049 9444
rect 18061 9412 18093 9444
rect 18105 9412 18137 9444
rect 18149 9412 18181 9444
rect 18017 9367 18049 9399
rect 18061 9367 18093 9399
rect 18105 9367 18137 9399
rect 18149 9367 18181 9399
rect -2142 9238 -2110 9270
rect -2098 9238 -2066 9270
rect -2054 9238 -2022 9270
rect -2010 9238 -1978 9270
rect -2142 9193 -2110 9225
rect -2098 9193 -2066 9225
rect -2054 9193 -2022 9225
rect -2010 9193 -1978 9225
rect -2142 9148 -2110 9180
rect -2098 9148 -2066 9180
rect -2054 9148 -2022 9180
rect -2010 9148 -1978 9180
rect 17722 9238 17754 9270
rect 17766 9238 17798 9270
rect 17810 9238 17842 9270
rect 17854 9238 17886 9270
rect 17722 9193 17754 9225
rect 17766 9193 17798 9225
rect 17810 9193 17842 9225
rect 17854 9193 17886 9225
rect 17722 9148 17754 9180
rect 17766 9148 17798 9180
rect 17810 9148 17842 9180
rect 17854 9148 17886 9180
rect -2143 8875 -1968 8877
rect -2143 8847 -1968 8875
rect -2143 8845 -1968 8847
rect 17712 8875 17887 8877
rect 17712 8847 17887 8875
rect 17712 8845 17887 8847
rect -2143 8435 -1968 8437
rect -2143 8407 -1968 8435
rect -2143 8405 -1968 8407
rect 17712 8435 17887 8437
rect 17712 8407 17887 8435
rect 17712 8405 17887 8407
rect -2143 7995 -1968 7997
rect -2143 7967 -1968 7995
rect -2143 7965 -1968 7967
rect 17712 7995 17887 7997
rect 17712 7967 17887 7995
rect 17712 7965 17887 7967
rect -2143 7555 -1968 7557
rect -2143 7527 -1968 7555
rect -2143 7525 -1968 7527
rect 17712 7555 17887 7557
rect 17712 7527 17887 7555
rect 17712 7525 17887 7527
rect -2143 7115 -1968 7117
rect -2143 7087 -1968 7115
rect -2143 7085 -1968 7087
rect 17712 7115 17887 7117
rect 17712 7087 17887 7115
rect 17712 7085 17887 7087
rect -2143 6675 -1968 6677
rect -2143 6647 -1968 6675
rect -2143 6645 -1968 6647
rect 17712 6675 17887 6677
rect 17712 6647 17887 6675
rect 17712 6645 17887 6647
rect -2143 6235 -1968 6237
rect -2143 6207 -1968 6235
rect -2143 6205 -1968 6207
rect 17712 6235 17887 6237
rect 17712 6207 17887 6235
rect 17712 6205 17887 6207
rect -2143 5795 -1968 5797
rect -2143 5767 -1968 5795
rect -2143 5765 -1968 5767
rect 17712 5795 17887 5797
rect 17712 5767 17887 5795
rect 17712 5765 17887 5767
rect -2143 5355 -1968 5357
rect -2143 5327 -1968 5355
rect -2143 5325 -1968 5327
rect 17712 5355 17887 5357
rect 17712 5327 17887 5355
rect 17712 5325 17887 5327
rect -2143 4915 -1968 4917
rect -2143 4887 -1968 4915
rect -2143 4885 -1968 4887
rect 17712 4915 17887 4917
rect 17712 4887 17887 4915
rect 17712 4885 17887 4887
rect -2143 4475 -1968 4477
rect -2143 4447 -1968 4475
rect -2143 4445 -1968 4447
rect 17712 4475 17887 4477
rect 17712 4447 17887 4475
rect 17712 4445 17887 4447
rect -2143 4035 -1968 4037
rect -2143 4007 -1968 4035
rect -2143 4005 -1968 4007
rect 17712 4035 17887 4037
rect 17712 4007 17887 4035
rect 17712 4005 17887 4007
rect -2143 3595 -1968 3597
rect -2143 3567 -1968 3595
rect -2143 3565 -1968 3567
rect 17712 3595 17887 3597
rect 17712 3567 17887 3595
rect 17712 3565 17887 3567
rect -2143 3155 -1968 3157
rect -2143 3127 -1968 3155
rect -2143 3125 -1968 3127
rect 17712 3155 17887 3157
rect 17712 3127 17887 3155
rect 17712 3125 17887 3127
rect -2143 2715 -1968 2717
rect -2143 2687 -1968 2715
rect -2143 2685 -1968 2687
rect 17712 2715 17887 2717
rect 17712 2687 17887 2715
rect 17712 2685 17887 2687
rect -2143 2275 -1968 2277
rect -2143 2247 -1968 2275
rect -2143 2245 -1968 2247
rect 17712 2275 17887 2277
rect 17712 2247 17887 2275
rect 17712 2245 17887 2247
rect -2143 1835 -1968 1837
rect -2143 1807 -1968 1835
rect -2143 1805 -1968 1807
rect 17712 1835 17887 1837
rect 17712 1807 17887 1835
rect 17712 1805 17887 1807
rect -2143 1395 -1968 1397
rect -2143 1367 -1968 1395
rect -2143 1365 -1968 1367
rect 17712 1395 17887 1397
rect 17712 1367 17887 1395
rect 17712 1365 17887 1367
rect -2143 955 -1968 957
rect -2143 927 -1968 955
rect -2143 925 -1968 927
rect 17712 955 17887 957
rect 17712 927 17887 955
rect 17712 925 17887 927
rect -2143 515 -1968 517
rect -2143 487 -1968 515
rect -2143 485 -1968 487
rect 17712 515 17887 517
rect 17712 487 17887 515
rect 17712 485 17887 487
rect -2143 75 -1968 77
rect -2143 47 -1968 75
rect -2143 45 -1968 47
rect 17712 75 17887 77
rect 17712 47 17887 75
rect 17712 45 17887 47
rect 17722 -58 17754 -26
rect 17766 -58 17798 -26
rect 17810 -58 17842 -26
rect 17854 -58 17886 -26
rect -2142 -123 -2110 -91
rect -2098 -123 -2066 -91
rect -2054 -123 -2022 -91
rect -2010 -123 -1978 -91
rect -2142 -168 -2110 -136
rect -2098 -168 -2066 -136
rect -2054 -168 -2022 -136
rect -2010 -168 -1978 -136
rect 17722 -103 17754 -71
rect 17766 -103 17798 -71
rect 17810 -103 17842 -71
rect 17854 -103 17886 -71
rect 17722 -148 17754 -116
rect 17766 -148 17798 -116
rect 17810 -148 17842 -116
rect 17854 -148 17886 -116
rect -2142 -213 -2110 -181
rect -2098 -213 -2066 -181
rect -2054 -213 -2022 -181
rect -2010 -213 -1978 -181
rect 18017 -277 18049 -245
rect 18061 -277 18093 -245
rect 18105 -277 18137 -245
rect 18149 -277 18181 -245
rect -2437 -342 -2405 -310
rect -2393 -342 -2361 -310
rect -2349 -342 -2317 -310
rect -2305 -342 -2273 -310
rect -2437 -387 -2405 -355
rect -2393 -387 -2361 -355
rect -2349 -387 -2317 -355
rect -2305 -387 -2273 -355
rect 18017 -322 18049 -290
rect 18061 -322 18093 -290
rect 18105 -322 18137 -290
rect 18149 -322 18181 -290
rect 18017 -367 18049 -335
rect 18061 -367 18093 -335
rect 18105 -367 18137 -335
rect 18149 -367 18181 -335
rect -2437 -432 -2405 -400
rect -2393 -432 -2361 -400
rect -2349 -432 -2317 -400
rect -2305 -432 -2273 -400
<< metal4 >>
rect -2452 9489 -2245 9494
rect -2452 9457 -2437 9489
rect -2405 9457 -2393 9489
rect -2361 9457 -2349 9489
rect -2317 9457 -2305 9489
rect -2273 9457 -2245 9489
rect -2452 9444 -2245 9457
rect -2452 9412 -2437 9444
rect -2405 9412 -2393 9444
rect -2361 9412 -2349 9444
rect -2317 9412 -2305 9444
rect -2273 9412 -2245 9444
rect -2452 9399 -2245 9412
rect -2452 9367 -2437 9399
rect -2405 9367 -2393 9399
rect -2361 9367 -2349 9399
rect -2317 9367 -2305 9399
rect -2273 9367 -2245 9399
rect -2452 -310 -2245 9367
rect -2157 9270 -1950 9494
rect -2157 9238 -2142 9270
rect -2110 9238 -2098 9270
rect -2066 9238 -2054 9270
rect -2022 9238 -2010 9270
rect -1978 9238 -1950 9270
rect -2157 9225 -1950 9238
rect -2157 9193 -2142 9225
rect -2110 9193 -2098 9225
rect -2066 9193 -2054 9225
rect -2022 9193 -2010 9225
rect -1978 9193 -1950 9225
rect -2157 9180 -1950 9193
rect -2157 9148 -2142 9180
rect -2110 9148 -2098 9180
rect -2066 9148 -2054 9180
rect -2022 9148 -2010 9180
rect -1978 9148 -1950 9180
rect -2157 8877 -1950 9148
rect -2157 8845 -2143 8877
rect -1968 8845 -1950 8877
rect -2157 8437 -1950 8845
rect 17694 9270 17901 9494
rect 17694 9238 17722 9270
rect 17754 9238 17766 9270
rect 17798 9238 17810 9270
rect 17842 9238 17854 9270
rect 17886 9238 17901 9270
rect 17694 9225 17901 9238
rect 17694 9193 17722 9225
rect 17754 9193 17766 9225
rect 17798 9193 17810 9225
rect 17842 9193 17854 9225
rect 17886 9193 17901 9225
rect 17694 9180 17901 9193
rect 17694 9148 17722 9180
rect 17754 9148 17766 9180
rect 17798 9148 17810 9180
rect 17842 9148 17854 9180
rect 17886 9148 17901 9180
rect 17694 8877 17901 9148
rect 17694 8845 17712 8877
rect 17887 8845 17901 8877
rect -2157 8405 -2143 8437
rect -1968 8405 -1950 8437
rect 969 8412 1039 8442
rect 1471 8412 1541 8442
rect 1973 8412 2043 8442
rect 2475 8412 2545 8442
rect 2977 8412 3047 8442
rect 3479 8412 3549 8442
rect 3981 8412 4051 8442
rect 4483 8412 4553 8442
rect 4985 8412 5055 8442
rect 5487 8412 5557 8442
rect 5989 8412 6059 8442
rect 6491 8412 6561 8442
rect 6993 8412 7063 8442
rect 7495 8412 7565 8442
rect 7997 8412 8067 8442
rect 8499 8412 8569 8442
rect 9001 8412 9071 8442
rect 9503 8412 9573 8442
rect 10005 8412 10075 8442
rect 10507 8412 10577 8442
rect 11009 8412 11079 8442
rect 11511 8412 11581 8442
rect 12013 8412 12083 8442
rect 12515 8412 12585 8442
rect 13017 8412 13087 8442
rect 13519 8412 13589 8442
rect 14021 8412 14091 8442
rect 14523 8412 14593 8442
rect 15025 8412 15095 8442
rect 15527 8412 15597 8442
rect 16029 8412 16099 8442
rect 17694 8437 17901 8845
rect -2157 7997 -1950 8405
rect 17694 8405 17712 8437
rect 17887 8405 17901 8437
rect 969 8124 1039 8154
rect 1471 8124 1541 8154
rect 1973 8124 2043 8154
rect 2475 8124 2545 8154
rect 2977 8124 3047 8154
rect 3479 8124 3549 8154
rect 3981 8124 4051 8154
rect 4483 8124 4553 8154
rect 4985 8124 5055 8154
rect 5487 8124 5557 8154
rect 5989 8124 6059 8154
rect 6491 8124 6561 8154
rect 6993 8124 7063 8154
rect 7495 8124 7565 8154
rect 7997 8124 8067 8154
rect 8499 8124 8569 8154
rect 9001 8124 9071 8154
rect 9503 8124 9573 8154
rect 10005 8124 10075 8154
rect 10507 8124 10577 8154
rect 11009 8124 11079 8154
rect 11511 8124 11581 8154
rect 12013 8124 12083 8154
rect 12515 8124 12585 8154
rect 13017 8124 13087 8154
rect 13519 8124 13589 8154
rect 14021 8124 14091 8154
rect 14523 8124 14593 8154
rect 15025 8124 15095 8154
rect 15527 8124 15597 8154
rect 16029 8124 16099 8154
rect 594 7997 624 8067
rect 882 7997 912 8067
rect 1096 7997 1126 8067
rect 1384 7997 1414 8067
rect 1598 7997 1628 8067
rect 1886 7997 1916 8067
rect 2100 7997 2130 8067
rect 2388 7997 2418 8067
rect 2602 7997 2632 8067
rect 2890 7997 2920 8067
rect 3104 7997 3134 8067
rect 3392 7997 3422 8067
rect 3606 7997 3636 8067
rect 3894 7997 3924 8067
rect 4108 7997 4138 8067
rect 4396 7997 4426 8067
rect 4610 7997 4640 8067
rect 4898 7997 4928 8067
rect 5112 7997 5142 8067
rect 5400 7997 5430 8067
rect 5614 7997 5644 8067
rect 5902 7997 5932 8067
rect 6116 7997 6146 8067
rect 6404 7997 6434 8067
rect 6618 7997 6648 8067
rect 6906 7997 6936 8067
rect 7120 7997 7150 8067
rect 7408 7997 7438 8067
rect 7622 7997 7652 8067
rect 7910 7997 7940 8067
rect 8124 7997 8154 8067
rect 8412 7997 8442 8067
rect 8626 7997 8656 8067
rect 8914 7997 8944 8067
rect 9128 7997 9158 8067
rect 9416 7997 9446 8067
rect 9630 7997 9660 8067
rect 9918 7997 9948 8067
rect 10132 7997 10162 8067
rect 10420 7997 10450 8067
rect 10634 7997 10664 8067
rect 10922 7997 10952 8067
rect 11136 7997 11166 8067
rect 11424 7997 11454 8067
rect 11638 7997 11668 8067
rect 11926 7997 11956 8067
rect 12140 7997 12170 8067
rect 12428 7997 12458 8067
rect 12642 7997 12672 8067
rect 12930 7997 12960 8067
rect 13144 7997 13174 8067
rect 13432 7997 13462 8067
rect 13646 7997 13676 8067
rect 13934 7997 13964 8067
rect 14148 7997 14178 8067
rect 14436 7997 14466 8067
rect 14650 7997 14680 8067
rect 14938 7997 14968 8067
rect 15152 7997 15182 8067
rect 15440 7997 15470 8067
rect 15654 7997 15684 8067
rect 15942 7997 15972 8067
rect 16156 7997 16186 8067
rect 16444 7997 16474 8067
rect 17694 7997 17901 8405
rect -2157 7965 -2143 7997
rect -1968 7965 -1950 7997
rect -2157 7557 -1950 7965
rect 17694 7965 17712 7997
rect 17887 7965 17901 7997
rect 969 7910 1039 7940
rect 1471 7910 1541 7940
rect 1973 7910 2043 7940
rect 2475 7910 2545 7940
rect 2977 7910 3047 7940
rect 3479 7910 3549 7940
rect 3981 7910 4051 7940
rect 4483 7910 4553 7940
rect 4985 7910 5055 7940
rect 5487 7910 5557 7940
rect 5989 7910 6059 7940
rect 6491 7910 6561 7940
rect 6993 7910 7063 7940
rect 7495 7910 7565 7940
rect 7997 7910 8067 7940
rect 8499 7910 8569 7940
rect 9001 7910 9071 7940
rect 9503 7910 9573 7940
rect 10005 7910 10075 7940
rect 10507 7910 10577 7940
rect 11009 7910 11079 7940
rect 11511 7910 11581 7940
rect 12013 7910 12083 7940
rect 12515 7910 12585 7940
rect 13017 7910 13087 7940
rect 13519 7910 13589 7940
rect 14021 7910 14091 7940
rect 14523 7910 14593 7940
rect 15025 7910 15095 7940
rect 15527 7910 15597 7940
rect 16029 7910 16099 7940
rect 969 7622 1039 7652
rect 1471 7622 1541 7652
rect 1973 7622 2043 7652
rect 2475 7622 2545 7652
rect 2977 7622 3047 7652
rect 3479 7622 3549 7652
rect 3981 7622 4051 7652
rect 4483 7622 4553 7652
rect 4985 7622 5055 7652
rect 5487 7622 5557 7652
rect 5989 7622 6059 7652
rect 6491 7622 6561 7652
rect 6993 7622 7063 7652
rect 7495 7622 7565 7652
rect 7997 7622 8067 7652
rect 8499 7622 8569 7652
rect 9001 7622 9071 7652
rect 9503 7622 9573 7652
rect 10005 7622 10075 7652
rect 10507 7622 10577 7652
rect 11009 7622 11079 7652
rect 11511 7622 11581 7652
rect 12013 7622 12083 7652
rect 12515 7622 12585 7652
rect 13017 7622 13087 7652
rect 13519 7622 13589 7652
rect 14021 7622 14091 7652
rect 14523 7622 14593 7652
rect 15025 7622 15095 7652
rect 15527 7622 15597 7652
rect 16029 7622 16099 7652
rect -2157 7525 -2143 7557
rect -1968 7525 -1950 7557
rect -2157 7117 -1950 7525
rect 594 7495 624 7565
rect 882 7495 912 7565
rect 1096 7495 1126 7565
rect 1384 7495 1414 7565
rect 1598 7495 1628 7565
rect 1886 7495 1916 7565
rect 2100 7495 2130 7565
rect 2388 7495 2418 7565
rect 2602 7495 2632 7565
rect 2890 7495 2920 7565
rect 3104 7495 3134 7565
rect 3392 7495 3422 7565
rect 3606 7495 3636 7565
rect 3894 7495 3924 7565
rect 4108 7495 4138 7565
rect 4396 7495 4426 7565
rect 4610 7495 4640 7565
rect 4898 7495 4928 7565
rect 5112 7495 5142 7565
rect 5400 7495 5430 7565
rect 5614 7495 5644 7565
rect 5902 7495 5932 7565
rect 6116 7495 6146 7565
rect 6404 7495 6434 7565
rect 6618 7495 6648 7565
rect 6906 7495 6936 7565
rect 7120 7495 7150 7565
rect 7408 7495 7438 7565
rect 7622 7495 7652 7565
rect 7910 7495 7940 7565
rect 8124 7495 8154 7565
rect 8412 7495 8442 7565
rect 8626 7495 8656 7565
rect 8914 7495 8944 7565
rect 9128 7495 9158 7565
rect 9416 7495 9446 7565
rect 9630 7495 9660 7565
rect 9918 7495 9948 7565
rect 10132 7495 10162 7565
rect 10420 7495 10450 7565
rect 10634 7495 10664 7565
rect 10922 7495 10952 7565
rect 11136 7495 11166 7565
rect 11424 7495 11454 7565
rect 11638 7495 11668 7565
rect 11926 7495 11956 7565
rect 12140 7495 12170 7565
rect 12428 7495 12458 7565
rect 12642 7495 12672 7565
rect 12930 7495 12960 7565
rect 13144 7495 13174 7565
rect 13432 7495 13462 7565
rect 13646 7495 13676 7565
rect 13934 7495 13964 7565
rect 14148 7495 14178 7565
rect 14436 7495 14466 7565
rect 14650 7495 14680 7565
rect 14938 7495 14968 7565
rect 15152 7495 15182 7565
rect 15440 7495 15470 7565
rect 15654 7495 15684 7565
rect 15942 7495 15972 7565
rect 16156 7495 16186 7565
rect 16444 7495 16474 7565
rect 17694 7557 17901 7965
rect 17694 7525 17712 7557
rect 17887 7525 17901 7557
rect 969 7408 1039 7438
rect 1471 7408 1541 7438
rect 1973 7408 2043 7438
rect 2475 7408 2545 7438
rect 2977 7408 3047 7438
rect 3479 7408 3549 7438
rect 3981 7408 4051 7438
rect 4483 7408 4553 7438
rect 4985 7408 5055 7438
rect 5487 7408 5557 7438
rect 5989 7408 6059 7438
rect 6491 7408 6561 7438
rect 6993 7408 7063 7438
rect 7495 7408 7565 7438
rect 7997 7408 8067 7438
rect 8499 7408 8569 7438
rect 9001 7408 9071 7438
rect 9503 7408 9573 7438
rect 10005 7408 10075 7438
rect 10507 7408 10577 7438
rect 11009 7408 11079 7438
rect 11511 7408 11581 7438
rect 12013 7408 12083 7438
rect 12515 7408 12585 7438
rect 13017 7408 13087 7438
rect 13519 7408 13589 7438
rect 14021 7408 14091 7438
rect 14523 7408 14593 7438
rect 15025 7408 15095 7438
rect 15527 7408 15597 7438
rect 16029 7408 16099 7438
rect 969 7120 1039 7150
rect 1471 7120 1541 7150
rect 1973 7120 2043 7150
rect 2475 7120 2545 7150
rect 2977 7120 3047 7150
rect 3479 7120 3549 7150
rect 3981 7120 4051 7150
rect 4483 7120 4553 7150
rect 4985 7120 5055 7150
rect 5487 7120 5557 7150
rect 5989 7120 6059 7150
rect 6491 7120 6561 7150
rect 6993 7120 7063 7150
rect 7495 7120 7565 7150
rect 7997 7120 8067 7150
rect 8499 7120 8569 7150
rect 9001 7120 9071 7150
rect 9503 7120 9573 7150
rect 10005 7120 10075 7150
rect 10507 7120 10577 7150
rect 11009 7120 11079 7150
rect 11511 7120 11581 7150
rect 12013 7120 12083 7150
rect 12515 7120 12585 7150
rect 13017 7120 13087 7150
rect 13519 7120 13589 7150
rect 14021 7120 14091 7150
rect 14523 7120 14593 7150
rect 15025 7120 15095 7150
rect 15527 7120 15597 7150
rect 16029 7120 16099 7150
rect -2157 7085 -2143 7117
rect -1968 7085 -1950 7117
rect -2157 6677 -1950 7085
rect 17694 7117 17901 7525
rect 17694 7085 17712 7117
rect 17887 7085 17901 7117
rect 594 6993 624 7063
rect 882 6993 912 7063
rect 1096 6993 1126 7063
rect 1384 6993 1414 7063
rect 1598 6993 1628 7063
rect 1886 6993 1916 7063
rect 2100 6993 2130 7063
rect 2388 6993 2418 7063
rect 2602 6993 2632 7063
rect 2890 6993 2920 7063
rect 3104 6993 3134 7063
rect 3392 6993 3422 7063
rect 3606 6993 3636 7063
rect 3894 6993 3924 7063
rect 4108 6993 4138 7063
rect 4396 6993 4426 7063
rect 4610 6993 4640 7063
rect 4898 6993 4928 7063
rect 5112 6993 5142 7063
rect 5400 6993 5430 7063
rect 5614 6993 5644 7063
rect 5902 6993 5932 7063
rect 6116 6993 6146 7063
rect 6404 6993 6434 7063
rect 6618 6993 6648 7063
rect 6906 6993 6936 7063
rect 7120 6993 7150 7063
rect 7408 6993 7438 7063
rect 7622 6993 7652 7063
rect 7910 6993 7940 7063
rect 8124 6993 8154 7063
rect 8412 6993 8442 7063
rect 8626 6993 8656 7063
rect 8914 6993 8944 7063
rect 9128 6993 9158 7063
rect 9416 6993 9446 7063
rect 9630 6993 9660 7063
rect 9918 6993 9948 7063
rect 10132 6993 10162 7063
rect 10420 6993 10450 7063
rect 10634 6993 10664 7063
rect 10922 6993 10952 7063
rect 11136 6993 11166 7063
rect 11424 6993 11454 7063
rect 11638 6993 11668 7063
rect 11926 6993 11956 7063
rect 12140 6993 12170 7063
rect 12428 6993 12458 7063
rect 12642 6993 12672 7063
rect 12930 6993 12960 7063
rect 13144 6993 13174 7063
rect 13432 6993 13462 7063
rect 13646 6993 13676 7063
rect 13934 6993 13964 7063
rect 14148 6993 14178 7063
rect 14436 6993 14466 7063
rect 14650 6993 14680 7063
rect 14938 6993 14968 7063
rect 15152 6993 15182 7063
rect 15440 6993 15470 7063
rect 15654 6993 15684 7063
rect 15942 6993 15972 7063
rect 16156 6993 16186 7063
rect 16444 6993 16474 7063
rect 969 6906 1039 6936
rect 1471 6906 1541 6936
rect 1973 6906 2043 6936
rect 2475 6906 2545 6936
rect 2977 6906 3047 6936
rect 3479 6906 3549 6936
rect 3981 6906 4051 6936
rect 4483 6906 4553 6936
rect 4985 6906 5055 6936
rect 5487 6906 5557 6936
rect 5989 6906 6059 6936
rect 6491 6906 6561 6936
rect 6993 6906 7063 6936
rect 7495 6906 7565 6936
rect 7997 6906 8067 6936
rect 8499 6906 8569 6936
rect 9001 6906 9071 6936
rect 9503 6906 9573 6936
rect 10005 6906 10075 6936
rect 10507 6906 10577 6936
rect 11009 6906 11079 6936
rect 11511 6906 11581 6936
rect 12013 6906 12083 6936
rect 12515 6906 12585 6936
rect 13017 6906 13087 6936
rect 13519 6906 13589 6936
rect 14021 6906 14091 6936
rect 14523 6906 14593 6936
rect 15025 6906 15095 6936
rect 15527 6906 15597 6936
rect 16029 6906 16099 6936
rect -2157 6645 -2143 6677
rect -1968 6645 -1950 6677
rect 17694 6677 17901 7085
rect -2157 6237 -1950 6645
rect 969 6618 1039 6648
rect 1471 6618 1541 6648
rect 1973 6618 2043 6648
rect 2475 6618 2545 6648
rect 2977 6618 3047 6648
rect 3479 6618 3549 6648
rect 3981 6618 4051 6648
rect 4483 6618 4553 6648
rect 4985 6618 5055 6648
rect 5487 6618 5557 6648
rect 5989 6618 6059 6648
rect 6491 6618 6561 6648
rect 6993 6618 7063 6648
rect 7495 6618 7565 6648
rect 7997 6618 8067 6648
rect 8499 6618 8569 6648
rect 9001 6618 9071 6648
rect 9503 6618 9573 6648
rect 10005 6618 10075 6648
rect 10507 6618 10577 6648
rect 11009 6618 11079 6648
rect 11511 6618 11581 6648
rect 12013 6618 12083 6648
rect 12515 6618 12585 6648
rect 13017 6618 13087 6648
rect 13519 6618 13589 6648
rect 14021 6618 14091 6648
rect 14523 6618 14593 6648
rect 15025 6618 15095 6648
rect 15527 6618 15597 6648
rect 16029 6618 16099 6648
rect 17694 6645 17712 6677
rect 17887 6645 17901 6677
rect 594 6491 624 6561
rect 882 6491 912 6561
rect 1096 6491 1126 6561
rect 1384 6491 1414 6561
rect 1598 6491 1628 6561
rect 1886 6491 1916 6561
rect 2100 6491 2130 6561
rect 2388 6491 2418 6561
rect 2602 6491 2632 6561
rect 2890 6491 2920 6561
rect 3104 6491 3134 6561
rect 3392 6491 3422 6561
rect 3606 6491 3636 6561
rect 3894 6491 3924 6561
rect 4108 6491 4138 6561
rect 4396 6491 4426 6561
rect 4610 6491 4640 6561
rect 4898 6491 4928 6561
rect 5112 6491 5142 6561
rect 5400 6491 5430 6561
rect 5614 6491 5644 6561
rect 5902 6491 5932 6561
rect 6116 6491 6146 6561
rect 6404 6491 6434 6561
rect 6618 6491 6648 6561
rect 6906 6491 6936 6561
rect 7120 6491 7150 6561
rect 7408 6491 7438 6561
rect 7622 6491 7652 6561
rect 7910 6491 7940 6561
rect 8124 6491 8154 6561
rect 8412 6491 8442 6561
rect 8626 6491 8656 6561
rect 8914 6491 8944 6561
rect 9128 6491 9158 6561
rect 9416 6491 9446 6561
rect 9630 6491 9660 6561
rect 9918 6491 9948 6561
rect 10132 6491 10162 6561
rect 10420 6491 10450 6561
rect 10634 6491 10664 6561
rect 10922 6491 10952 6561
rect 11136 6491 11166 6561
rect 11424 6491 11454 6561
rect 11638 6491 11668 6561
rect 11926 6491 11956 6561
rect 12140 6491 12170 6561
rect 12428 6491 12458 6561
rect 12642 6491 12672 6561
rect 12930 6491 12960 6561
rect 13144 6491 13174 6561
rect 13432 6491 13462 6561
rect 13646 6491 13676 6561
rect 13934 6491 13964 6561
rect 14148 6491 14178 6561
rect 14436 6491 14466 6561
rect 14650 6491 14680 6561
rect 14938 6491 14968 6561
rect 15152 6491 15182 6561
rect 15440 6491 15470 6561
rect 15654 6491 15684 6561
rect 15942 6491 15972 6561
rect 16156 6491 16186 6561
rect 16444 6491 16474 6561
rect 969 6404 1039 6434
rect 1471 6404 1541 6434
rect 1973 6404 2043 6434
rect 2475 6404 2545 6434
rect 2977 6404 3047 6434
rect 3479 6404 3549 6434
rect 3981 6404 4051 6434
rect 4483 6404 4553 6434
rect 4985 6404 5055 6434
rect 5487 6404 5557 6434
rect 5989 6404 6059 6434
rect 6491 6404 6561 6434
rect 6993 6404 7063 6434
rect 7495 6404 7565 6434
rect 7997 6404 8067 6434
rect 8499 6404 8569 6434
rect 9001 6404 9071 6434
rect 9503 6404 9573 6434
rect 10005 6404 10075 6434
rect 10507 6404 10577 6434
rect 11009 6404 11079 6434
rect 11511 6404 11581 6434
rect 12013 6404 12083 6434
rect 12515 6404 12585 6434
rect 13017 6404 13087 6434
rect 13519 6404 13589 6434
rect 14021 6404 14091 6434
rect 14523 6404 14593 6434
rect 15025 6404 15095 6434
rect 15527 6404 15597 6434
rect 16029 6404 16099 6434
rect -2157 6205 -2143 6237
rect -1968 6205 -1950 6237
rect -2157 5797 -1950 6205
rect 17694 6237 17901 6645
rect 17694 6205 17712 6237
rect 17887 6205 17901 6237
rect 969 6116 1039 6146
rect 1471 6116 1541 6146
rect 1973 6116 2043 6146
rect 2475 6116 2545 6146
rect 2977 6116 3047 6146
rect 3479 6116 3549 6146
rect 3981 6116 4051 6146
rect 4483 6116 4553 6146
rect 4985 6116 5055 6146
rect 5487 6116 5557 6146
rect 5989 6116 6059 6146
rect 6491 6116 6561 6146
rect 6993 6116 7063 6146
rect 7495 6116 7565 6146
rect 7997 6116 8067 6146
rect 8499 6116 8569 6146
rect 9001 6116 9071 6146
rect 9503 6116 9573 6146
rect 10005 6116 10075 6146
rect 10507 6116 10577 6146
rect 11009 6116 11079 6146
rect 11511 6116 11581 6146
rect 12013 6116 12083 6146
rect 12515 6116 12585 6146
rect 13017 6116 13087 6146
rect 13519 6116 13589 6146
rect 14021 6116 14091 6146
rect 14523 6116 14593 6146
rect 15025 6116 15095 6146
rect 15527 6116 15597 6146
rect 16029 6116 16099 6146
rect 594 5989 624 6059
rect 882 5989 912 6059
rect 1096 5989 1126 6059
rect 1384 5989 1414 6059
rect 1598 5989 1628 6059
rect 1886 5989 1916 6059
rect 2100 5989 2130 6059
rect 2388 5989 2418 6059
rect 2602 5989 2632 6059
rect 2890 5989 2920 6059
rect 3104 5989 3134 6059
rect 3392 5989 3422 6059
rect 3606 5989 3636 6059
rect 3894 5989 3924 6059
rect 4108 5989 4138 6059
rect 4396 5989 4426 6059
rect 4610 5989 4640 6059
rect 4898 5989 4928 6059
rect 5112 5989 5142 6059
rect 5400 5989 5430 6059
rect 5614 5989 5644 6059
rect 5902 5989 5932 6059
rect 6116 5989 6146 6059
rect 6404 5989 6434 6059
rect 6618 5989 6648 6059
rect 6906 5989 6936 6059
rect 7120 5989 7150 6059
rect 7408 5989 7438 6059
rect 7622 5989 7652 6059
rect 7910 5989 7940 6059
rect 8124 5989 8154 6059
rect 8412 5989 8442 6059
rect 8626 5989 8656 6059
rect 8914 5989 8944 6059
rect 9128 5989 9158 6059
rect 9416 5989 9446 6059
rect 9630 5989 9660 6059
rect 9918 5989 9948 6059
rect 10132 5989 10162 6059
rect 10420 5989 10450 6059
rect 10634 5989 10664 6059
rect 10922 5989 10952 6059
rect 11136 5989 11166 6059
rect 11424 5989 11454 6059
rect 11638 5989 11668 6059
rect 11926 5989 11956 6059
rect 12140 5989 12170 6059
rect 12428 5989 12458 6059
rect 12642 5989 12672 6059
rect 12930 5989 12960 6059
rect 13144 5989 13174 6059
rect 13432 5989 13462 6059
rect 13646 5989 13676 6059
rect 13934 5989 13964 6059
rect 14148 5989 14178 6059
rect 14436 5989 14466 6059
rect 14650 5989 14680 6059
rect 14938 5989 14968 6059
rect 15152 5989 15182 6059
rect 15440 5989 15470 6059
rect 15654 5989 15684 6059
rect 15942 5989 15972 6059
rect 16156 5989 16186 6059
rect 16444 5989 16474 6059
rect 969 5902 1039 5932
rect 1471 5902 1541 5932
rect 1973 5902 2043 5932
rect 2475 5902 2545 5932
rect 2977 5902 3047 5932
rect 3479 5902 3549 5932
rect 3981 5902 4051 5932
rect 4483 5902 4553 5932
rect 4985 5902 5055 5932
rect 5487 5902 5557 5932
rect 5989 5902 6059 5932
rect 6491 5902 6561 5932
rect 6993 5902 7063 5932
rect 7495 5902 7565 5932
rect 7997 5902 8067 5932
rect 8499 5902 8569 5932
rect 9001 5902 9071 5932
rect 9503 5902 9573 5932
rect 10005 5902 10075 5932
rect 10507 5902 10577 5932
rect 11009 5902 11079 5932
rect 11511 5902 11581 5932
rect 12013 5902 12083 5932
rect 12515 5902 12585 5932
rect 13017 5902 13087 5932
rect 13519 5902 13589 5932
rect 14021 5902 14091 5932
rect 14523 5902 14593 5932
rect 15025 5902 15095 5932
rect 15527 5902 15597 5932
rect 16029 5902 16099 5932
rect -2157 5765 -2143 5797
rect -1968 5765 -1950 5797
rect -2157 5357 -1950 5765
rect 17694 5797 17901 6205
rect 17694 5765 17712 5797
rect 17887 5765 17901 5797
rect 969 5614 1039 5644
rect 1471 5614 1541 5644
rect 1973 5614 2043 5644
rect 2475 5614 2545 5644
rect 2977 5614 3047 5644
rect 3479 5614 3549 5644
rect 3981 5614 4051 5644
rect 4483 5614 4553 5644
rect 4985 5614 5055 5644
rect 5487 5614 5557 5644
rect 5989 5614 6059 5644
rect 6491 5614 6561 5644
rect 6993 5614 7063 5644
rect 7495 5614 7565 5644
rect 7997 5614 8067 5644
rect 8499 5614 8569 5644
rect 9001 5614 9071 5644
rect 9503 5614 9573 5644
rect 10005 5614 10075 5644
rect 10507 5614 10577 5644
rect 11009 5614 11079 5644
rect 11511 5614 11581 5644
rect 12013 5614 12083 5644
rect 12515 5614 12585 5644
rect 13017 5614 13087 5644
rect 13519 5614 13589 5644
rect 14021 5614 14091 5644
rect 14523 5614 14593 5644
rect 15025 5614 15095 5644
rect 15527 5614 15597 5644
rect 16029 5614 16099 5644
rect 594 5487 624 5557
rect 882 5487 912 5557
rect 1096 5487 1126 5557
rect 1384 5487 1414 5557
rect 1598 5487 1628 5557
rect 1886 5487 1916 5557
rect 2100 5487 2130 5557
rect 2388 5487 2418 5557
rect 2602 5487 2632 5557
rect 2890 5487 2920 5557
rect 3104 5487 3134 5557
rect 3392 5487 3422 5557
rect 3606 5487 3636 5557
rect 3894 5487 3924 5557
rect 4108 5487 4138 5557
rect 4396 5487 4426 5557
rect 4610 5487 4640 5557
rect 4898 5487 4928 5557
rect 5112 5487 5142 5557
rect 5400 5487 5430 5557
rect 5614 5487 5644 5557
rect 5902 5487 5932 5557
rect 6116 5487 6146 5557
rect 6404 5487 6434 5557
rect 6618 5487 6648 5557
rect 6906 5487 6936 5557
rect 7120 5487 7150 5557
rect 7408 5487 7438 5557
rect 7622 5487 7652 5557
rect 7910 5487 7940 5557
rect 8124 5487 8154 5557
rect 8412 5487 8442 5557
rect 8626 5487 8656 5557
rect 8914 5487 8944 5557
rect 9128 5487 9158 5557
rect 9416 5487 9446 5557
rect 9630 5487 9660 5557
rect 9918 5487 9948 5557
rect 10132 5487 10162 5557
rect 10420 5487 10450 5557
rect 10634 5487 10664 5557
rect 10922 5487 10952 5557
rect 11136 5487 11166 5557
rect 11424 5487 11454 5557
rect 11638 5487 11668 5557
rect 11926 5487 11956 5557
rect 12140 5487 12170 5557
rect 12428 5487 12458 5557
rect 12642 5487 12672 5557
rect 12930 5487 12960 5557
rect 13144 5487 13174 5557
rect 13432 5487 13462 5557
rect 13646 5487 13676 5557
rect 13934 5487 13964 5557
rect 14148 5487 14178 5557
rect 14436 5487 14466 5557
rect 14650 5487 14680 5557
rect 14938 5487 14968 5557
rect 15152 5487 15182 5557
rect 15440 5487 15470 5557
rect 15654 5487 15684 5557
rect 15942 5487 15972 5557
rect 16156 5487 16186 5557
rect 16444 5487 16474 5557
rect 969 5400 1039 5430
rect 1471 5400 1541 5430
rect 1973 5400 2043 5430
rect 2475 5400 2545 5430
rect 2977 5400 3047 5430
rect 3479 5400 3549 5430
rect 3981 5400 4051 5430
rect 4483 5400 4553 5430
rect 4985 5400 5055 5430
rect 5487 5400 5557 5430
rect 5989 5400 6059 5430
rect 6491 5400 6561 5430
rect 6993 5400 7063 5430
rect 7495 5400 7565 5430
rect 7997 5400 8067 5430
rect 8499 5400 8569 5430
rect 9001 5400 9071 5430
rect 9503 5400 9573 5430
rect 10005 5400 10075 5430
rect 10507 5400 10577 5430
rect 11009 5400 11079 5430
rect 11511 5400 11581 5430
rect 12013 5400 12083 5430
rect 12515 5400 12585 5430
rect 13017 5400 13087 5430
rect 13519 5400 13589 5430
rect 14021 5400 14091 5430
rect 14523 5400 14593 5430
rect 15025 5400 15095 5430
rect 15527 5400 15597 5430
rect 16029 5400 16099 5430
rect -2157 5325 -2143 5357
rect -1968 5325 -1950 5357
rect -2157 4917 -1950 5325
rect 17694 5357 17901 5765
rect 17694 5325 17712 5357
rect 17887 5325 17901 5357
rect 969 5112 1039 5142
rect 1471 5112 1541 5142
rect 1973 5112 2043 5142
rect 2475 5112 2545 5142
rect 2977 5112 3047 5142
rect 3479 5112 3549 5142
rect 3981 5112 4051 5142
rect 4483 5112 4553 5142
rect 4985 5112 5055 5142
rect 5487 5112 5557 5142
rect 5989 5112 6059 5142
rect 6491 5112 6561 5142
rect 6993 5112 7063 5142
rect 7495 5112 7565 5142
rect 7997 5112 8067 5142
rect 8499 5112 8569 5142
rect 9001 5112 9071 5142
rect 9503 5112 9573 5142
rect 10005 5112 10075 5142
rect 10507 5112 10577 5142
rect 11009 5112 11079 5142
rect 11511 5112 11581 5142
rect 12013 5112 12083 5142
rect 12515 5112 12585 5142
rect 13017 5112 13087 5142
rect 13519 5112 13589 5142
rect 14021 5112 14091 5142
rect 14523 5112 14593 5142
rect 15025 5112 15095 5142
rect 15527 5112 15597 5142
rect 16029 5112 16099 5142
rect 594 4985 624 5055
rect 882 4985 912 5055
rect 1096 4985 1126 5055
rect 1384 4985 1414 5055
rect 1598 4985 1628 5055
rect 1886 4985 1916 5055
rect 2100 4985 2130 5055
rect 2388 4985 2418 5055
rect 2602 4985 2632 5055
rect 2890 4985 2920 5055
rect 3104 4985 3134 5055
rect 3392 4985 3422 5055
rect 3606 4985 3636 5055
rect 3894 4985 3924 5055
rect 4108 4985 4138 5055
rect 4396 4985 4426 5055
rect 4610 4985 4640 5055
rect 4898 4985 4928 5055
rect 5112 4985 5142 5055
rect 5400 4985 5430 5055
rect 5614 4985 5644 5055
rect 5902 4985 5932 5055
rect 6116 4985 6146 5055
rect 6404 4985 6434 5055
rect 6618 4985 6648 5055
rect 6906 4985 6936 5055
rect 7120 4985 7150 5055
rect 7408 4985 7438 5055
rect 7622 4985 7652 5055
rect 7910 4985 7940 5055
rect 8124 4985 8154 5055
rect 8412 4985 8442 5055
rect 8626 4985 8656 5055
rect 8914 4985 8944 5055
rect 9128 4985 9158 5055
rect 9416 4985 9446 5055
rect 9630 4985 9660 5055
rect 9918 4985 9948 5055
rect 10132 4985 10162 5055
rect 10420 4985 10450 5055
rect 10634 4985 10664 5055
rect 10922 4985 10952 5055
rect 11136 4985 11166 5055
rect 11424 4985 11454 5055
rect 11638 4985 11668 5055
rect 11926 4985 11956 5055
rect 12140 4985 12170 5055
rect 12428 4985 12458 5055
rect 12642 4985 12672 5055
rect 12930 4985 12960 5055
rect 13144 4985 13174 5055
rect 13432 4985 13462 5055
rect 13646 4985 13676 5055
rect 13934 4985 13964 5055
rect 14148 4985 14178 5055
rect 14436 4985 14466 5055
rect 14650 4985 14680 5055
rect 14938 4985 14968 5055
rect 15152 4985 15182 5055
rect 15440 4985 15470 5055
rect 15654 4985 15684 5055
rect 15942 4985 15972 5055
rect 16156 4985 16186 5055
rect 16444 4985 16474 5055
rect -2157 4885 -2143 4917
rect -1968 4885 -1950 4917
rect 969 4898 1039 4928
rect 1471 4898 1541 4928
rect 1973 4898 2043 4928
rect 2475 4898 2545 4928
rect 2977 4898 3047 4928
rect 3479 4898 3549 4928
rect 3981 4898 4051 4928
rect 4483 4898 4553 4928
rect 4985 4898 5055 4928
rect 5487 4898 5557 4928
rect 5989 4898 6059 4928
rect 6491 4898 6561 4928
rect 6993 4898 7063 4928
rect 7495 4898 7565 4928
rect 7997 4898 8067 4928
rect 8499 4898 8569 4928
rect 9001 4898 9071 4928
rect 9503 4898 9573 4928
rect 10005 4898 10075 4928
rect 10507 4898 10577 4928
rect 11009 4898 11079 4928
rect 11511 4898 11581 4928
rect 12013 4898 12083 4928
rect 12515 4898 12585 4928
rect 13017 4898 13087 4928
rect 13519 4898 13589 4928
rect 14021 4898 14091 4928
rect 14523 4898 14593 4928
rect 15025 4898 15095 4928
rect 15527 4898 15597 4928
rect 16029 4898 16099 4928
rect 17694 4917 17901 5325
rect -2157 4477 -1950 4885
rect 17694 4885 17712 4917
rect 17887 4885 17901 4917
rect 969 4610 1039 4640
rect 1471 4610 1541 4640
rect 1973 4610 2043 4640
rect 2475 4610 2545 4640
rect 2977 4610 3047 4640
rect 3479 4610 3549 4640
rect 3981 4610 4051 4640
rect 4483 4610 4553 4640
rect 4985 4610 5055 4640
rect 5487 4610 5557 4640
rect 5989 4610 6059 4640
rect 6491 4610 6561 4640
rect 6993 4610 7063 4640
rect 7495 4610 7565 4640
rect 7997 4610 8067 4640
rect 8499 4610 8569 4640
rect 9001 4610 9071 4640
rect 9503 4610 9573 4640
rect 10005 4610 10075 4640
rect 10507 4610 10577 4640
rect 11009 4610 11079 4640
rect 11511 4610 11581 4640
rect 12013 4610 12083 4640
rect 12515 4610 12585 4640
rect 13017 4610 13087 4640
rect 13519 4610 13589 4640
rect 14021 4610 14091 4640
rect 14523 4610 14593 4640
rect 15025 4610 15095 4640
rect 15527 4610 15597 4640
rect 16029 4610 16099 4640
rect 594 4483 624 4553
rect 882 4483 912 4553
rect 1096 4483 1126 4553
rect 1384 4483 1414 4553
rect 1598 4483 1628 4553
rect 1886 4483 1916 4553
rect 2100 4483 2130 4553
rect 2388 4483 2418 4553
rect 2602 4483 2632 4553
rect 2890 4483 2920 4553
rect 3104 4483 3134 4553
rect 3392 4483 3422 4553
rect 3606 4483 3636 4553
rect 3894 4483 3924 4553
rect 4108 4483 4138 4553
rect 4396 4483 4426 4553
rect 4610 4483 4640 4553
rect 4898 4483 4928 4553
rect 5112 4483 5142 4553
rect 5400 4483 5430 4553
rect 5614 4483 5644 4553
rect 5902 4483 5932 4553
rect 6116 4483 6146 4553
rect 6404 4483 6434 4553
rect 6618 4483 6648 4553
rect 6906 4483 6936 4553
rect 7120 4483 7150 4553
rect 7408 4483 7438 4553
rect 7622 4483 7652 4553
rect 7910 4483 7940 4553
rect 8124 4483 8154 4553
rect 8412 4483 8442 4553
rect 8626 4483 8656 4553
rect 8914 4483 8944 4553
rect 9128 4483 9158 4553
rect 9416 4483 9446 4553
rect 9630 4483 9660 4553
rect 9918 4483 9948 4553
rect 10132 4483 10162 4553
rect 10420 4483 10450 4553
rect 10634 4483 10664 4553
rect 10922 4483 10952 4553
rect 11136 4483 11166 4553
rect 11424 4483 11454 4553
rect 11638 4483 11668 4553
rect 11926 4483 11956 4553
rect 12140 4483 12170 4553
rect 12428 4483 12458 4553
rect 12642 4483 12672 4553
rect 12930 4483 12960 4553
rect 13144 4483 13174 4553
rect 13432 4483 13462 4553
rect 13646 4483 13676 4553
rect 13934 4483 13964 4553
rect 14148 4483 14178 4553
rect 14436 4483 14466 4553
rect 14650 4483 14680 4553
rect 14938 4483 14968 4553
rect 15152 4483 15182 4553
rect 15440 4483 15470 4553
rect 15654 4483 15684 4553
rect 15942 4483 15972 4553
rect 16156 4483 16186 4553
rect 16444 4483 16474 4553
rect -2157 4445 -2143 4477
rect -1968 4445 -1950 4477
rect -2157 4037 -1950 4445
rect 17694 4477 17901 4885
rect 17694 4445 17712 4477
rect 17887 4445 17901 4477
rect 969 4396 1039 4426
rect 1471 4396 1541 4426
rect 1973 4396 2043 4426
rect 2475 4396 2545 4426
rect 2977 4396 3047 4426
rect 3479 4396 3549 4426
rect 3981 4396 4051 4426
rect 4483 4396 4553 4426
rect 4985 4396 5055 4426
rect 5487 4396 5557 4426
rect 5989 4396 6059 4426
rect 6491 4396 6561 4426
rect 6993 4396 7063 4426
rect 7495 4396 7565 4426
rect 7997 4396 8067 4426
rect 8499 4396 8569 4426
rect 9001 4396 9071 4426
rect 9503 4396 9573 4426
rect 10005 4396 10075 4426
rect 10507 4396 10577 4426
rect 11009 4396 11079 4426
rect 11511 4396 11581 4426
rect 12013 4396 12083 4426
rect 12515 4396 12585 4426
rect 13017 4396 13087 4426
rect 13519 4396 13589 4426
rect 14021 4396 14091 4426
rect 14523 4396 14593 4426
rect 15025 4396 15095 4426
rect 15527 4396 15597 4426
rect 16029 4396 16099 4426
rect 969 4108 1039 4138
rect 1471 4108 1541 4138
rect 1973 4108 2043 4138
rect 2475 4108 2545 4138
rect 2977 4108 3047 4138
rect 3479 4108 3549 4138
rect 3981 4108 4051 4138
rect 4483 4108 4553 4138
rect 4985 4108 5055 4138
rect 5487 4108 5557 4138
rect 5989 4108 6059 4138
rect 6491 4108 6561 4138
rect 6993 4108 7063 4138
rect 7495 4108 7565 4138
rect 7997 4108 8067 4138
rect 8499 4108 8569 4138
rect 9001 4108 9071 4138
rect 9503 4108 9573 4138
rect 10005 4108 10075 4138
rect 10507 4108 10577 4138
rect 11009 4108 11079 4138
rect 11511 4108 11581 4138
rect 12013 4108 12083 4138
rect 12515 4108 12585 4138
rect 13017 4108 13087 4138
rect 13519 4108 13589 4138
rect 14021 4108 14091 4138
rect 14523 4108 14593 4138
rect 15025 4108 15095 4138
rect 15527 4108 15597 4138
rect 16029 4108 16099 4138
rect -2157 4005 -2143 4037
rect -1968 4005 -1950 4037
rect -2157 3597 -1950 4005
rect 594 3981 624 4051
rect 882 3981 912 4051
rect 1096 3981 1126 4051
rect 1384 3981 1414 4051
rect 1598 3981 1628 4051
rect 1886 3981 1916 4051
rect 2100 3981 2130 4051
rect 2388 3981 2418 4051
rect 2602 3981 2632 4051
rect 2890 3981 2920 4051
rect 3104 3981 3134 4051
rect 3392 3981 3422 4051
rect 3606 3981 3636 4051
rect 3894 3981 3924 4051
rect 4108 3981 4138 4051
rect 4396 3981 4426 4051
rect 4610 3981 4640 4051
rect 4898 3981 4928 4051
rect 5112 3981 5142 4051
rect 5400 3981 5430 4051
rect 5614 3981 5644 4051
rect 5902 3981 5932 4051
rect 6116 3981 6146 4051
rect 6404 3981 6434 4051
rect 6618 3981 6648 4051
rect 6906 3981 6936 4051
rect 7120 3981 7150 4051
rect 7408 3981 7438 4051
rect 7622 3981 7652 4051
rect 7910 3981 7940 4051
rect 8124 3981 8154 4051
rect 8412 3981 8442 4051
rect 8626 3981 8656 4051
rect 8914 3981 8944 4051
rect 9128 3981 9158 4051
rect 9416 3981 9446 4051
rect 9630 3981 9660 4051
rect 9918 3981 9948 4051
rect 10132 3981 10162 4051
rect 10420 3981 10450 4051
rect 10634 3981 10664 4051
rect 10922 3981 10952 4051
rect 11136 3981 11166 4051
rect 11424 3981 11454 4051
rect 11638 3981 11668 4051
rect 11926 3981 11956 4051
rect 12140 3981 12170 4051
rect 12428 3981 12458 4051
rect 12642 3981 12672 4051
rect 12930 3981 12960 4051
rect 13144 3981 13174 4051
rect 13432 3981 13462 4051
rect 13646 3981 13676 4051
rect 13934 3981 13964 4051
rect 14148 3981 14178 4051
rect 14436 3981 14466 4051
rect 14650 3981 14680 4051
rect 14938 3981 14968 4051
rect 15152 3981 15182 4051
rect 15440 3981 15470 4051
rect 15654 3981 15684 4051
rect 15942 3981 15972 4051
rect 16156 3981 16186 4051
rect 16444 3981 16474 4051
rect 17694 4037 17901 4445
rect 17694 4005 17712 4037
rect 17887 4005 17901 4037
rect 969 3894 1039 3924
rect 1471 3894 1541 3924
rect 1973 3894 2043 3924
rect 2475 3894 2545 3924
rect 2977 3894 3047 3924
rect 3479 3894 3549 3924
rect 3981 3894 4051 3924
rect 4483 3894 4553 3924
rect 4985 3894 5055 3924
rect 5487 3894 5557 3924
rect 5989 3894 6059 3924
rect 6491 3894 6561 3924
rect 6993 3894 7063 3924
rect 7495 3894 7565 3924
rect 7997 3894 8067 3924
rect 8499 3894 8569 3924
rect 9001 3894 9071 3924
rect 9503 3894 9573 3924
rect 10005 3894 10075 3924
rect 10507 3894 10577 3924
rect 11009 3894 11079 3924
rect 11511 3894 11581 3924
rect 12013 3894 12083 3924
rect 12515 3894 12585 3924
rect 13017 3894 13087 3924
rect 13519 3894 13589 3924
rect 14021 3894 14091 3924
rect 14523 3894 14593 3924
rect 15025 3894 15095 3924
rect 15527 3894 15597 3924
rect 16029 3894 16099 3924
rect 969 3606 1039 3636
rect 1471 3606 1541 3636
rect 1973 3606 2043 3636
rect 2475 3606 2545 3636
rect 2977 3606 3047 3636
rect 3479 3606 3549 3636
rect 3981 3606 4051 3636
rect 4483 3606 4553 3636
rect 4985 3606 5055 3636
rect 5487 3606 5557 3636
rect 5989 3606 6059 3636
rect 6491 3606 6561 3636
rect 6993 3606 7063 3636
rect 7495 3606 7565 3636
rect 7997 3606 8067 3636
rect 8499 3606 8569 3636
rect 9001 3606 9071 3636
rect 9503 3606 9573 3636
rect 10005 3606 10075 3636
rect 10507 3606 10577 3636
rect 11009 3606 11079 3636
rect 11511 3606 11581 3636
rect 12013 3606 12083 3636
rect 12515 3606 12585 3636
rect 13017 3606 13087 3636
rect 13519 3606 13589 3636
rect 14021 3606 14091 3636
rect 14523 3606 14593 3636
rect 15025 3606 15095 3636
rect 15527 3606 15597 3636
rect 16029 3606 16099 3636
rect -2157 3565 -2143 3597
rect -1968 3565 -1950 3597
rect -2157 3157 -1950 3565
rect 17694 3597 17901 4005
rect 17694 3565 17712 3597
rect 17887 3565 17901 3597
rect 594 3479 624 3549
rect 882 3479 912 3549
rect 1096 3479 1126 3549
rect 1384 3479 1414 3549
rect 1598 3479 1628 3549
rect 1886 3479 1916 3549
rect 2100 3479 2130 3549
rect 2388 3479 2418 3549
rect 2602 3479 2632 3549
rect 2890 3479 2920 3549
rect 3104 3479 3134 3549
rect 3392 3479 3422 3549
rect 3606 3479 3636 3549
rect 3894 3479 3924 3549
rect 4108 3479 4138 3549
rect 4396 3479 4426 3549
rect 4610 3479 4640 3549
rect 4898 3479 4928 3549
rect 5112 3479 5142 3549
rect 5400 3479 5430 3549
rect 5614 3479 5644 3549
rect 5902 3479 5932 3549
rect 6116 3479 6146 3549
rect 6404 3479 6434 3549
rect 6618 3479 6648 3549
rect 6906 3479 6936 3549
rect 7120 3479 7150 3549
rect 7408 3479 7438 3549
rect 7622 3479 7652 3549
rect 7910 3479 7940 3549
rect 8124 3479 8154 3549
rect 8412 3479 8442 3549
rect 8626 3479 8656 3549
rect 8914 3479 8944 3549
rect 9128 3479 9158 3549
rect 9416 3479 9446 3549
rect 9630 3479 9660 3549
rect 9918 3479 9948 3549
rect 10132 3479 10162 3549
rect 10420 3479 10450 3549
rect 10634 3479 10664 3549
rect 10922 3479 10952 3549
rect 11136 3479 11166 3549
rect 11424 3479 11454 3549
rect 11638 3479 11668 3549
rect 11926 3479 11956 3549
rect 12140 3479 12170 3549
rect 12428 3479 12458 3549
rect 12642 3479 12672 3549
rect 12930 3479 12960 3549
rect 13144 3479 13174 3549
rect 13432 3479 13462 3549
rect 13646 3479 13676 3549
rect 13934 3479 13964 3549
rect 14148 3479 14178 3549
rect 14436 3479 14466 3549
rect 14650 3479 14680 3549
rect 14938 3479 14968 3549
rect 15152 3479 15182 3549
rect 15440 3479 15470 3549
rect 15654 3479 15684 3549
rect 15942 3479 15972 3549
rect 16156 3479 16186 3549
rect 16444 3479 16474 3549
rect 969 3392 1039 3422
rect 1471 3392 1541 3422
rect 1973 3392 2043 3422
rect 2475 3392 2545 3422
rect 2977 3392 3047 3422
rect 3479 3392 3549 3422
rect 3981 3392 4051 3422
rect 4483 3392 4553 3422
rect 4985 3392 5055 3422
rect 5487 3392 5557 3422
rect 5989 3392 6059 3422
rect 6491 3392 6561 3422
rect 6993 3392 7063 3422
rect 7495 3392 7565 3422
rect 7997 3392 8067 3422
rect 8499 3392 8569 3422
rect 9001 3392 9071 3422
rect 9503 3392 9573 3422
rect 10005 3392 10075 3422
rect 10507 3392 10577 3422
rect 11009 3392 11079 3422
rect 11511 3392 11581 3422
rect 12013 3392 12083 3422
rect 12515 3392 12585 3422
rect 13017 3392 13087 3422
rect 13519 3392 13589 3422
rect 14021 3392 14091 3422
rect 14523 3392 14593 3422
rect 15025 3392 15095 3422
rect 15527 3392 15597 3422
rect 16029 3392 16099 3422
rect -2157 3125 -2143 3157
rect -1968 3125 -1950 3157
rect 17694 3157 17901 3565
rect -2157 2717 -1950 3125
rect 969 3104 1039 3134
rect 1471 3104 1541 3134
rect 1973 3104 2043 3134
rect 2475 3104 2545 3134
rect 2977 3104 3047 3134
rect 3479 3104 3549 3134
rect 3981 3104 4051 3134
rect 4483 3104 4553 3134
rect 4985 3104 5055 3134
rect 5487 3104 5557 3134
rect 5989 3104 6059 3134
rect 6491 3104 6561 3134
rect 6993 3104 7063 3134
rect 7495 3104 7565 3134
rect 7997 3104 8067 3134
rect 8499 3104 8569 3134
rect 9001 3104 9071 3134
rect 9503 3104 9573 3134
rect 10005 3104 10075 3134
rect 10507 3104 10577 3134
rect 11009 3104 11079 3134
rect 11511 3104 11581 3134
rect 12013 3104 12083 3134
rect 12515 3104 12585 3134
rect 13017 3104 13087 3134
rect 13519 3104 13589 3134
rect 14021 3104 14091 3134
rect 14523 3104 14593 3134
rect 15025 3104 15095 3134
rect 15527 3104 15597 3134
rect 16029 3104 16099 3134
rect 17694 3125 17712 3157
rect 17887 3125 17901 3157
rect 594 2977 624 3047
rect 882 2977 912 3047
rect 1096 2977 1126 3047
rect 1384 2977 1414 3047
rect 1598 2977 1628 3047
rect 1886 2977 1916 3047
rect 2100 2977 2130 3047
rect 2388 2977 2418 3047
rect 2602 2977 2632 3047
rect 2890 2977 2920 3047
rect 3104 2977 3134 3047
rect 3392 2977 3422 3047
rect 3606 2977 3636 3047
rect 3894 2977 3924 3047
rect 4108 2977 4138 3047
rect 4396 2977 4426 3047
rect 4610 2977 4640 3047
rect 4898 2977 4928 3047
rect 5112 2977 5142 3047
rect 5400 2977 5430 3047
rect 5614 2977 5644 3047
rect 5902 2977 5932 3047
rect 6116 2977 6146 3047
rect 6404 2977 6434 3047
rect 6618 2977 6648 3047
rect 6906 2977 6936 3047
rect 7120 2977 7150 3047
rect 7408 2977 7438 3047
rect 7622 2977 7652 3047
rect 7910 2977 7940 3047
rect 8124 2977 8154 3047
rect 8412 2977 8442 3047
rect 8626 2977 8656 3047
rect 8914 2977 8944 3047
rect 9128 2977 9158 3047
rect 9416 2977 9446 3047
rect 9630 2977 9660 3047
rect 9918 2977 9948 3047
rect 10132 2977 10162 3047
rect 10420 2977 10450 3047
rect 10634 2977 10664 3047
rect 10922 2977 10952 3047
rect 11136 2977 11166 3047
rect 11424 2977 11454 3047
rect 11638 2977 11668 3047
rect 11926 2977 11956 3047
rect 12140 2977 12170 3047
rect 12428 2977 12458 3047
rect 12642 2977 12672 3047
rect 12930 2977 12960 3047
rect 13144 2977 13174 3047
rect 13432 2977 13462 3047
rect 13646 2977 13676 3047
rect 13934 2977 13964 3047
rect 14148 2977 14178 3047
rect 14436 2977 14466 3047
rect 14650 2977 14680 3047
rect 14938 2977 14968 3047
rect 15152 2977 15182 3047
rect 15440 2977 15470 3047
rect 15654 2977 15684 3047
rect 15942 2977 15972 3047
rect 16156 2977 16186 3047
rect 16444 2977 16474 3047
rect 969 2890 1039 2920
rect 1471 2890 1541 2920
rect 1973 2890 2043 2920
rect 2475 2890 2545 2920
rect 2977 2890 3047 2920
rect 3479 2890 3549 2920
rect 3981 2890 4051 2920
rect 4483 2890 4553 2920
rect 4985 2890 5055 2920
rect 5487 2890 5557 2920
rect 5989 2890 6059 2920
rect 6491 2890 6561 2920
rect 6993 2890 7063 2920
rect 7495 2890 7565 2920
rect 7997 2890 8067 2920
rect 8499 2890 8569 2920
rect 9001 2890 9071 2920
rect 9503 2890 9573 2920
rect 10005 2890 10075 2920
rect 10507 2890 10577 2920
rect 11009 2890 11079 2920
rect 11511 2890 11581 2920
rect 12013 2890 12083 2920
rect 12515 2890 12585 2920
rect 13017 2890 13087 2920
rect 13519 2890 13589 2920
rect 14021 2890 14091 2920
rect 14523 2890 14593 2920
rect 15025 2890 15095 2920
rect 15527 2890 15597 2920
rect 16029 2890 16099 2920
rect -2157 2685 -2143 2717
rect -1968 2685 -1950 2717
rect -2157 2277 -1950 2685
rect 17694 2717 17901 3125
rect 17694 2685 17712 2717
rect 17887 2685 17901 2717
rect 969 2602 1039 2632
rect 1471 2602 1541 2632
rect 1973 2602 2043 2632
rect 2475 2602 2545 2632
rect 2977 2602 3047 2632
rect 3479 2602 3549 2632
rect 3981 2602 4051 2632
rect 4483 2602 4553 2632
rect 4985 2602 5055 2632
rect 5487 2602 5557 2632
rect 5989 2602 6059 2632
rect 6491 2602 6561 2632
rect 6993 2602 7063 2632
rect 7495 2602 7565 2632
rect 7997 2602 8067 2632
rect 8499 2602 8569 2632
rect 9001 2602 9071 2632
rect 9503 2602 9573 2632
rect 10005 2602 10075 2632
rect 10507 2602 10577 2632
rect 11009 2602 11079 2632
rect 11511 2602 11581 2632
rect 12013 2602 12083 2632
rect 12515 2602 12585 2632
rect 13017 2602 13087 2632
rect 13519 2602 13589 2632
rect 14021 2602 14091 2632
rect 14523 2602 14593 2632
rect 15025 2602 15095 2632
rect 15527 2602 15597 2632
rect 16029 2602 16099 2632
rect 594 2475 624 2545
rect 882 2475 912 2545
rect 1096 2475 1126 2545
rect 1384 2475 1414 2545
rect 1598 2475 1628 2545
rect 1886 2475 1916 2545
rect 2100 2475 2130 2545
rect 2388 2475 2418 2545
rect 2602 2475 2632 2545
rect 2890 2475 2920 2545
rect 3104 2475 3134 2545
rect 3392 2475 3422 2545
rect 3606 2475 3636 2545
rect 3894 2475 3924 2545
rect 4108 2475 4138 2545
rect 4396 2475 4426 2545
rect 4610 2475 4640 2545
rect 4898 2475 4928 2545
rect 5112 2475 5142 2545
rect 5400 2475 5430 2545
rect 5614 2475 5644 2545
rect 5902 2475 5932 2545
rect 6116 2475 6146 2545
rect 6404 2475 6434 2545
rect 6618 2475 6648 2545
rect 6906 2475 6936 2545
rect 7120 2475 7150 2545
rect 7408 2475 7438 2545
rect 7622 2475 7652 2545
rect 7910 2475 7940 2545
rect 8124 2475 8154 2545
rect 8412 2475 8442 2545
rect 8626 2475 8656 2545
rect 8914 2475 8944 2545
rect 9128 2475 9158 2545
rect 9416 2475 9446 2545
rect 9630 2475 9660 2545
rect 9918 2475 9948 2545
rect 10132 2475 10162 2545
rect 10420 2475 10450 2545
rect 10634 2475 10664 2545
rect 10922 2475 10952 2545
rect 11136 2475 11166 2545
rect 11424 2475 11454 2545
rect 11638 2475 11668 2545
rect 11926 2475 11956 2545
rect 12140 2475 12170 2545
rect 12428 2475 12458 2545
rect 12642 2475 12672 2545
rect 12930 2475 12960 2545
rect 13144 2475 13174 2545
rect 13432 2475 13462 2545
rect 13646 2475 13676 2545
rect 13934 2475 13964 2545
rect 14148 2475 14178 2545
rect 14436 2475 14466 2545
rect 14650 2475 14680 2545
rect 14938 2475 14968 2545
rect 15152 2475 15182 2545
rect 15440 2475 15470 2545
rect 15654 2475 15684 2545
rect 15942 2475 15972 2545
rect 16156 2475 16186 2545
rect 16444 2475 16474 2545
rect 969 2388 1039 2418
rect 1471 2388 1541 2418
rect 1973 2388 2043 2418
rect 2475 2388 2545 2418
rect 2977 2388 3047 2418
rect 3479 2388 3549 2418
rect 3981 2388 4051 2418
rect 4483 2388 4553 2418
rect 4985 2388 5055 2418
rect 5487 2388 5557 2418
rect 5989 2388 6059 2418
rect 6491 2388 6561 2418
rect 6993 2388 7063 2418
rect 7495 2388 7565 2418
rect 7997 2388 8067 2418
rect 8499 2388 8569 2418
rect 9001 2388 9071 2418
rect 9503 2388 9573 2418
rect 10005 2388 10075 2418
rect 10507 2388 10577 2418
rect 11009 2388 11079 2418
rect 11511 2388 11581 2418
rect 12013 2388 12083 2418
rect 12515 2388 12585 2418
rect 13017 2388 13087 2418
rect 13519 2388 13589 2418
rect 14021 2388 14091 2418
rect 14523 2388 14593 2418
rect 15025 2388 15095 2418
rect 15527 2388 15597 2418
rect 16029 2388 16099 2418
rect -2157 2245 -2143 2277
rect -1968 2245 -1950 2277
rect -2157 1837 -1950 2245
rect 17694 2277 17901 2685
rect 17694 2245 17712 2277
rect 17887 2245 17901 2277
rect 969 2100 1039 2130
rect 1471 2100 1541 2130
rect 1973 2100 2043 2130
rect 2475 2100 2545 2130
rect 2977 2100 3047 2130
rect 3479 2100 3549 2130
rect 3981 2100 4051 2130
rect 4483 2100 4553 2130
rect 4985 2100 5055 2130
rect 5487 2100 5557 2130
rect 5989 2100 6059 2130
rect 6491 2100 6561 2130
rect 6993 2100 7063 2130
rect 7495 2100 7565 2130
rect 7997 2100 8067 2130
rect 8499 2100 8569 2130
rect 9001 2100 9071 2130
rect 9503 2100 9573 2130
rect 10005 2100 10075 2130
rect 10507 2100 10577 2130
rect 11009 2100 11079 2130
rect 11511 2100 11581 2130
rect 12013 2100 12083 2130
rect 12515 2100 12585 2130
rect 13017 2100 13087 2130
rect 13519 2100 13589 2130
rect 14021 2100 14091 2130
rect 14523 2100 14593 2130
rect 15025 2100 15095 2130
rect 15527 2100 15597 2130
rect 16029 2100 16099 2130
rect 594 1973 624 2043
rect 882 1973 912 2043
rect 1096 1973 1126 2043
rect 1384 1973 1414 2043
rect 1598 1973 1628 2043
rect 1886 1973 1916 2043
rect 2100 1973 2130 2043
rect 2388 1973 2418 2043
rect 2602 1973 2632 2043
rect 2890 1973 2920 2043
rect 3104 1973 3134 2043
rect 3392 1973 3422 2043
rect 3606 1973 3636 2043
rect 3894 1973 3924 2043
rect 4108 1973 4138 2043
rect 4396 1973 4426 2043
rect 4610 1973 4640 2043
rect 4898 1973 4928 2043
rect 5112 1973 5142 2043
rect 5400 1973 5430 2043
rect 5614 1973 5644 2043
rect 5902 1973 5932 2043
rect 6116 1973 6146 2043
rect 6404 1973 6434 2043
rect 6618 1973 6648 2043
rect 6906 1973 6936 2043
rect 7120 1973 7150 2043
rect 7408 1973 7438 2043
rect 7622 1973 7652 2043
rect 7910 1973 7940 2043
rect 8124 1973 8154 2043
rect 8412 1973 8442 2043
rect 8626 1973 8656 2043
rect 8914 1973 8944 2043
rect 9128 1973 9158 2043
rect 9416 1973 9446 2043
rect 9630 1973 9660 2043
rect 9918 1973 9948 2043
rect 10132 1973 10162 2043
rect 10420 1973 10450 2043
rect 10634 1973 10664 2043
rect 10922 1973 10952 2043
rect 11136 1973 11166 2043
rect 11424 1973 11454 2043
rect 11638 1973 11668 2043
rect 11926 1973 11956 2043
rect 12140 1973 12170 2043
rect 12428 1973 12458 2043
rect 12642 1973 12672 2043
rect 12930 1973 12960 2043
rect 13144 1973 13174 2043
rect 13432 1973 13462 2043
rect 13646 1973 13676 2043
rect 13934 1973 13964 2043
rect 14148 1973 14178 2043
rect 14436 1973 14466 2043
rect 14650 1973 14680 2043
rect 14938 1973 14968 2043
rect 15152 1973 15182 2043
rect 15440 1973 15470 2043
rect 15654 1973 15684 2043
rect 15942 1973 15972 2043
rect 16156 1973 16186 2043
rect 16444 1973 16474 2043
rect 969 1886 1039 1916
rect 1471 1886 1541 1916
rect 1973 1886 2043 1916
rect 2475 1886 2545 1916
rect 2977 1886 3047 1916
rect 3479 1886 3549 1916
rect 3981 1886 4051 1916
rect 4483 1886 4553 1916
rect 4985 1886 5055 1916
rect 5487 1886 5557 1916
rect 5989 1886 6059 1916
rect 6491 1886 6561 1916
rect 6993 1886 7063 1916
rect 7495 1886 7565 1916
rect 7997 1886 8067 1916
rect 8499 1886 8569 1916
rect 9001 1886 9071 1916
rect 9503 1886 9573 1916
rect 10005 1886 10075 1916
rect 10507 1886 10577 1916
rect 11009 1886 11079 1916
rect 11511 1886 11581 1916
rect 12013 1886 12083 1916
rect 12515 1886 12585 1916
rect 13017 1886 13087 1916
rect 13519 1886 13589 1916
rect 14021 1886 14091 1916
rect 14523 1886 14593 1916
rect 15025 1886 15095 1916
rect 15527 1886 15597 1916
rect 16029 1886 16099 1916
rect -2157 1805 -2143 1837
rect -1968 1805 -1950 1837
rect -2157 1397 -1950 1805
rect 17694 1837 17901 2245
rect 17694 1805 17712 1837
rect 17887 1805 17901 1837
rect 969 1598 1039 1628
rect 1471 1598 1541 1628
rect 1973 1598 2043 1628
rect 2475 1598 2545 1628
rect 2977 1598 3047 1628
rect 3479 1598 3549 1628
rect 3981 1598 4051 1628
rect 4483 1598 4553 1628
rect 4985 1598 5055 1628
rect 5487 1598 5557 1628
rect 5989 1598 6059 1628
rect 6491 1598 6561 1628
rect 6993 1598 7063 1628
rect 7495 1598 7565 1628
rect 7997 1598 8067 1628
rect 8499 1598 8569 1628
rect 9001 1598 9071 1628
rect 9503 1598 9573 1628
rect 10005 1598 10075 1628
rect 10507 1598 10577 1628
rect 11009 1598 11079 1628
rect 11511 1598 11581 1628
rect 12013 1598 12083 1628
rect 12515 1598 12585 1628
rect 13017 1598 13087 1628
rect 13519 1598 13589 1628
rect 14021 1598 14091 1628
rect 14523 1598 14593 1628
rect 15025 1598 15095 1628
rect 15527 1598 15597 1628
rect 16029 1598 16099 1628
rect 594 1471 624 1541
rect 882 1471 912 1541
rect 1096 1471 1126 1541
rect 1384 1471 1414 1541
rect 1598 1471 1628 1541
rect 1886 1471 1916 1541
rect 2100 1471 2130 1541
rect 2388 1471 2418 1541
rect 2602 1471 2632 1541
rect 2890 1471 2920 1541
rect 3104 1471 3134 1541
rect 3392 1471 3422 1541
rect 3606 1471 3636 1541
rect 3894 1471 3924 1541
rect 4108 1471 4138 1541
rect 4396 1471 4426 1541
rect 4610 1471 4640 1541
rect 4898 1471 4928 1541
rect 5112 1471 5142 1541
rect 5400 1471 5430 1541
rect 5614 1471 5644 1541
rect 5902 1471 5932 1541
rect 6116 1471 6146 1541
rect 6404 1471 6434 1541
rect 6618 1471 6648 1541
rect 6906 1471 6936 1541
rect 7120 1471 7150 1541
rect 7408 1471 7438 1541
rect 7622 1471 7652 1541
rect 7910 1471 7940 1541
rect 8124 1471 8154 1541
rect 8412 1471 8442 1541
rect 8626 1471 8656 1541
rect 8914 1471 8944 1541
rect 9128 1471 9158 1541
rect 9416 1471 9446 1541
rect 9630 1471 9660 1541
rect 9918 1471 9948 1541
rect 10132 1471 10162 1541
rect 10420 1471 10450 1541
rect 10634 1471 10664 1541
rect 10922 1471 10952 1541
rect 11136 1471 11166 1541
rect 11424 1471 11454 1541
rect 11638 1471 11668 1541
rect 11926 1471 11956 1541
rect 12140 1471 12170 1541
rect 12428 1471 12458 1541
rect 12642 1471 12672 1541
rect 12930 1471 12960 1541
rect 13144 1471 13174 1541
rect 13432 1471 13462 1541
rect 13646 1471 13676 1541
rect 13934 1471 13964 1541
rect 14148 1471 14178 1541
rect 14436 1471 14466 1541
rect 14650 1471 14680 1541
rect 14938 1471 14968 1541
rect 15152 1471 15182 1541
rect 15440 1471 15470 1541
rect 15654 1471 15684 1541
rect 15942 1471 15972 1541
rect 16156 1471 16186 1541
rect 16444 1471 16474 1541
rect -2157 1365 -2143 1397
rect -1968 1365 -1950 1397
rect 969 1384 1039 1414
rect 1471 1384 1541 1414
rect 1973 1384 2043 1414
rect 2475 1384 2545 1414
rect 2977 1384 3047 1414
rect 3479 1384 3549 1414
rect 3981 1384 4051 1414
rect 4483 1384 4553 1414
rect 4985 1384 5055 1414
rect 5487 1384 5557 1414
rect 5989 1384 6059 1414
rect 6491 1384 6561 1414
rect 6993 1384 7063 1414
rect 7495 1384 7565 1414
rect 7997 1384 8067 1414
rect 8499 1384 8569 1414
rect 9001 1384 9071 1414
rect 9503 1384 9573 1414
rect 10005 1384 10075 1414
rect 10507 1384 10577 1414
rect 11009 1384 11079 1414
rect 11511 1384 11581 1414
rect 12013 1384 12083 1414
rect 12515 1384 12585 1414
rect 13017 1384 13087 1414
rect 13519 1384 13589 1414
rect 14021 1384 14091 1414
rect 14523 1384 14593 1414
rect 15025 1384 15095 1414
rect 15527 1384 15597 1414
rect 16029 1384 16099 1414
rect 17694 1397 17901 1805
rect -2157 957 -1950 1365
rect 17694 1365 17712 1397
rect 17887 1365 17901 1397
rect 969 1096 1039 1126
rect 1471 1096 1541 1126
rect 1973 1096 2043 1126
rect 2475 1096 2545 1126
rect 2977 1096 3047 1126
rect 3479 1096 3549 1126
rect 3981 1096 4051 1126
rect 4483 1096 4553 1126
rect 4985 1096 5055 1126
rect 5487 1096 5557 1126
rect 5989 1096 6059 1126
rect 6491 1096 6561 1126
rect 6993 1096 7063 1126
rect 7495 1096 7565 1126
rect 7997 1096 8067 1126
rect 8499 1096 8569 1126
rect 9001 1096 9071 1126
rect 9503 1096 9573 1126
rect 10005 1096 10075 1126
rect 10507 1096 10577 1126
rect 11009 1096 11079 1126
rect 11511 1096 11581 1126
rect 12013 1096 12083 1126
rect 12515 1096 12585 1126
rect 13017 1096 13087 1126
rect 13519 1096 13589 1126
rect 14021 1096 14091 1126
rect 14523 1096 14593 1126
rect 15025 1096 15095 1126
rect 15527 1096 15597 1126
rect 16029 1096 16099 1126
rect 594 969 624 1039
rect 882 969 912 1039
rect 1096 969 1126 1039
rect 1384 969 1414 1039
rect 1598 969 1628 1039
rect 1886 969 1916 1039
rect 2100 969 2130 1039
rect 2388 969 2418 1039
rect 2602 969 2632 1039
rect 2890 969 2920 1039
rect 3104 969 3134 1039
rect 3392 969 3422 1039
rect 3606 969 3636 1039
rect 3894 969 3924 1039
rect 4108 969 4138 1039
rect 4396 969 4426 1039
rect 4610 969 4640 1039
rect 4898 969 4928 1039
rect 5112 969 5142 1039
rect 5400 969 5430 1039
rect 5614 969 5644 1039
rect 5902 969 5932 1039
rect 6116 969 6146 1039
rect 6404 969 6434 1039
rect 6618 969 6648 1039
rect 6906 969 6936 1039
rect 7120 969 7150 1039
rect 7408 969 7438 1039
rect 7622 969 7652 1039
rect 7910 969 7940 1039
rect 8124 969 8154 1039
rect 8412 969 8442 1039
rect 8626 969 8656 1039
rect 8914 969 8944 1039
rect 9128 969 9158 1039
rect 9416 969 9446 1039
rect 9630 969 9660 1039
rect 9918 969 9948 1039
rect 10132 969 10162 1039
rect 10420 969 10450 1039
rect 10634 969 10664 1039
rect 10922 969 10952 1039
rect 11136 969 11166 1039
rect 11424 969 11454 1039
rect 11638 969 11668 1039
rect 11926 969 11956 1039
rect 12140 969 12170 1039
rect 12428 969 12458 1039
rect 12642 969 12672 1039
rect 12930 969 12960 1039
rect 13144 969 13174 1039
rect 13432 969 13462 1039
rect 13646 969 13676 1039
rect 13934 969 13964 1039
rect 14148 969 14178 1039
rect 14436 969 14466 1039
rect 14650 969 14680 1039
rect 14938 969 14968 1039
rect 15152 969 15182 1039
rect 15440 969 15470 1039
rect 15654 969 15684 1039
rect 15942 969 15972 1039
rect 16156 969 16186 1039
rect 16444 969 16474 1039
rect -2157 925 -2143 957
rect -1968 925 -1950 957
rect -2157 517 -1950 925
rect 17694 957 17901 1365
rect 17694 925 17712 957
rect 17887 925 17901 957
rect 969 882 1039 912
rect 1471 882 1541 912
rect 1973 882 2043 912
rect 2475 882 2545 912
rect 2977 882 3047 912
rect 3479 882 3549 912
rect 3981 882 4051 912
rect 4483 882 4553 912
rect 4985 882 5055 912
rect 5487 882 5557 912
rect 5989 882 6059 912
rect 6491 882 6561 912
rect 6993 882 7063 912
rect 7495 882 7565 912
rect 7997 882 8067 912
rect 8499 882 8569 912
rect 9001 882 9071 912
rect 9503 882 9573 912
rect 10005 882 10075 912
rect 10507 882 10577 912
rect 11009 882 11079 912
rect 11511 882 11581 912
rect 12013 882 12083 912
rect 12515 882 12585 912
rect 13017 882 13087 912
rect 13519 882 13589 912
rect 14021 882 14091 912
rect 14523 882 14593 912
rect 15025 882 15095 912
rect 15527 882 15597 912
rect 16029 882 16099 912
rect 969 594 1039 624
rect 1471 594 1541 624
rect 1973 594 2043 624
rect 2475 594 2545 624
rect 2977 594 3047 624
rect 3479 594 3549 624
rect 3981 594 4051 624
rect 4483 594 4553 624
rect 4985 594 5055 624
rect 5487 594 5557 624
rect 5989 594 6059 624
rect 6491 594 6561 624
rect 6993 594 7063 624
rect 7495 594 7565 624
rect 7997 594 8067 624
rect 8499 594 8569 624
rect 9001 594 9071 624
rect 9503 594 9573 624
rect 10005 594 10075 624
rect 10507 594 10577 624
rect 11009 594 11079 624
rect 11511 594 11581 624
rect 12013 594 12083 624
rect 12515 594 12585 624
rect 13017 594 13087 624
rect 13519 594 13589 624
rect 14021 594 14091 624
rect 14523 594 14593 624
rect 15025 594 15095 624
rect 15527 594 15597 624
rect 16029 594 16099 624
rect -2157 485 -2143 517
rect -1968 485 -1950 517
rect -2157 77 -1950 485
rect 4610 467 4640 537
rect 4898 467 4928 537
rect 6762 467 6792 537
rect 8626 467 8656 537
rect 8770 467 8800 537
rect 12642 467 12672 537
rect 14292 467 14322 537
rect 17694 517 17901 925
rect 17694 485 17712 517
rect 17887 485 17901 517
rect 4518 380 4553 410
rect 4985 380 5020 410
rect -2157 45 -2143 77
rect -1968 45 -1950 77
rect -2157 -91 -1950 45
rect 17694 77 17901 485
rect 17694 45 17712 77
rect 17887 45 17901 77
rect -2157 -123 -2142 -91
rect -2110 -123 -2098 -91
rect -2066 -123 -2054 -91
rect -2022 -123 -2010 -91
rect -1978 -123 -1950 -91
rect -2157 -136 -1950 -123
rect -2157 -168 -2142 -136
rect -2110 -168 -2098 -136
rect -2066 -168 -2054 -136
rect -2022 -168 -2010 -136
rect -1978 -168 -1950 -136
rect -2157 -181 -1950 -168
rect -2157 -213 -2142 -181
rect -2110 -213 -2098 -181
rect -2066 -213 -2054 -181
rect -2022 -213 -2010 -181
rect -1978 -213 -1950 -181
rect -2157 -217 -1950 -213
rect -2452 -342 -2437 -310
rect -2405 -342 -2393 -310
rect -2361 -342 -2349 -310
rect -2317 -342 -2305 -310
rect -2273 -342 -2245 -310
rect -2452 -355 -2245 -342
rect -2452 -387 -2437 -355
rect -2405 -387 -2393 -355
rect -2361 -387 -2349 -355
rect -2317 -387 -2305 -355
rect -2273 -387 -2245 -355
rect -2452 -400 -2245 -387
rect -2452 -432 -2437 -400
rect -2405 -432 -2393 -400
rect -2361 -432 -2349 -400
rect -2317 -432 -2305 -400
rect -2273 -432 -2245 -400
rect -2452 -436 -2245 -432
rect 16300 -456 16330 0
rect 17694 -26 17901 45
rect 17694 -58 17722 -26
rect 17754 -58 17766 -26
rect 17798 -58 17810 -26
rect 17842 -58 17854 -26
rect 17886 -58 17901 -26
rect 17694 -71 17901 -58
rect 17694 -103 17722 -71
rect 17754 -103 17766 -71
rect 17798 -103 17810 -71
rect 17842 -103 17854 -71
rect 17886 -103 17901 -71
rect 17694 -116 17901 -103
rect 17694 -148 17722 -116
rect 17754 -148 17766 -116
rect 17798 -148 17810 -116
rect 17842 -148 17854 -116
rect 17886 -148 17901 -116
rect 17694 -152 17901 -148
rect 17989 9489 18196 9494
rect 17989 9457 18017 9489
rect 18049 9457 18061 9489
rect 18093 9457 18105 9489
rect 18137 9457 18149 9489
rect 18181 9457 18196 9489
rect 17989 9444 18196 9457
rect 17989 9412 18017 9444
rect 18049 9412 18061 9444
rect 18093 9412 18105 9444
rect 18137 9412 18149 9444
rect 18181 9412 18196 9444
rect 17989 9399 18196 9412
rect 17989 9367 18017 9399
rect 18049 9367 18061 9399
rect 18093 9367 18105 9399
rect 18137 9367 18149 9399
rect 18181 9367 18196 9399
rect 17989 -245 18196 9367
rect 17989 -277 18017 -245
rect 18049 -277 18061 -245
rect 18093 -277 18105 -245
rect 18137 -277 18149 -245
rect 18181 -277 18196 -245
rect 17989 -290 18196 -277
rect 17989 -322 18017 -290
rect 18049 -322 18061 -290
rect 18093 -322 18105 -290
rect 18137 -322 18149 -290
rect 18181 -322 18196 -290
rect 17989 -335 18196 -322
rect 17989 -367 18017 -335
rect 18049 -367 18061 -335
rect 18093 -367 18105 -335
rect 18137 -367 18149 -335
rect 18181 -367 18196 -335
rect 17989 -371 18196 -367
use adc_array_wafflecap_8_1  adc_array_wafflecap_8_1_0 ../adc_array_cap
timestamp 1662987872
transform 1 0 12550 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_2  adc_array_wafflecap_8_2_0 ../adc_array_cap
timestamp 1662983799
transform 1 0 8534 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_4  adc_array_wafflecap_8_4_0 ../adc_array_cap
timestamp 1662985026
transform 1 0 4518 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_8  adc_array_wafflecap_8_8_0 ../adc_array_cap
array 0 31 502 0 15 502
timestamp 1662984960
transform 1 0 502 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8_Drv  adc_array_wafflecap_8_Drv_0 ../adc_array_cap
array 0 0 502 0 15 502
timestamp 1663073688
transform 1 0 0 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_0 ../adc_array_cap
array 0 8 502 0 0 502
timestamp 1663073688
transform 1 0 0 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_1
array 0 6 502 0 0 502
timestamp 1663073688
transform 1 0 5020 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_2
array 0 6 502 0 0 502
timestamp 1663073688
transform 1 0 9036 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_3
array 0 5 502 0 0 502
timestamp 1663073688
transform 1 0 13052 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_4
array 0 33 502 0 0 502
timestamp 1663073688
transform 1 0 0 0 1 8534
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_5
array 0 0 502 0 15 502
timestamp 1663073688
transform 1 0 16566 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_6
timestamp 1663073688
transform 1 0 16566 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Gate  adc_array_wafflecap_8_Gate_0 ../adc_array_cap
timestamp 1663061126
transform 1 0 16064 0 1 0
box 0 0 502 502
<< labels >>
flabel locali s -1914 -457 -1895 -436 5 FreeSans 40 0 0 0 colon_n[0]
port 12 s
flabel locali s -1878 -457 -1859 -436 5 FreeSans 40 0 0 0 colon_n[1]
port 13 s
flabel locali s -1842 -457 -1823 -436 5 FreeSans 40 0 0 0 colon_n[2]
port 14 s
flabel locali s -1806 -457 -1787 -436 5 FreeSans 40 0 0 0 colon_n[3]
port 15 s
flabel locali s -1770 -457 -1751 -436 5 FreeSans 40 0 0 0 colon_n[4]
port 16 s
flabel locali s -1734 -457 -1715 -436 5 FreeSans 40 0 0 0 colon_n[5]
port 17 s
flabel locali s -1698 -457 -1679 -436 5 FreeSans 40 0 0 0 colon_n[6]
port 18 s
flabel locali s -1662 -457 -1643 -436 5 FreeSans 40 0 0 0 colon_n[7]
port 19 s
flabel locali s -1626 -457 -1607 -436 5 FreeSans 40 0 0 0 colon_n[8]
port 20 s
flabel locali s -1590 -457 -1571 -436 5 FreeSans 40 0 0 0 colon_n[9]
port 21 s
flabel locali s -1554 -457 -1535 -436 5 FreeSans 40 0 0 0 colon_n[10]
port 22 s
flabel locali s -1518 -457 -1499 -436 5 FreeSans 40 0 0 0 colon_n[11]
port 23 s
flabel locali s -1482 -457 -1463 -436 5 FreeSans 40 0 0 0 colon_n[12]
port 24 s
flabel locali s -1446 -457 -1427 -436 5 FreeSans 40 0 0 0 colon_n[13]
port 25 s
flabel locali s -1410 -457 -1391 -436 5 FreeSans 40 0 0 0 colon_n[14]
port 26 s
flabel locali s -1374 -457 -1355 -436 5 FreeSans 40 0 0 0 colon_n[15]
port 27 s
flabel locali s -1302 -457 -1283 -436 5 FreeSans 40 0 0 0 col_n[0]
port 28 s
flabel locali s -1266 -457 -1247 -436 5 FreeSans 40 0 0 0 col_n[1]
port 29 s
flabel locali s -1230 -457 -1211 -436 5 FreeSans 40 0 0 0 col_n[2]
port 30 s
flabel locali s -1194 -457 -1175 -436 5 FreeSans 40 0 0 0 col_n[3]
port 31 s
flabel locali s -1158 -457 -1139 -436 5 FreeSans 40 0 0 0 col_n[4]
port 32 s
flabel locali s -1122 -457 -1103 -436 5 FreeSans 40 0 0 0 col_n[5]
port 33 s
flabel locali s -1086 -457 -1067 -436 5 FreeSans 40 0 0 0 col_n[6]
port 34 s
flabel locali s -1050 -457 -1031 -436 5 FreeSans 40 0 0 0 col_n[7]
port 35 s
flabel locali s -1014 -457 -995 -436 5 FreeSans 40 0 0 0 col_n[8]
port 36 s
flabel locali s -978 -457 -959 -436 5 FreeSans 40 0 0 0 col_n[9]
port 37 s
flabel locali s -942 -457 -923 -436 5 FreeSans 40 0 0 0 col_n[10]
port 38 s
flabel locali s -906 -457 -887 -436 5 FreeSans 40 0 0 0 col_n[11]
port 39 s
flabel locali s -870 -457 -851 -436 5 FreeSans 40 0 0 0 col_n[12]
port 40 s
flabel locali s -834 -457 -815 -436 5 FreeSans 40 0 0 0 col_n[13]
port 41 s
flabel locali s -798 -457 -779 -436 5 FreeSans 40 0 0 0 col_n[14]
port 42 s
flabel locali s -762 -457 -743 -436 5 FreeSans 40 0 0 0 col_n[15]
port 43 s
flabel locali s -659 -457 -625 -436 5 FreeSans 40 0 0 0 sample_n
port 44 s
flabel locali s -605 -457 -571 -436 5 FreeSans 40 0 0 0 sample
port 45 s
flabel locali s -551 -457 -483 -436 5 FreeSans 40 0 0 0 vcom
port 46 s
flabel locali s -440 -457 -294 -436 5 FreeSans 40 0 0 0 VDD
port 61 s
flabel metal4 s -2452 -436 -2245 9494 0 FreeSans 800 90 0 0 VDD
port 61 nsew
flabel metal4 s -2157 -217 -1950 9494 0 FreeSans 800 90 0 0 VSS
port 62 nsew
flabel locali s -251 -457 -105 -436 5 FreeSans 40 0 0 0 VSS
port 62 s
flabel locali s 929 -457 946 -436 5 FreeSans 80 0 0 0 row_n[0]
port 70 s
flabel locali s 1431 -457 1448 -436 5 FreeSans 80 0 0 0 row_n[1]
port 71 s
flabel locali s 1933 -457 1950 -436 5 FreeSans 80 0 0 0 row_n[2]
port 72 s
flabel locali s 2435 -457 2452 -436 5 FreeSans 80 0 0 0 row_n[3]
port 73 s
flabel locali s 2937 -457 2954 -436 5 FreeSans 80 0 0 0 row_n[4]
port 74 s
flabel locali s 3439 -457 3456 -436 5 FreeSans 80 0 0 0 row_n[5]
port 75 s
flabel locali s 3941 -457 3958 -436 5 FreeSans 80 0 0 0 row_n[6]
port 76 s
flabel locali s 4443 -457 4460 -436 5 FreeSans 80 0 0 0 row_n[7]
port 77 s
flabel locali s 4945 -457 4962 -436 5 FreeSans 80 0 0 0 row_n[8]
port 78 s
flabel locali s 5447 -457 5464 -436 5 FreeSans 80 0 0 0 row_n[9]
port 79 s
flabel locali s 5949 -457 5966 -436 5 FreeSans 80 0 0 0 row_n[10]
port 80 s
flabel locali s 6451 -457 6468 -436 5 FreeSans 80 0 0 0 row_n[11]
port 81 s
flabel locali s 6953 -457 6970 -436 5 FreeSans 80 0 0 0 row_n[12]
port 82 s
flabel locali s 7455 -457 7472 -436 5 FreeSans 80 0 0 0 row_n[13]
port 83 s
flabel locali s 7957 -457 7974 -436 5 FreeSans 80 0 0 0 row_n[14]
port 84 s
flabel locali s 8459 -457 8476 -436 5 FreeSans 80 0 0 0 row_n[15]
port 85 s
flabel locali s 8961 -457 8978 -436 5 FreeSans 80 0 0 0 row_n[16]
port 86 s
flabel locali s 9463 -457 9480 -436 5 FreeSans 80 0 0 0 row_n[17]
port 87 s
flabel locali s 9965 -457 9982 -436 5 FreeSans 80 0 0 0 row_n[18]
port 88 s
flabel locali s 10467 -457 10484 -436 5 FreeSans 80 0 0 0 row_n[19]
port 89 s
flabel locali s 10969 -457 10986 -436 5 FreeSans 80 0 0 0 row_n[20]
port 90 s
flabel locali s 11471 -457 11488 -436 5 FreeSans 80 0 0 0 row_n[21]
port 91 s
flabel locali s 11973 -457 11990 -436 5 FreeSans 80 0 0 0 row_n[22]
port 92 s
flabel locali s 12475 -457 12492 -436 5 FreeSans 80 0 0 0 row_n[23]
port 93 s
flabel locali s 12977 -457 12994 -436 5 FreeSans 80 0 0 0 row_n[24]
port 94 s
flabel locali s 4779 -457 4796 -436 5 FreeSans 80 0 0 0 en_n_bit[2]
port 102 s
flabel locali s 8795 -457 8812 -436 5 FreeSans 80 0 0 0 en_n_bit[1]
port 103 s
flabel locali s 12811 -457 12828 -436 5 FreeSans 80 0 0 0 en_n_bit[0]
port 104 s
flabel locali s 13079 -457 13096 -436 5 FreeSans 80 0 0 0 row_n[25]
port 95 s
flabel locali s 13181 -457 13198 -436 5 FreeSans 80 0 0 0 row_n[26]
port 96 s
flabel locali s 13283 -457 13300 -436 5 FreeSans 80 0 0 0 row_n[27]
port 97 s
flabel locali s 13385 -457 13402 -436 5 FreeSans 80 0 0 0 row_n[28]
port 98 s
flabel locali s 13487 -457 13504 -436 5 FreeSans 80 0 0 0 row_n[29]
port 99 s
flabel locali s 13589 -457 13606 -436 5 FreeSans 80 0 0 0 row_n[30]
port 100 s
flabel locali s 13691 -457 13708 -436 5 FreeSans 80 0 0 0 row_n[31]
port 101 s
flabel locali s 16043 -456 16060 -435 5 FreeSans 80 90 0 0 sw_n
port 110 s
flabel locali s 16104 -456 16121 -435 5 FreeSans 80 90 0 0 sw
port 111 s
flabel metal4 s 16300 -456 16330 -427 5 FreeSans 80 0 0 0 ctop
port 115 s
flabel locali s 17167 -392 17315 -370 0 FreeSans 160 0 0 0 VSS
port 62 nsew
flabel locali s 17355 -392 17503 -370 0 FreeSans 160 0 0 0 VDD
port 61 nsew
flabel metal4 s 17989 -371 18196 9495 0 FreeSans 800 90 0 0 VDD
port 117 nsew
flabel metal4 s 17694 -152 17901 9494 0 FreeSans 800 90 0 0 VSS
port 119 nsew
flabel metal1 s 18102 -453 18196 -429 0 FreeSans 80 0 0 0 analog_in
port 122 nsew
<< end >>
