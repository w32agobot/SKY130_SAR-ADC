magic
tech sky130A
timestamp 1658934595
<< metal2 >>
rect 7 530 397 540
rect 7 502 18 530
rect 46 502 358 530
rect 386 502 397 530
rect 7 411 397 502
rect 7 380 18 411
rect 46 380 358 411
rect 386 380 397 411
rect 7 289 397 380
rect 7 258 18 289
rect 46 258 358 289
rect 386 258 397 289
rect 7 168 397 258
rect 7 137 18 168
rect 46 137 397 168
rect 7 46 397 137
rect 7 18 18 46
rect 46 18 358 46
rect 386 18 397 46
rect 7 7 397 18
<< via2 >>
rect 18 502 46 530
rect 358 502 386 530
rect 18 380 46 411
rect 358 380 386 411
rect 18 258 46 289
rect 358 258 386 289
rect 18 137 46 168
rect 18 18 46 46
rect 358 18 386 46
<< metal3 >>
rect 15 530 389 533
rect 15 502 18 530
rect 46 503 358 530
rect 46 502 49 503
rect 15 499 49 502
rect 355 502 358 503
rect 386 502 389 530
rect 355 499 389 502
rect 15 415 45 499
rect 75 441 155 473
rect 187 441 217 473
rect 249 441 328 473
rect 359 415 389 499
rect 15 411 49 415
rect 355 411 389 415
rect 15 380 18 411
rect 46 381 358 411
rect 46 380 49 381
rect 15 377 49 380
rect 355 380 358 381
rect 386 380 389 411
rect 355 377 389 380
rect 15 293 45 377
rect 75 319 155 351
rect 187 319 217 351
rect 249 319 328 351
rect 359 293 389 377
rect 15 289 49 293
rect 355 289 389 293
rect 15 258 18 289
rect 46 259 358 289
rect 46 258 49 259
rect 15 255 49 258
rect 355 258 358 259
rect 386 258 389 289
rect 355 255 389 258
rect 15 171 45 255
rect 75 197 155 229
rect 187 197 217 229
rect 249 197 328 229
rect 359 171 389 255
rect 15 168 49 171
rect 15 137 18 168
rect 46 167 49 168
rect 355 167 389 171
rect 46 137 389 167
rect 15 133 49 137
rect 355 133 389 137
rect 15 49 45 133
rect 75 75 155 107
rect 187 75 217 107
rect 249 75 328 107
rect 359 49 389 133
rect 15 46 49 49
rect 15 18 18 46
rect 46 45 49 46
rect 355 46 389 49
rect 355 45 358 46
rect 46 18 358 45
rect 386 18 389 46
rect 15 15 389 18
<< via3 >>
rect 155 441 187 473
rect 217 441 249 473
rect 155 319 187 351
rect 217 319 249 351
rect 155 197 187 229
rect 217 197 249 229
rect 155 75 187 107
rect 217 75 249 107
<< metal4 >>
rect 7 543 397 573
rect 187 474 217 543
rect 154 473 250 474
rect 154 441 155 473
rect 187 441 217 473
rect 249 441 250 473
rect 154 440 250 441
rect 187 352 217 440
rect 154 351 250 352
rect 154 319 155 351
rect 187 319 217 351
rect 249 319 250 351
rect 154 318 250 319
rect 187 230 217 318
rect 154 229 250 230
rect 154 197 155 229
rect 187 197 217 229
rect 249 197 250 229
rect 154 196 250 197
rect 187 108 217 196
rect 154 107 250 108
rect 154 75 155 107
rect 187 75 217 107
rect 249 75 250 107
rect 154 74 250 75
rect 187 4 217 74
rect 7 -26 397 4
<< comment >>
rect 0 364 15 379
rect 389 364 404 379
rect 0 0 15 15
rect 389 0 404 15
<< labels >>
rlabel metal4 7 -26 7 -26 1 ctop
rlabel metal2 7 33 7 33 1 cbot
<< end >>
