magic
tech sky130A
magscale 1 2
timestamp 1663935139
<< nwell >>
rect 3676 3604 5258 3608
rect 1318 3200 5258 3604
rect 1318 3182 3610 3200
rect 1844 3180 2086 3182
rect 2452 2832 3610 3182
rect 4248 3152 5258 3200
rect 846 2414 1288 2812
rect 4408 2460 4922 2512
rect 3712 2056 4922 2460
<< pwell >>
rect 1464 5198 1944 5378
rect 4044 5198 4524 5378
rect 1004 5118 2254 5198
rect 2904 5118 3084 5198
rect 3734 5118 4984 5198
rect 1004 4058 4984 5118
rect 1004 3978 2254 4058
rect 2904 3978 3084 4058
rect 3734 3978 4984 4058
rect 1464 3798 1944 3978
rect 4044 3798 4524 3978
rect 1464 1608 1944 1788
rect 4044 1608 4524 1788
rect 1004 1528 2254 1608
rect 2904 1528 3084 1608
rect 3734 1528 4984 1608
rect 1004 468 4984 1528
rect 1004 388 2254 468
rect 2904 388 3084 468
rect 3734 388 4984 468
rect 1464 208 1944 388
rect 4044 208 4524 388
<< nmos >>
rect 1154 4198 4834 4978
rect 3810 2936 3840 3036
rect 3906 2936 3936 3036
rect 4002 2936 4032 3036
rect 4346 3000 4376 3084
rect 4442 3000 4472 3084
rect 4842 3000 4872 3084
rect 4938 3000 4968 3084
rect 1418 2468 1448 2868
rect 1514 2468 1544 2868
rect 1610 2468 1640 2868
rect 1706 2468 1736 2868
rect 1802 2468 1832 2868
rect 1898 2468 1928 2868
rect 1994 2468 2024 2868
rect 2090 2468 2120 2868
rect 908 2258 992 2288
rect 1142 2258 1226 2288
rect 1418 2208 1448 2308
rect 1514 2208 1544 2308
rect 1610 2208 1640 2308
rect 1706 2208 1736 2308
rect 1802 2208 1832 2308
rect 1898 2208 1928 2308
rect 1994 2208 2024 2308
rect 2090 2208 2120 2308
rect 2872 2202 2902 2602
rect 2968 2202 2998 2602
rect 3064 2202 3094 2602
rect 3160 2202 3190 2602
rect 3810 2624 3840 2724
rect 3906 2624 3936 2724
rect 4002 2624 4032 2724
rect 4506 2580 4536 2664
rect 4602 2580 4632 2664
rect 1154 608 4834 1388
<< pmos >>
rect 1418 3282 1448 3382
rect 1514 3282 1544 3382
rect 1610 3282 1640 3382
rect 1706 3282 1736 3382
rect 1802 3282 1832 3382
rect 1898 3282 1928 3382
rect 1994 3282 2024 3382
rect 2090 3282 2120 3382
rect 2550 2932 2580 3332
rect 2646 2932 2676 3332
rect 2872 2932 2902 3332
rect 2968 2932 2998 3332
rect 3064 2932 3094 3332
rect 3160 2932 3190 3332
rect 3386 2932 3416 3332
rect 3482 2932 3512 3332
rect 3810 3262 3840 3462
rect 3906 3262 3936 3462
rect 4002 3262 4032 3462
rect 4346 3254 4376 3414
rect 4442 3254 4472 3414
rect 4538 3254 4568 3414
rect 4634 3254 4664 3414
rect 4842 3254 4872 3414
rect 4938 3254 4968 3414
rect 5034 3254 5064 3414
rect 5130 3254 5160 3414
rect 908 2600 996 2630
rect 1142 2600 1230 2630
rect 908 2508 996 2538
rect 1142 2508 1230 2538
rect 3810 2198 3840 2398
rect 3906 2198 3936 2398
rect 4002 2198 4032 2398
rect 4506 2250 4536 2410
rect 4602 2250 4632 2410
rect 4698 2250 4728 2410
rect 4794 2250 4824 2410
<< ndiff >>
rect 1154 5098 4834 5118
rect 1154 4998 1164 5098
rect 1284 4998 1324 5098
rect 1444 4998 1484 5098
rect 1604 4998 1644 5098
rect 1764 4998 1804 5098
rect 1924 4998 1964 5098
rect 2084 4998 2124 5098
rect 2244 4998 3744 5098
rect 3864 4998 3904 5098
rect 4024 4998 4064 5098
rect 4184 4998 4224 5098
rect 4344 4998 4384 5098
rect 4504 4998 4544 5098
rect 4664 4998 4704 5098
rect 4824 4998 4834 5098
rect 1154 4978 4834 4998
rect 1154 4178 4834 4198
rect 1154 4078 1164 4178
rect 1284 4078 1324 4178
rect 1444 4078 1484 4178
rect 1604 4078 1644 4178
rect 1764 4078 1804 4178
rect 1924 4078 1964 4178
rect 2084 4078 2124 4178
rect 2244 4078 3744 4178
rect 3864 4078 3904 4178
rect 4024 4078 4064 4178
rect 4184 4078 4224 4178
rect 4344 4078 4384 4178
rect 4504 4078 4544 4178
rect 4664 4078 4704 4178
rect 4824 4078 4834 4178
rect 1154 4058 4834 4078
rect 3748 3024 3810 3036
rect 3748 2948 3760 3024
rect 3794 2948 3810 3024
rect 3748 2936 3810 2948
rect 3840 3024 3906 3036
rect 3840 2948 3856 3024
rect 3890 2948 3906 3024
rect 3840 2936 3906 2948
rect 3936 3024 4002 3036
rect 3936 2948 3952 3024
rect 3986 2948 4002 3024
rect 3936 2936 4002 2948
rect 4032 3024 4094 3036
rect 4032 2948 4048 3024
rect 4082 2948 4094 3024
rect 4032 2936 4094 2948
rect 4284 3072 4346 3084
rect 4284 3012 4296 3072
rect 4330 3012 4346 3072
rect 4284 3000 4346 3012
rect 4376 3072 4442 3084
rect 4376 3012 4392 3072
rect 4426 3012 4442 3072
rect 4376 3000 4442 3012
rect 4472 3072 4534 3084
rect 4472 3012 4488 3072
rect 4522 3012 4534 3072
rect 4472 3000 4534 3012
rect 4780 3072 4842 3084
rect 4780 3012 4792 3072
rect 4826 3012 4842 3072
rect 4780 3000 4842 3012
rect 4872 3072 4938 3084
rect 4872 3012 4888 3072
rect 4922 3012 4938 3072
rect 4872 3000 4938 3012
rect 4968 3072 5030 3084
rect 4968 3012 4984 3072
rect 5018 3012 5030 3072
rect 4968 3000 5030 3012
rect 1356 2856 1418 2868
rect 1356 2480 1368 2856
rect 1402 2480 1418 2856
rect 1356 2468 1418 2480
rect 1448 2856 1514 2868
rect 1448 2480 1464 2856
rect 1498 2480 1514 2856
rect 1448 2468 1514 2480
rect 1544 2856 1610 2868
rect 1544 2480 1560 2856
rect 1594 2480 1610 2856
rect 1544 2468 1610 2480
rect 1640 2856 1706 2868
rect 1640 2480 1656 2856
rect 1690 2480 1706 2856
rect 1640 2468 1706 2480
rect 1736 2856 1802 2868
rect 1736 2480 1752 2856
rect 1786 2480 1802 2856
rect 1736 2468 1802 2480
rect 1832 2856 1898 2868
rect 1832 2480 1848 2856
rect 1882 2480 1898 2856
rect 1832 2468 1898 2480
rect 1928 2856 1994 2868
rect 1928 2480 1944 2856
rect 1978 2480 1994 2856
rect 1928 2468 1994 2480
rect 2024 2856 2090 2868
rect 2024 2480 2040 2856
rect 2074 2480 2090 2856
rect 2024 2468 2090 2480
rect 2120 2856 2182 2868
rect 2120 2480 2136 2856
rect 2170 2480 2182 2856
rect 2120 2468 2182 2480
rect 2810 2590 2872 2602
rect 908 2334 992 2346
rect 908 2300 920 2334
rect 980 2300 992 2334
rect 908 2288 992 2300
rect 1142 2334 1226 2346
rect 1142 2300 1154 2334
rect 1214 2300 1226 2334
rect 1142 2288 1226 2300
rect 1356 2296 1418 2308
rect 908 2246 992 2258
rect 908 2212 920 2246
rect 980 2212 992 2246
rect 908 2200 992 2212
rect 1142 2246 1226 2258
rect 1142 2212 1154 2246
rect 1214 2212 1226 2246
rect 1142 2200 1226 2212
rect 1356 2220 1368 2296
rect 1402 2220 1418 2296
rect 1356 2208 1418 2220
rect 1448 2296 1514 2308
rect 1448 2220 1464 2296
rect 1498 2220 1514 2296
rect 1448 2208 1514 2220
rect 1544 2296 1610 2308
rect 1544 2220 1560 2296
rect 1594 2220 1610 2296
rect 1544 2208 1610 2220
rect 1640 2296 1706 2308
rect 1640 2220 1656 2296
rect 1690 2220 1706 2296
rect 1640 2208 1706 2220
rect 1736 2296 1802 2308
rect 1736 2220 1752 2296
rect 1786 2220 1802 2296
rect 1736 2208 1802 2220
rect 1832 2296 1898 2308
rect 1832 2220 1848 2296
rect 1882 2220 1898 2296
rect 1832 2208 1898 2220
rect 1928 2296 1994 2308
rect 1928 2220 1944 2296
rect 1978 2220 1994 2296
rect 1928 2208 1994 2220
rect 2024 2296 2090 2308
rect 2024 2220 2040 2296
rect 2074 2220 2090 2296
rect 2024 2208 2090 2220
rect 2120 2296 2182 2308
rect 2120 2220 2136 2296
rect 2170 2220 2182 2296
rect 2120 2208 2182 2220
rect 2810 2214 2822 2590
rect 2856 2214 2872 2590
rect 2810 2202 2872 2214
rect 2902 2590 2968 2602
rect 2902 2214 2918 2590
rect 2952 2214 2968 2590
rect 2902 2202 2968 2214
rect 2998 2590 3064 2602
rect 2998 2214 3014 2590
rect 3048 2214 3064 2590
rect 2998 2202 3064 2214
rect 3094 2590 3160 2602
rect 3094 2214 3110 2590
rect 3144 2214 3160 2590
rect 3094 2202 3160 2214
rect 3190 2590 3252 2602
rect 3190 2214 3206 2590
rect 3240 2214 3252 2590
rect 3748 2712 3810 2724
rect 3748 2636 3760 2712
rect 3794 2636 3810 2712
rect 3748 2624 3810 2636
rect 3840 2712 3906 2724
rect 3840 2636 3856 2712
rect 3890 2636 3906 2712
rect 3840 2624 3906 2636
rect 3936 2712 4002 2724
rect 3936 2636 3952 2712
rect 3986 2636 4002 2712
rect 3936 2624 4002 2636
rect 4032 2712 4094 2724
rect 4032 2636 4048 2712
rect 4082 2636 4094 2712
rect 4032 2624 4094 2636
rect 4444 2652 4506 2664
rect 4444 2592 4456 2652
rect 4490 2592 4506 2652
rect 4444 2580 4506 2592
rect 4536 2652 4602 2664
rect 4536 2592 4552 2652
rect 4586 2592 4602 2652
rect 4536 2580 4602 2592
rect 4632 2652 4694 2664
rect 4632 2592 4648 2652
rect 4682 2592 4694 2652
rect 4632 2580 4694 2592
rect 3190 2202 3252 2214
rect 1154 1508 4834 1528
rect 1154 1408 1164 1508
rect 1284 1408 1324 1508
rect 1444 1408 1484 1508
rect 1604 1408 1644 1508
rect 1764 1408 1804 1508
rect 1924 1408 1964 1508
rect 2084 1408 2124 1508
rect 2244 1408 3744 1508
rect 3864 1408 3904 1508
rect 4024 1408 4064 1508
rect 4184 1408 4224 1508
rect 4344 1408 4384 1508
rect 4504 1408 4544 1508
rect 4664 1408 4704 1508
rect 4824 1408 4834 1508
rect 1154 1388 4834 1408
rect 1154 588 4834 608
rect 1154 488 1164 588
rect 1284 488 1324 588
rect 1444 488 1484 588
rect 1604 488 1644 588
rect 1764 488 1804 588
rect 1924 488 1964 588
rect 2084 488 2124 588
rect 2244 488 3744 588
rect 3864 488 3904 588
rect 4024 488 4064 588
rect 4184 488 4224 588
rect 4344 488 4384 588
rect 4504 488 4544 588
rect 4664 488 4704 588
rect 4824 488 4834 588
rect 1154 468 4834 488
<< pdiff >>
rect 3748 3450 3810 3462
rect 1356 3370 1418 3382
rect 1356 3294 1368 3370
rect 1402 3294 1418 3370
rect 1356 3282 1418 3294
rect 1448 3370 1514 3382
rect 1448 3294 1464 3370
rect 1498 3294 1514 3370
rect 1448 3282 1514 3294
rect 1544 3370 1610 3382
rect 1544 3294 1560 3370
rect 1594 3294 1610 3370
rect 1544 3282 1610 3294
rect 1640 3370 1706 3382
rect 1640 3294 1656 3370
rect 1690 3294 1706 3370
rect 1640 3282 1706 3294
rect 1736 3370 1802 3382
rect 1736 3294 1752 3370
rect 1786 3294 1802 3370
rect 1736 3282 1802 3294
rect 1832 3370 1898 3382
rect 1832 3294 1848 3370
rect 1882 3294 1898 3370
rect 1832 3282 1898 3294
rect 1928 3370 1994 3382
rect 1928 3294 1944 3370
rect 1978 3294 1994 3370
rect 1928 3282 1994 3294
rect 2024 3370 2090 3382
rect 2024 3294 2040 3370
rect 2074 3294 2090 3370
rect 2024 3282 2090 3294
rect 2120 3370 2182 3382
rect 2120 3294 2136 3370
rect 2170 3294 2182 3370
rect 2120 3282 2182 3294
rect 2488 3320 2550 3332
rect 2488 2944 2500 3320
rect 2534 2944 2550 3320
rect 2488 2932 2550 2944
rect 2580 3320 2646 3332
rect 2580 2944 2596 3320
rect 2630 2944 2646 3320
rect 2580 2932 2646 2944
rect 2676 3320 2738 3332
rect 2676 2944 2692 3320
rect 2726 2944 2738 3320
rect 2676 2932 2738 2944
rect 2810 3320 2872 3332
rect 2810 2944 2822 3320
rect 2856 2944 2872 3320
rect 2810 2932 2872 2944
rect 2902 3320 2968 3332
rect 2902 2944 2918 3320
rect 2952 2944 2968 3320
rect 2902 2932 2968 2944
rect 2998 3320 3064 3332
rect 2998 2944 3014 3320
rect 3048 2944 3064 3320
rect 2998 2932 3064 2944
rect 3094 3320 3160 3332
rect 3094 2944 3110 3320
rect 3144 2944 3160 3320
rect 3094 2932 3160 2944
rect 3190 3320 3252 3332
rect 3190 2944 3206 3320
rect 3240 2944 3252 3320
rect 3190 2932 3252 2944
rect 3324 3320 3386 3332
rect 3324 2944 3336 3320
rect 3370 2944 3386 3320
rect 3324 2932 3386 2944
rect 3416 3320 3482 3332
rect 3416 2944 3432 3320
rect 3466 2944 3482 3320
rect 3416 2932 3482 2944
rect 3512 3320 3574 3332
rect 3512 2944 3528 3320
rect 3562 2944 3574 3320
rect 3748 3274 3760 3450
rect 3794 3274 3810 3450
rect 3748 3262 3810 3274
rect 3840 3450 3906 3462
rect 3840 3274 3856 3450
rect 3890 3274 3906 3450
rect 3840 3262 3906 3274
rect 3936 3450 4002 3462
rect 3936 3274 3952 3450
rect 3986 3274 4002 3450
rect 3936 3262 4002 3274
rect 4032 3450 4094 3462
rect 4032 3274 4048 3450
rect 4082 3274 4094 3450
rect 4032 3262 4094 3274
rect 4284 3402 4346 3414
rect 4284 3266 4296 3402
rect 4330 3266 4346 3402
rect 4284 3254 4346 3266
rect 4376 3402 4442 3414
rect 4376 3266 4392 3402
rect 4426 3266 4442 3402
rect 4376 3254 4442 3266
rect 4472 3402 4538 3414
rect 4472 3266 4488 3402
rect 4522 3266 4538 3402
rect 4472 3254 4538 3266
rect 4568 3402 4634 3414
rect 4568 3266 4584 3402
rect 4618 3266 4634 3402
rect 4568 3254 4634 3266
rect 4664 3402 4726 3414
rect 4664 3266 4680 3402
rect 4714 3266 4726 3402
rect 4664 3254 4726 3266
rect 4780 3402 4842 3414
rect 4780 3266 4792 3402
rect 4826 3266 4842 3402
rect 4780 3254 4842 3266
rect 4872 3402 4938 3414
rect 4872 3266 4888 3402
rect 4922 3266 4938 3402
rect 4872 3254 4938 3266
rect 4968 3402 5034 3414
rect 4968 3266 4984 3402
rect 5018 3266 5034 3402
rect 4968 3254 5034 3266
rect 5064 3402 5130 3414
rect 5064 3266 5080 3402
rect 5114 3266 5130 3402
rect 5064 3254 5130 3266
rect 5160 3402 5222 3414
rect 5160 3266 5176 3402
rect 5210 3266 5222 3402
rect 5160 3254 5222 3266
rect 3512 2932 3574 2944
rect 908 2678 996 2686
rect 908 2644 920 2678
rect 980 2644 996 2678
rect 908 2630 996 2644
rect 1142 2678 1230 2686
rect 1142 2644 1154 2678
rect 1214 2644 1230 2678
rect 1142 2630 1230 2644
rect 908 2586 996 2600
rect 908 2552 920 2586
rect 980 2552 996 2586
rect 908 2538 996 2552
rect 1142 2586 1230 2600
rect 1142 2552 1154 2586
rect 1214 2552 1230 2586
rect 1142 2538 1230 2552
rect 908 2496 996 2508
rect 908 2462 920 2496
rect 980 2462 996 2496
rect 908 2450 996 2462
rect 1142 2496 1230 2508
rect 1142 2462 1154 2496
rect 1214 2462 1230 2496
rect 1142 2450 1230 2462
rect 4444 2398 4506 2410
rect 3748 2386 3810 2398
rect 3748 2210 3760 2386
rect 3794 2210 3810 2386
rect 3748 2198 3810 2210
rect 3840 2386 3906 2398
rect 3840 2210 3856 2386
rect 3890 2210 3906 2386
rect 3840 2198 3906 2210
rect 3936 2386 4002 2398
rect 3936 2210 3952 2386
rect 3986 2210 4002 2386
rect 3936 2198 4002 2210
rect 4032 2386 4094 2398
rect 4032 2210 4048 2386
rect 4082 2210 4094 2386
rect 4444 2262 4456 2398
rect 4490 2262 4506 2398
rect 4444 2250 4506 2262
rect 4536 2398 4602 2410
rect 4536 2262 4552 2398
rect 4586 2262 4602 2398
rect 4536 2250 4602 2262
rect 4632 2398 4698 2410
rect 4632 2262 4648 2398
rect 4682 2262 4698 2398
rect 4632 2250 4698 2262
rect 4728 2398 4794 2410
rect 4728 2262 4744 2398
rect 4778 2262 4794 2398
rect 4728 2250 4794 2262
rect 4824 2398 4886 2410
rect 4824 2262 4840 2398
rect 4874 2262 4886 2398
rect 4824 2250 4886 2262
rect 4032 2198 4094 2210
<< ndiffc >>
rect 1164 4998 1284 5098
rect 1324 4998 1444 5098
rect 1484 4998 1604 5098
rect 1644 4998 1764 5098
rect 1804 4998 1924 5098
rect 1964 4998 2084 5098
rect 2124 4998 2244 5098
rect 3744 4998 3864 5098
rect 3904 4998 4024 5098
rect 4064 4998 4184 5098
rect 4224 4998 4344 5098
rect 4384 4998 4504 5098
rect 4544 4998 4664 5098
rect 4704 4998 4824 5098
rect 1164 4078 1284 4178
rect 1324 4078 1444 4178
rect 1484 4078 1604 4178
rect 1644 4078 1764 4178
rect 1804 4078 1924 4178
rect 1964 4078 2084 4178
rect 2124 4078 2244 4178
rect 3744 4078 3864 4178
rect 3904 4078 4024 4178
rect 4064 4078 4184 4178
rect 4224 4078 4344 4178
rect 4384 4078 4504 4178
rect 4544 4078 4664 4178
rect 4704 4078 4824 4178
rect 3760 2948 3794 3024
rect 3856 2948 3890 3024
rect 3952 2948 3986 3024
rect 4048 2948 4082 3024
rect 4296 3012 4330 3072
rect 4392 3012 4426 3072
rect 4488 3012 4522 3072
rect 4792 3012 4826 3072
rect 4888 3012 4922 3072
rect 4984 3012 5018 3072
rect 1368 2480 1402 2856
rect 1464 2480 1498 2856
rect 1560 2480 1594 2856
rect 1656 2480 1690 2856
rect 1752 2480 1786 2856
rect 1848 2480 1882 2856
rect 1944 2480 1978 2856
rect 2040 2480 2074 2856
rect 2136 2480 2170 2856
rect 920 2300 980 2334
rect 1154 2300 1214 2334
rect 920 2212 980 2246
rect 1154 2212 1214 2246
rect 1368 2220 1402 2296
rect 1464 2220 1498 2296
rect 1560 2220 1594 2296
rect 1656 2220 1690 2296
rect 1752 2220 1786 2296
rect 1848 2220 1882 2296
rect 1944 2220 1978 2296
rect 2040 2220 2074 2296
rect 2136 2220 2170 2296
rect 2822 2214 2856 2590
rect 2918 2214 2952 2590
rect 3014 2214 3048 2590
rect 3110 2214 3144 2590
rect 3206 2214 3240 2590
rect 3760 2636 3794 2712
rect 3856 2636 3890 2712
rect 3952 2636 3986 2712
rect 4048 2636 4082 2712
rect 4456 2592 4490 2652
rect 4552 2592 4586 2652
rect 4648 2592 4682 2652
rect 1164 1408 1284 1508
rect 1324 1408 1444 1508
rect 1484 1408 1604 1508
rect 1644 1408 1764 1508
rect 1804 1408 1924 1508
rect 1964 1408 2084 1508
rect 2124 1408 2244 1508
rect 3744 1408 3864 1508
rect 3904 1408 4024 1508
rect 4064 1408 4184 1508
rect 4224 1408 4344 1508
rect 4384 1408 4504 1508
rect 4544 1408 4664 1508
rect 4704 1408 4824 1508
rect 1164 488 1284 588
rect 1324 488 1444 588
rect 1484 488 1604 588
rect 1644 488 1764 588
rect 1804 488 1924 588
rect 1964 488 2084 588
rect 2124 488 2244 588
rect 3744 488 3864 588
rect 3904 488 4024 588
rect 4064 488 4184 588
rect 4224 488 4344 588
rect 4384 488 4504 588
rect 4544 488 4664 588
rect 4704 488 4824 588
<< pdiffc >>
rect 1368 3294 1402 3370
rect 1464 3294 1498 3370
rect 1560 3294 1594 3370
rect 1656 3294 1690 3370
rect 1752 3294 1786 3370
rect 1848 3294 1882 3370
rect 1944 3294 1978 3370
rect 2040 3294 2074 3370
rect 2136 3294 2170 3370
rect 2500 2944 2534 3320
rect 2596 2944 2630 3320
rect 2692 2944 2726 3320
rect 2822 2944 2856 3320
rect 2918 2944 2952 3320
rect 3014 2944 3048 3320
rect 3110 2944 3144 3320
rect 3206 2944 3240 3320
rect 3336 2944 3370 3320
rect 3432 2944 3466 3320
rect 3528 2944 3562 3320
rect 3760 3274 3794 3450
rect 3856 3274 3890 3450
rect 3952 3274 3986 3450
rect 4048 3274 4082 3450
rect 4296 3266 4330 3402
rect 4392 3266 4426 3402
rect 4488 3266 4522 3402
rect 4584 3266 4618 3402
rect 4680 3266 4714 3402
rect 4792 3266 4826 3402
rect 4888 3266 4922 3402
rect 4984 3266 5018 3402
rect 5080 3266 5114 3402
rect 5176 3266 5210 3402
rect 920 2644 980 2678
rect 1154 2644 1214 2678
rect 920 2552 980 2586
rect 1154 2552 1214 2586
rect 920 2462 980 2496
rect 1154 2462 1214 2496
rect 3760 2210 3794 2386
rect 3856 2210 3890 2386
rect 3952 2210 3986 2386
rect 4048 2210 4082 2386
rect 4456 2262 4490 2398
rect 4552 2262 4586 2398
rect 4648 2262 4682 2398
rect 4744 2262 4778 2398
rect 4840 2262 4874 2398
<< psubdiff >>
rect 988 5540 1110 5566
rect 988 5466 1012 5540
rect 1086 5466 1110 5540
rect 988 5442 1110 5466
rect 1536 5540 1658 5566
rect 1536 5466 1560 5540
rect 1634 5466 1658 5540
rect 1536 5442 1658 5466
rect 2084 5540 2206 5566
rect 2084 5466 2108 5540
rect 2182 5466 2206 5540
rect 2084 5442 2206 5466
rect 2632 5540 2754 5566
rect 2632 5466 2656 5540
rect 2730 5466 2754 5540
rect 2632 5442 2754 5466
rect 3180 5540 3302 5566
rect 3180 5466 3204 5540
rect 3278 5466 3302 5540
rect 3180 5442 3302 5466
rect 3710 5540 3832 5566
rect 3710 5466 3734 5540
rect 3808 5466 3832 5540
rect 3710 5442 3832 5466
rect 4258 5540 4380 5566
rect 4258 5466 4282 5540
rect 4356 5466 4380 5540
rect 4258 5442 4380 5466
rect 4808 5540 4930 5566
rect 4808 5466 4832 5540
rect 4906 5466 4930 5540
rect 4808 5442 4930 5466
rect 622 5398 744 5424
rect 622 5324 646 5398
rect 720 5324 744 5398
rect 622 5300 744 5324
rect 5304 5328 5426 5354
rect 1474 5278 1934 5298
rect 1474 5228 1504 5278
rect 1904 5228 1934 5278
rect 1474 5208 1934 5228
rect 4054 5278 4514 5298
rect 4054 5228 4084 5278
rect 4484 5228 4514 5278
rect 5304 5254 5328 5328
rect 5402 5254 5426 5328
rect 5304 5230 5426 5254
rect 4054 5208 4514 5228
rect 622 4924 744 4950
rect 622 4850 646 4924
rect 720 4850 744 4924
rect 622 4826 744 4850
rect 622 4450 744 4476
rect 622 4376 646 4450
rect 720 4376 744 4450
rect 622 4352 744 4376
rect 5304 4852 5426 4878
rect 5304 4778 5328 4852
rect 5402 4778 5426 4852
rect 5304 4754 5426 4778
rect 5304 4378 5426 4404
rect 5304 4304 5328 4378
rect 5402 4304 5426 4378
rect 5304 4280 5426 4304
rect 622 3976 744 4002
rect 622 3902 646 3976
rect 720 3902 744 3976
rect 622 3878 744 3902
rect 1474 3948 1934 3968
rect 1474 3898 1504 3948
rect 1904 3898 1934 3948
rect 1474 3878 1934 3898
rect 4054 3948 4514 3968
rect 4054 3898 4084 3948
rect 4484 3898 4514 3948
rect 4054 3878 4514 3898
rect 5302 3904 5424 3930
rect 5302 3830 5326 3904
rect 5400 3830 5424 3904
rect 5302 3812 5424 3830
rect 622 3290 744 3316
rect 622 3216 646 3290
rect 720 3216 744 3290
rect 622 3192 744 3216
rect 5302 3292 5424 3318
rect 5302 3218 5326 3292
rect 5400 3218 5424 3292
rect 5302 3194 5424 3218
rect 614 2764 736 2790
rect 614 2690 638 2764
rect 712 2690 736 2764
rect 614 2666 736 2690
rect 4368 2912 4392 2946
rect 4426 2912 4454 2946
rect 4864 2912 4888 2946
rect 4922 2912 4950 2946
rect 3748 2848 3774 2882
rect 3808 2848 3842 2882
rect 3876 2848 3910 2882
rect 3944 2848 3978 2882
rect 4012 2848 4046 2882
rect 4080 2848 4104 2882
rect 3748 2812 4104 2848
rect 3748 2778 3774 2812
rect 3808 2778 3842 2812
rect 3876 2778 3910 2812
rect 3944 2778 3978 2812
rect 4012 2778 4046 2812
rect 4080 2778 4104 2812
rect 5302 2818 5424 2844
rect 614 2290 736 2316
rect 614 2216 638 2290
rect 712 2216 736 2290
rect 614 2192 736 2216
rect 4528 2718 4552 2752
rect 4586 2718 4614 2752
rect 5302 2744 5326 2818
rect 5400 2744 5424 2818
rect 5302 2720 5424 2744
rect 908 2112 932 2146
rect 968 2112 992 2146
rect 908 2106 992 2112
rect 1142 2112 1166 2146
rect 1202 2112 1226 2146
rect 5302 2344 5424 2370
rect 5302 2270 5326 2344
rect 5400 2270 5424 2344
rect 5302 2246 5424 2270
rect 1142 2106 1226 2112
rect 2816 2054 2840 2090
rect 2876 2054 2932 2090
rect 2968 2054 3024 2090
rect 3060 2054 3116 2090
rect 3152 2054 3208 2090
rect 3244 2054 3268 2090
rect 2816 2052 3268 2054
rect 1350 2046 2168 2048
rect 1350 2010 1374 2046
rect 1410 2010 1492 2046
rect 1528 2010 1610 2046
rect 1646 2010 1728 2046
rect 1764 2010 1846 2046
rect 1882 2010 1964 2046
rect 2000 2010 2082 2046
rect 2118 2010 2168 2046
rect 1350 2006 2168 2010
rect 1474 1688 1934 1708
rect 628 1638 750 1664
rect 628 1564 652 1638
rect 726 1564 750 1638
rect 1474 1638 1504 1688
rect 1904 1638 1934 1688
rect 1474 1618 1934 1638
rect 4054 1688 4514 1708
rect 4054 1638 4084 1688
rect 4484 1638 4514 1688
rect 4054 1618 4514 1638
rect 628 1540 750 1564
rect 5302 1608 5424 1634
rect 5302 1534 5326 1608
rect 5400 1534 5424 1608
rect 5302 1510 5424 1534
rect 628 1164 750 1190
rect 628 1090 652 1164
rect 726 1090 750 1164
rect 628 1066 750 1090
rect 628 690 750 716
rect 628 616 652 690
rect 726 616 750 690
rect 628 592 750 616
rect 5302 1134 5424 1160
rect 5302 1060 5326 1134
rect 5400 1060 5424 1134
rect 5302 1036 5424 1060
rect 5302 660 5424 686
rect 5302 586 5326 660
rect 5400 586 5424 660
rect 5302 562 5424 586
rect 1474 358 1934 378
rect 1474 308 1504 358
rect 1904 308 1934 358
rect 1474 288 1934 308
rect 4054 358 4514 378
rect 4054 308 4084 358
rect 4484 308 4514 358
rect 4054 288 4514 308
rect 1158 130 1280 156
rect 1158 56 1182 130
rect 1256 56 1280 130
rect 1158 32 1280 56
rect 1706 130 1828 156
rect 1706 56 1730 130
rect 1804 56 1828 130
rect 1706 32 1828 56
rect 2254 130 2376 156
rect 2254 56 2278 130
rect 2352 56 2376 130
rect 2254 32 2376 56
rect 2802 130 2924 156
rect 2802 56 2826 130
rect 2900 56 2924 130
rect 2802 32 2924 56
rect 3350 130 3472 156
rect 3350 56 3374 130
rect 3448 56 3472 130
rect 3350 32 3472 56
rect 3898 130 4020 156
rect 3898 56 3922 130
rect 3996 56 4020 130
rect 3898 32 4020 56
rect 4448 130 4570 156
rect 4448 56 4472 130
rect 4546 56 4570 130
rect 4448 32 4570 56
<< nsubdiff >>
rect 3748 3530 3772 3568
rect 3810 3530 3848 3568
rect 3886 3530 3924 3568
rect 3962 3530 4000 3568
rect 4038 3530 4094 3568
rect 4322 3538 4352 3572
rect 4386 3538 4420 3572
rect 4454 3538 4488 3572
rect 4522 3538 4556 3572
rect 4590 3538 4624 3572
rect 4658 3538 4700 3572
rect 4818 3538 4848 3572
rect 4882 3538 4916 3572
rect 4950 3538 4984 3572
rect 5018 3538 5052 3572
rect 5086 3538 5120 3572
rect 5154 3538 5196 3572
rect 2656 3488 3380 3496
rect 1356 3478 2212 3486
rect 1356 3444 1386 3478
rect 1420 3444 1470 3478
rect 1504 3444 1554 3478
rect 1588 3444 1638 3478
rect 1672 3444 1722 3478
rect 1756 3444 1806 3478
rect 1840 3444 1890 3478
rect 1924 3444 1974 3478
rect 2008 3444 2058 3478
rect 2092 3444 2148 3478
rect 2182 3444 2212 3478
rect 2656 3454 2694 3488
rect 2728 3454 2778 3488
rect 2812 3454 2862 3488
rect 2896 3454 2946 3488
rect 2980 3454 3030 3488
rect 3064 3454 3114 3488
rect 3148 3454 3198 3488
rect 3232 3454 3282 3488
rect 3316 3454 3380 3488
rect 2656 3448 3380 3454
rect 1356 3438 2212 3444
rect 908 2740 932 2776
rect 968 2740 992 2776
rect 1142 2740 1166 2776
rect 1202 2740 1226 2776
rect 3748 2092 3772 2130
rect 3810 2092 3848 2130
rect 3886 2092 3924 2130
rect 3962 2092 4000 2130
rect 4038 2092 4094 2130
rect 4482 2092 4512 2126
rect 4546 2092 4580 2126
rect 4614 2092 4648 2126
rect 4682 2092 4716 2126
rect 4750 2092 4784 2126
rect 4818 2092 4860 2126
<< psubdiffcont >>
rect 1012 5466 1086 5540
rect 1560 5466 1634 5540
rect 2108 5466 2182 5540
rect 2656 5466 2730 5540
rect 3204 5466 3278 5540
rect 3734 5466 3808 5540
rect 4282 5466 4356 5540
rect 4832 5466 4906 5540
rect 646 5324 720 5398
rect 1504 5228 1904 5278
rect 4084 5228 4484 5278
rect 5328 5254 5402 5328
rect 646 4850 720 4924
rect 646 4376 720 4450
rect 5328 4778 5402 4852
rect 5328 4304 5402 4378
rect 646 3902 720 3976
rect 1504 3898 1904 3948
rect 4084 3898 4484 3948
rect 5326 3830 5400 3904
rect 646 3216 720 3290
rect 5326 3218 5400 3292
rect 638 2690 712 2764
rect 4392 2912 4426 2946
rect 4888 2912 4922 2946
rect 3774 2848 3808 2882
rect 3842 2848 3876 2882
rect 3910 2848 3944 2882
rect 3978 2848 4012 2882
rect 4046 2848 4080 2882
rect 3774 2778 3808 2812
rect 3842 2778 3876 2812
rect 3910 2778 3944 2812
rect 3978 2778 4012 2812
rect 4046 2778 4080 2812
rect 638 2216 712 2290
rect 4552 2718 4586 2752
rect 5326 2744 5400 2818
rect 932 2112 968 2146
rect 1166 2112 1202 2146
rect 5326 2270 5400 2344
rect 2840 2054 2876 2090
rect 2932 2054 2968 2090
rect 3024 2054 3060 2090
rect 3116 2054 3152 2090
rect 3208 2054 3244 2090
rect 1374 2010 1410 2046
rect 1492 2010 1528 2046
rect 1610 2010 1646 2046
rect 1728 2010 1764 2046
rect 1846 2010 1882 2046
rect 1964 2010 2000 2046
rect 2082 2010 2118 2046
rect 652 1564 726 1638
rect 1504 1638 1904 1688
rect 4084 1638 4484 1688
rect 5326 1534 5400 1608
rect 652 1090 726 1164
rect 652 616 726 690
rect 5326 1060 5400 1134
rect 5326 586 5400 660
rect 1504 308 1904 358
rect 4084 308 4484 358
rect 1182 56 1256 130
rect 1730 56 1804 130
rect 2278 56 2352 130
rect 2826 56 2900 130
rect 3374 56 3448 130
rect 3922 56 3996 130
rect 4472 56 4546 130
<< nsubdiffcont >>
rect 3772 3530 3810 3568
rect 3848 3530 3886 3568
rect 3924 3530 3962 3568
rect 4000 3530 4038 3568
rect 4352 3538 4386 3572
rect 4420 3538 4454 3572
rect 4488 3538 4522 3572
rect 4556 3538 4590 3572
rect 4624 3538 4658 3572
rect 4848 3538 4882 3572
rect 4916 3538 4950 3572
rect 4984 3538 5018 3572
rect 5052 3538 5086 3572
rect 5120 3538 5154 3572
rect 1386 3444 1420 3478
rect 1470 3444 1504 3478
rect 1554 3444 1588 3478
rect 1638 3444 1672 3478
rect 1722 3444 1756 3478
rect 1806 3444 1840 3478
rect 1890 3444 1924 3478
rect 1974 3444 2008 3478
rect 2058 3444 2092 3478
rect 2148 3444 2182 3478
rect 2694 3454 2728 3488
rect 2778 3454 2812 3488
rect 2862 3454 2896 3488
rect 2946 3454 2980 3488
rect 3030 3454 3064 3488
rect 3114 3454 3148 3488
rect 3198 3454 3232 3488
rect 3282 3454 3316 3488
rect 932 2740 968 2776
rect 1166 2740 1202 2776
rect 3772 2092 3810 2130
rect 3848 2092 3886 2130
rect 3924 2092 3962 2130
rect 4000 2092 4038 2130
rect 4512 2092 4546 2126
rect 4580 2092 4614 2126
rect 4648 2092 4682 2126
rect 4716 2092 4750 2126
rect 4784 2092 4818 2126
<< poly >>
rect 1034 4848 1154 4978
rect 1034 4798 1064 4848
rect 1114 4798 1154 4848
rect 1034 4758 1154 4798
rect 1034 4708 1064 4758
rect 1114 4708 1154 4758
rect 1034 4668 1154 4708
rect 1034 4618 1064 4668
rect 1114 4618 1154 4668
rect 1034 4568 1154 4618
rect 1034 4518 1064 4568
rect 1114 4518 1154 4568
rect 1034 4478 1154 4518
rect 1034 4428 1064 4478
rect 1114 4428 1154 4478
rect 1034 4388 1154 4428
rect 1034 4338 1064 4388
rect 1114 4338 1154 4388
rect 1034 4198 1154 4338
rect 4834 4838 4944 4978
rect 4834 4788 4874 4838
rect 4924 4788 4944 4838
rect 4834 4748 4944 4788
rect 4834 4698 4874 4748
rect 4924 4698 4944 4748
rect 4834 4658 4944 4698
rect 4834 4608 4874 4658
rect 4924 4628 4944 4658
rect 4924 4608 4954 4628
rect 4834 4558 4954 4608
rect 4834 4508 4874 4558
rect 4924 4548 4954 4558
rect 4924 4508 4944 4548
rect 4834 4468 4944 4508
rect 4834 4418 4874 4468
rect 4924 4418 4944 4468
rect 4834 4378 4944 4418
rect 4834 4328 4874 4378
rect 4924 4328 4944 4378
rect 4834 4198 4944 4328
rect 3906 3488 4032 3518
rect 3810 3462 3840 3488
rect 3906 3462 3936 3488
rect 4002 3462 4032 3488
rect 4302 3496 4568 3512
rect 4302 3462 4312 3496
rect 4346 3482 4568 3496
rect 4346 3462 4376 3482
rect 1418 3382 1448 3408
rect 1514 3382 1544 3408
rect 1610 3382 1640 3408
rect 1706 3382 1736 3408
rect 1802 3382 1832 3408
rect 1898 3382 1928 3408
rect 1994 3382 2024 3408
rect 2090 3382 2120 3408
rect 2550 3332 2580 3358
rect 2646 3332 2676 3358
rect 2872 3332 2902 3358
rect 2968 3332 2998 3358
rect 3064 3332 3094 3358
rect 3160 3332 3190 3358
rect 3386 3332 3416 3358
rect 3482 3332 3512 3358
rect 1418 3256 1448 3282
rect 1514 3256 1544 3282
rect 1610 3256 1640 3282
rect 1706 3256 1736 3282
rect 1802 3256 1832 3282
rect 1898 3256 1928 3282
rect 1994 3256 2024 3282
rect 2090 3256 2120 3282
rect 1418 3224 2120 3256
rect 1740 3182 1798 3224
rect 1260 3172 1798 3182
rect 1260 3138 1276 3172
rect 1310 3146 1798 3172
rect 1310 3138 1326 3146
rect 1260 3124 1326 3138
rect 1926 3094 1998 3104
rect 1926 3054 1942 3094
rect 1982 3054 1998 3094
rect 1534 3044 1606 3054
rect 1926 3044 1998 3054
rect 2374 3084 2442 3094
rect 2374 3048 2390 3084
rect 2426 3048 2442 3084
rect 1534 3004 1550 3044
rect 1590 3004 1606 3044
rect 1534 2994 1606 3004
rect 1558 2924 1596 2994
rect 1942 2924 1980 3044
rect 2374 3010 2442 3048
rect 2374 2974 2390 3010
rect 2426 2974 2442 3010
rect 2374 2936 2442 2974
rect 1418 2894 1736 2924
rect 1418 2868 1448 2894
rect 1514 2868 1544 2894
rect 1610 2868 1640 2894
rect 1706 2868 1736 2894
rect 1802 2894 2120 2924
rect 1802 2868 1832 2894
rect 1898 2868 1928 2894
rect 1994 2868 2024 2894
rect 2090 2868 2120 2894
rect 2374 2900 2390 2936
rect 2426 2916 2442 2936
rect 4302 3446 4376 3462
rect 4346 3414 4376 3446
rect 4442 3414 4472 3440
rect 4538 3414 4568 3482
rect 4798 3496 5064 3512
rect 4798 3462 4808 3496
rect 4842 3482 5064 3496
rect 4842 3462 4872 3482
rect 4798 3446 4872 3462
rect 4634 3414 4664 3440
rect 4842 3414 4872 3446
rect 4938 3414 4968 3440
rect 5034 3414 5064 3482
rect 5130 3414 5160 3440
rect 3810 3236 3840 3262
rect 3798 3212 3840 3236
rect 3670 3174 3744 3190
rect 3670 3140 3684 3174
rect 3720 3140 3744 3174
rect 3670 3122 3744 3140
rect 3798 3122 3830 3212
rect 3906 3180 3936 3262
rect 4002 3236 4032 3262
rect 3670 3102 3830 3122
rect 3872 3163 3936 3180
rect 3872 3129 3882 3163
rect 3916 3129 3936 3163
rect 4346 3140 4376 3254
rect 4442 3222 4472 3254
rect 4538 3228 4568 3254
rect 4418 3206 4472 3222
rect 4418 3172 4428 3206
rect 4462 3186 4472 3206
rect 4634 3186 4664 3254
rect 4462 3172 4664 3186
rect 4418 3156 4664 3172
rect 3872 3112 3936 3129
rect 3670 3068 3684 3102
rect 3720 3086 3830 3102
rect 3720 3068 3744 3086
rect 3670 3052 3744 3068
rect 3798 3084 3830 3086
rect 3798 3060 3840 3084
rect 3810 3036 3840 3060
rect 3906 3082 3936 3112
rect 4238 3108 4376 3140
rect 3906 3052 4032 3082
rect 3906 3036 3936 3052
rect 4002 3036 4032 3052
rect 4238 2948 4268 3108
rect 4346 3084 4376 3108
rect 4442 3084 4472 3156
rect 4842 3084 4872 3254
rect 4938 3222 4968 3254
rect 5034 3228 5064 3254
rect 4914 3206 4968 3222
rect 4914 3172 4924 3206
rect 4958 3186 4968 3206
rect 5130 3186 5160 3254
rect 4958 3172 5160 3186
rect 4914 3156 5160 3172
rect 4938 3084 4968 3156
rect 4346 2974 4376 3000
rect 4442 2974 4472 3000
rect 4842 2974 4872 3000
rect 4938 2974 4968 3000
rect 2550 2916 2580 2932
rect 2646 2916 2676 2932
rect 2426 2900 2676 2916
rect 2374 2886 2676 2900
rect 2872 2916 2902 2932
rect 2968 2916 2998 2932
rect 2872 2886 2998 2916
rect 862 2600 908 2630
rect 996 2600 1022 2630
rect 1096 2600 1142 2630
rect 1230 2600 1256 2630
rect 862 2538 892 2600
rect 1096 2538 1126 2600
rect 862 2508 908 2538
rect 996 2508 1022 2538
rect 1096 2508 1142 2538
rect 1230 2508 1256 2538
rect 862 2424 892 2508
rect 1096 2424 1126 2508
rect 2964 2820 2998 2886
rect 2932 2810 2998 2820
rect 2932 2776 2948 2810
rect 2982 2776 2998 2810
rect 2932 2766 2998 2776
rect 2872 2602 2902 2628
rect 2968 2602 2998 2766
rect 3064 2916 3094 2932
rect 3160 2916 3190 2932
rect 3064 2886 3190 2916
rect 3386 2916 3416 2932
rect 3482 2916 3512 2932
rect 3386 2886 3512 2916
rect 3810 2910 3840 2936
rect 3906 2910 3936 2936
rect 4002 2910 4032 2936
rect 4238 2930 4312 2948
rect 3064 2752 3098 2886
rect 3064 2742 3324 2752
rect 3064 2708 3082 2742
rect 3116 2708 3324 2742
rect 3478 2710 3512 2886
rect 4238 2896 4268 2930
rect 4302 2896 4312 2930
rect 4238 2880 4312 2896
rect 3810 2724 3840 2750
rect 3906 2724 3936 2750
rect 4002 2724 4032 2750
rect 3064 2698 3324 2708
rect 3064 2602 3094 2698
rect 3160 2602 3190 2628
rect 1418 2440 1448 2468
rect 1514 2440 1544 2468
rect 1610 2440 1640 2468
rect 1706 2440 1736 2468
rect 1802 2440 1832 2468
rect 1898 2440 1928 2468
rect 1994 2440 2024 2468
rect 2090 2440 2120 2468
rect 820 2408 892 2424
rect 820 2374 836 2408
rect 870 2374 892 2408
rect 820 2358 892 2374
rect 1054 2408 1126 2424
rect 1054 2374 1070 2408
rect 1104 2374 1126 2408
rect 1054 2358 1126 2374
rect 862 2288 892 2358
rect 1096 2288 1126 2358
rect 1268 2374 1334 2384
rect 1268 2340 1284 2374
rect 1318 2364 1334 2374
rect 1318 2340 2120 2364
rect 1268 2334 2120 2340
rect 1268 2330 1334 2334
rect 1418 2308 1448 2334
rect 1514 2308 1544 2334
rect 1610 2308 1640 2334
rect 1706 2308 1736 2334
rect 1802 2308 1832 2334
rect 1898 2308 1928 2334
rect 1994 2308 2024 2334
rect 2090 2308 2120 2334
rect 862 2258 908 2288
rect 992 2258 1018 2288
rect 1096 2258 1142 2288
rect 1226 2258 1252 2288
rect 1418 2182 1448 2208
rect 1514 2182 1544 2208
rect 1610 2182 1640 2208
rect 1706 2182 1736 2208
rect 1802 2182 1832 2208
rect 1898 2182 1928 2208
rect 1994 2182 2024 2208
rect 2090 2182 2120 2208
rect 3268 2582 3324 2698
rect 3382 2694 3512 2710
rect 3382 2658 3392 2694
rect 3428 2658 3466 2694
rect 3502 2658 3512 2694
rect 3382 2642 3512 2658
rect 4506 2664 4536 2690
rect 4602 2664 4632 2690
rect 3810 2600 3840 2624
rect 3268 2574 3744 2582
rect 3798 2576 3840 2600
rect 3906 2608 3936 2624
rect 4002 2608 4032 2624
rect 3906 2578 4032 2608
rect 3798 2574 3830 2576
rect 3268 2538 3830 2574
rect 3906 2548 3936 2578
rect 3268 2526 3744 2538
rect 3798 2448 3830 2538
rect 3872 2531 3936 2548
rect 3872 2497 3882 2531
rect 3916 2497 3936 2531
rect 3872 2480 3936 2497
rect 3798 2424 3840 2448
rect 3810 2398 3840 2424
rect 3906 2398 3936 2480
rect 4002 2398 4032 2424
rect 4506 2410 4536 2580
rect 4602 2508 4632 2580
rect 4578 2492 4824 2508
rect 4578 2458 4588 2492
rect 4622 2478 4824 2492
rect 4622 2458 4632 2478
rect 4578 2442 4632 2458
rect 4602 2410 4632 2442
rect 4698 2410 4728 2436
rect 4794 2410 4824 2478
rect 2872 2134 2902 2202
rect 2968 2176 2998 2202
rect 3064 2176 3094 2202
rect 3160 2134 3190 2202
rect 4506 2218 4536 2250
rect 4602 2224 4632 2250
rect 4462 2202 4536 2218
rect 3810 2172 3840 2198
rect 3906 2172 3936 2198
rect 4002 2172 4032 2198
rect 3906 2142 4032 2172
rect 4462 2168 4472 2202
rect 4506 2182 4536 2202
rect 4698 2182 4728 2250
rect 4794 2224 4824 2250
rect 4506 2168 4728 2182
rect 4462 2152 4728 2168
rect 2636 2124 3190 2134
rect 2636 2090 2652 2124
rect 2686 2090 2730 2124
rect 2764 2104 3190 2124
rect 2764 2090 2780 2104
rect 2636 2080 2780 2090
rect 1034 1258 1154 1388
rect 1034 1208 1064 1258
rect 1114 1208 1154 1258
rect 1034 1168 1154 1208
rect 1034 1118 1064 1168
rect 1114 1118 1154 1168
rect 1034 1078 1154 1118
rect 1034 1028 1064 1078
rect 1114 1028 1154 1078
rect 1034 978 1154 1028
rect 1034 928 1064 978
rect 1114 928 1154 978
rect 1034 888 1154 928
rect 1034 838 1064 888
rect 1114 838 1154 888
rect 1034 798 1154 838
rect 1034 748 1064 798
rect 1114 748 1154 798
rect 1034 608 1154 748
rect 4834 1248 4944 1388
rect 4834 1198 4874 1248
rect 4924 1198 4944 1248
rect 4834 1158 4944 1198
rect 4834 1108 4874 1158
rect 4924 1108 4944 1158
rect 4834 1068 4944 1108
rect 4834 1018 4874 1068
rect 4924 1038 4944 1068
rect 4924 1018 4954 1038
rect 4834 968 4954 1018
rect 4834 918 4874 968
rect 4924 958 4954 968
rect 4924 918 4944 958
rect 4834 878 4944 918
rect 4834 828 4874 878
rect 4924 828 4944 878
rect 4834 788 4944 828
rect 4834 738 4874 788
rect 4924 738 4944 788
rect 4834 608 4944 738
<< polycont >>
rect 1064 4798 1114 4848
rect 1064 4708 1114 4758
rect 1064 4618 1114 4668
rect 1064 4518 1114 4568
rect 1064 4428 1114 4478
rect 1064 4338 1114 4388
rect 4874 4788 4924 4838
rect 4874 4698 4924 4748
rect 4874 4608 4924 4658
rect 4874 4508 4924 4558
rect 4874 4418 4924 4468
rect 4874 4328 4924 4378
rect 4312 3462 4346 3496
rect 1276 3138 1310 3172
rect 1942 3054 1982 3094
rect 2390 3048 2426 3084
rect 1550 3004 1590 3044
rect 2390 2974 2426 3010
rect 2390 2900 2426 2936
rect 4808 3462 4842 3496
rect 3684 3140 3720 3174
rect 3882 3129 3916 3163
rect 4428 3172 4462 3206
rect 3684 3068 3720 3102
rect 4924 3172 4958 3206
rect 2948 2776 2982 2810
rect 3082 2708 3116 2742
rect 4268 2896 4302 2930
rect 836 2374 870 2408
rect 1070 2374 1104 2408
rect 1284 2340 1318 2374
rect 3392 2658 3428 2694
rect 3466 2658 3502 2694
rect 3882 2497 3916 2531
rect 4588 2458 4622 2492
rect 4472 2168 4506 2202
rect 2652 2090 2686 2124
rect 2730 2090 2764 2124
rect 1064 1208 1114 1258
rect 1064 1118 1114 1168
rect 1064 1028 1114 1078
rect 1064 928 1114 978
rect 1064 838 1114 888
rect 1064 748 1114 798
rect 4874 1198 4924 1248
rect 4874 1108 4924 1158
rect 4874 1018 4924 1068
rect 4874 918 4924 968
rect 4874 828 4924 878
rect 4874 738 4924 788
<< locali >>
rect 588 5540 5466 5596
rect 588 5466 1012 5540
rect 1086 5466 1560 5540
rect 1634 5466 2108 5540
rect 2182 5466 2656 5540
rect 2730 5466 3204 5540
rect 3278 5466 3734 5540
rect 3808 5466 4282 5540
rect 4356 5466 4832 5540
rect 4906 5466 5466 5540
rect 588 5398 5466 5466
rect 588 5348 646 5398
rect 720 5348 824 5398
rect 588 4948 624 5348
rect 754 4948 824 5348
rect 1474 5298 1934 5398
rect 4054 5298 4514 5398
rect 5268 5328 5466 5398
rect 588 4924 824 4948
rect 588 4850 646 4924
rect 720 4908 824 4924
rect 904 5278 5084 5298
rect 904 5228 1504 5278
rect 1904 5228 4084 5278
rect 4484 5228 5084 5278
rect 904 5218 5084 5228
rect 720 4850 786 4908
rect 588 4808 786 4850
rect 588 4368 608 4808
rect 744 4368 786 4808
rect 588 4248 786 4368
rect 588 3818 608 4248
rect 764 3818 786 4248
rect 904 3958 984 5218
rect 1474 5208 1934 5218
rect 4054 5208 4514 5218
rect 1144 4998 1164 5098
rect 1284 4998 1324 5098
rect 1444 4998 1484 5098
rect 1604 4998 1644 5098
rect 1764 4998 1804 5098
rect 1924 4998 1964 5098
rect 2084 4998 2124 5098
rect 2244 4998 3744 5098
rect 3864 4998 3904 5098
rect 4024 4998 4064 5098
rect 4184 4998 4224 5098
rect 4344 4998 4384 5098
rect 4504 4998 4544 5098
rect 4664 4998 4704 5098
rect 4824 4998 4844 5098
rect 1144 4978 4844 4998
rect 1064 4898 1624 4938
rect 1064 4848 1174 4898
rect 1664 4858 1734 4978
rect 1114 4798 1174 4848
rect 1214 4818 1734 4858
rect 1064 4778 1174 4798
rect 1064 4758 1624 4778
rect 1134 4738 1624 4758
rect 1134 4708 1174 4738
rect 1064 4668 1174 4708
rect 1664 4698 1734 4818
rect 1134 4618 1174 4668
rect 1214 4658 1734 4698
rect 1774 4628 1814 4938
rect 1854 4678 1894 4978
rect 1934 4628 1974 4938
rect 2014 4678 2054 4978
rect 2094 4628 2134 4938
rect 2174 4678 2214 4978
rect 2254 4628 2294 4938
rect 2334 4678 2374 4978
rect 2414 4628 2454 4938
rect 2494 4678 2534 4978
rect 2574 4628 2614 4938
rect 2654 4678 2694 4978
rect 2734 4628 2774 4938
rect 2814 4678 2854 4978
rect 2894 4628 2934 4938
rect 2974 4678 3014 4978
rect 3054 4628 3094 4938
rect 3134 4678 3174 4978
rect 3214 4628 3254 4938
rect 3294 4678 3334 4978
rect 3374 4628 3414 4938
rect 3454 4678 3494 4978
rect 3534 4628 3574 4938
rect 3614 4678 3654 4978
rect 3694 4628 3734 4938
rect 3774 4678 3814 4978
rect 3854 4628 3894 4938
rect 3934 4678 3974 4978
rect 4014 4628 4054 4938
rect 4094 4678 4134 4978
rect 4174 4628 4214 4938
rect 4254 4858 4324 4978
rect 4364 4898 4924 4938
rect 4254 4818 4774 4858
rect 4814 4838 4924 4898
rect 4254 4698 4324 4818
rect 4814 4788 4874 4838
rect 4814 4778 4924 4788
rect 4364 4748 4924 4778
rect 4364 4738 4854 4748
rect 4814 4698 4854 4738
rect 4254 4658 4764 4698
rect 4814 4658 4924 4698
rect 1774 4618 4214 4628
rect 4814 4618 4854 4658
rect 1064 4608 4854 4618
rect 1064 4568 4924 4608
rect 1134 4558 4924 4568
rect 1134 4518 1174 4558
rect 1774 4548 4214 4558
rect 1064 4478 1174 4518
rect 1214 4478 1734 4518
rect 1134 4438 1174 4478
rect 1134 4428 1624 4438
rect 1064 4398 1624 4428
rect 1064 4388 1174 4398
rect 1114 4338 1174 4388
rect 1664 4358 1734 4478
rect 1064 4278 1174 4338
rect 1214 4318 1734 4358
rect 1064 4238 1624 4278
rect 1664 4198 1734 4318
rect 1774 4238 1814 4548
rect 1854 4198 1894 4498
rect 1934 4238 1974 4548
rect 2014 4198 2054 4498
rect 2094 4238 2134 4548
rect 2174 4198 2214 4498
rect 2254 4238 2294 4548
rect 2334 4198 2374 4498
rect 2414 4238 2454 4548
rect 2494 4198 2534 4498
rect 2574 4238 2614 4548
rect 2654 4198 2694 4498
rect 2734 4238 2774 4548
rect 2814 4198 2854 4498
rect 2894 4248 2934 4548
rect 2974 4198 3014 4498
rect 3054 4248 3094 4548
rect 3134 4198 3174 4498
rect 3214 4238 3254 4548
rect 3294 4198 3334 4498
rect 3374 4238 3414 4548
rect 3454 4198 3494 4498
rect 3534 4238 3574 4548
rect 3614 4198 3654 4498
rect 3694 4238 3734 4548
rect 3774 4198 3814 4498
rect 3854 4238 3894 4548
rect 3934 4198 3974 4498
rect 4014 4238 4054 4548
rect 4094 4198 4134 4498
rect 4174 4238 4214 4548
rect 4254 4478 4764 4518
rect 4814 4508 4854 4558
rect 4254 4358 4324 4478
rect 4814 4468 4924 4508
rect 4814 4438 4854 4468
rect 4364 4418 4854 4438
rect 4364 4398 4924 4418
rect 4814 4378 4924 4398
rect 4254 4318 4774 4358
rect 4814 4328 4874 4378
rect 4254 4198 4324 4318
rect 4814 4278 4924 4328
rect 4364 4238 4924 4278
rect 1144 4178 4844 4198
rect 1144 4078 1164 4178
rect 1284 4078 1324 4178
rect 1444 4078 1484 4178
rect 1604 4078 1644 4178
rect 1764 4078 1804 4178
rect 1924 4078 1964 4178
rect 2084 4078 2124 4178
rect 2244 4078 3744 4178
rect 3864 4078 3904 4178
rect 4024 4078 4064 4178
rect 4184 4078 4224 4178
rect 4344 4078 4384 4178
rect 4504 4078 4544 4178
rect 4664 4078 4704 4178
rect 4824 4078 4844 4178
rect 1474 3958 1934 3968
rect 4054 3958 4514 3968
rect 5004 3958 5084 5218
rect 904 3948 5084 3958
rect 904 3898 1504 3948
rect 1904 3898 4084 3948
rect 4484 3898 5084 3948
rect 904 3878 5084 3898
rect 5268 5254 5328 5328
rect 5402 5254 5466 5328
rect 5268 4852 5466 5254
rect 5268 4778 5328 4852
rect 5402 4778 5466 4852
rect 5268 4378 5466 4778
rect 5268 4304 5328 4378
rect 5402 4304 5466 4378
rect 5268 3904 5466 4304
rect 588 3290 786 3818
rect 1474 3798 1934 3878
rect 4054 3798 4514 3878
rect 5268 3830 5326 3904
rect 5400 3830 5466 3904
rect 3678 3608 4226 3628
rect 3678 3572 3772 3608
rect 3808 3572 3848 3608
rect 3884 3572 3924 3608
rect 3960 3572 4000 3608
rect 4036 3572 4076 3608
rect 4112 3572 4152 3608
rect 4188 3572 4226 3608
rect 3678 3568 4226 3572
rect 3678 3530 3772 3568
rect 3810 3530 3848 3568
rect 3886 3530 3924 3568
rect 3962 3530 4000 3568
rect 4038 3530 4226 3568
rect 4336 3538 4352 3572
rect 4386 3538 4420 3572
rect 4454 3538 4488 3572
rect 4522 3538 4556 3572
rect 4590 3538 4624 3572
rect 4658 3538 4848 3572
rect 4882 3538 4916 3572
rect 4950 3538 4984 3572
rect 5018 3538 5052 3572
rect 5086 3538 5120 3572
rect 5154 3538 5182 3572
rect 2656 3488 3380 3496
rect 588 3216 646 3290
rect 720 3216 786 3290
rect 588 2764 786 3216
rect 1140 3480 2212 3486
rect 1140 3444 1152 3480
rect 1186 3444 1230 3480
rect 1264 3444 1302 3480
rect 1336 3478 2212 3480
rect 1336 3444 1386 3478
rect 1420 3444 1470 3478
rect 1504 3444 1554 3478
rect 1588 3444 1638 3478
rect 1672 3444 1722 3478
rect 1756 3444 1806 3478
rect 1840 3444 1890 3478
rect 1924 3444 1974 3478
rect 2008 3444 2058 3478
rect 2092 3444 2148 3478
rect 2182 3444 2212 3478
rect 2656 3454 2694 3488
rect 2728 3454 2778 3488
rect 2812 3454 2862 3488
rect 2896 3454 2946 3488
rect 2980 3454 3030 3488
rect 3064 3454 3114 3488
rect 3148 3454 3198 3488
rect 3232 3454 3282 3488
rect 3316 3454 3380 3488
rect 2656 3448 3380 3454
rect 3760 3450 3794 3466
rect 1140 3438 2212 3444
rect 1140 2812 1226 3438
rect 1368 3420 2170 3438
rect 1368 3370 1402 3420
rect 1368 3278 1402 3294
rect 1464 3370 1498 3386
rect 1464 3218 1498 3294
rect 1560 3370 1594 3420
rect 1560 3278 1594 3294
rect 1656 3370 1690 3386
rect 1656 3218 1690 3294
rect 1752 3370 1786 3420
rect 1752 3278 1786 3294
rect 1848 3370 1882 3386
rect 1464 3184 1690 3218
rect 1848 3218 1882 3294
rect 1944 3370 1978 3420
rect 1944 3278 1978 3294
rect 2040 3370 2074 3386
rect 2040 3218 2074 3294
rect 2136 3370 2170 3420
rect 2136 3278 2170 3294
rect 2264 3428 2454 3448
rect 2264 3278 2284 3428
rect 2434 3278 2454 3428
rect 2992 3414 3082 3448
rect 2264 3258 2454 3278
rect 2500 3370 2726 3404
rect 2500 3320 2534 3370
rect 1848 3184 2074 3218
rect 1260 3172 1326 3182
rect 1260 3138 1276 3172
rect 1310 3138 1326 3172
rect 1260 3124 1326 3138
rect 588 2690 638 2764
rect 712 2690 786 2764
rect 588 2290 786 2690
rect 820 2778 932 2812
rect 968 2778 1166 2812
rect 1202 2778 1226 2812
rect 820 2776 1226 2778
rect 820 2772 932 2776
rect 820 2588 856 2772
rect 908 2740 932 2772
rect 968 2772 1166 2776
rect 968 2740 992 2772
rect 908 2680 996 2686
rect 904 2678 1000 2680
rect 904 2644 920 2678
rect 980 2644 1000 2678
rect 904 2642 1000 2644
rect 1046 2588 1090 2772
rect 1142 2740 1166 2772
rect 1202 2740 1226 2776
rect 1142 2680 1230 2686
rect 1138 2678 1234 2680
rect 1138 2644 1154 2678
rect 1214 2644 1234 2678
rect 1138 2642 1234 2644
rect 820 2586 1000 2588
rect 820 2552 920 2586
rect 980 2552 1000 2586
rect 820 2550 1000 2552
rect 1046 2586 1234 2588
rect 1046 2552 1154 2586
rect 1214 2552 1234 2586
rect 1046 2550 1234 2552
rect 904 2462 920 2496
rect 980 2462 1000 2496
rect 1138 2462 1154 2496
rect 1214 2462 1234 2496
rect 908 2450 996 2462
rect 1142 2450 1230 2462
rect 820 2408 874 2424
rect 820 2374 836 2408
rect 870 2374 874 2408
rect 820 2358 874 2374
rect 908 2414 992 2450
rect 1054 2414 1108 2424
rect 908 2408 1108 2414
rect 908 2374 1070 2408
rect 1104 2374 1108 2408
rect 908 2368 1108 2374
rect 908 2334 992 2368
rect 1054 2358 1108 2368
rect 1142 2414 1226 2450
rect 1280 2414 1326 3124
rect 1464 2960 1498 3184
rect 1534 3044 1606 3054
rect 1534 3004 1550 3044
rect 1590 3004 1606 3044
rect 1534 2994 1606 3004
rect 1642 3014 1690 3020
rect 1642 2978 1648 3014
rect 1684 2978 1690 3014
rect 1642 2960 1690 2978
rect 1464 2926 1690 2960
rect 1142 2384 1326 2414
rect 1368 2856 1402 2872
rect 1368 2430 1402 2480
rect 1464 2856 1498 2926
rect 1464 2464 1498 2480
rect 1560 2856 1594 2872
rect 1560 2430 1594 2480
rect 1656 2856 1690 2926
rect 1848 2962 1882 3184
rect 1926 3094 1998 3104
rect 1926 3054 1942 3094
rect 1982 3054 1998 3094
rect 1926 3044 1998 3054
rect 2370 3084 2446 3258
rect 2370 3048 2390 3084
rect 2426 3048 2446 3084
rect 2370 3010 2446 3048
rect 2370 2974 2390 3010
rect 2426 2974 2446 3010
rect 1848 2928 2324 2962
rect 1656 2464 1690 2480
rect 1752 2856 1786 2872
rect 1752 2430 1786 2480
rect 1848 2856 1882 2928
rect 1848 2464 1882 2480
rect 1944 2856 1978 2872
rect 1944 2430 1978 2480
rect 2040 2856 2074 2928
rect 2040 2464 2074 2480
rect 2136 2856 2170 2872
rect 2248 2838 2324 2928
rect 2370 2936 2446 2974
rect 2370 2900 2390 2936
rect 2426 2900 2446 2936
rect 2370 2872 2446 2900
rect 2248 2826 2446 2838
rect 2248 2790 2390 2826
rect 2426 2790 2446 2826
rect 2500 2810 2534 2944
rect 2596 3320 2630 3336
rect 2596 2878 2630 2944
rect 2692 3320 2726 3370
rect 2692 2928 2726 2944
rect 2822 3380 3240 3414
rect 2822 3320 2856 3380
rect 2822 2928 2856 2944
rect 2918 3320 2952 3336
rect 2918 2878 2952 2944
rect 3014 3320 3048 3380
rect 3014 2928 3048 2944
rect 3110 3320 3144 3336
rect 2596 2844 2952 2878
rect 3110 2878 3144 2944
rect 3206 3320 3240 3380
rect 3206 2928 3240 2944
rect 3336 3370 3562 3404
rect 3336 3320 3370 3370
rect 3336 2928 3370 2944
rect 3432 3320 3466 3336
rect 3432 2878 3466 2944
rect 3110 2844 3466 2878
rect 3528 3320 3562 3370
rect 3562 3174 3726 3190
rect 3562 3140 3684 3174
rect 3720 3140 3726 3174
rect 3562 3102 3726 3140
rect 3562 3068 3684 3102
rect 3720 3068 3726 3102
rect 3562 3052 3726 3068
rect 3760 3180 3794 3274
rect 3856 3450 3890 3530
rect 3856 3258 3890 3274
rect 3952 3450 3986 3466
rect 3760 3163 3918 3180
rect 3760 3129 3882 3163
rect 3916 3129 3918 3163
rect 3760 3112 3918 3129
rect 3952 3144 3986 3274
rect 4048 3450 4082 3530
rect 4048 3258 4082 3274
rect 4060 3144 4120 3154
rect 3952 3142 4134 3144
rect 3528 2810 3562 2944
rect 3760 3024 3794 3112
rect 3952 3106 4066 3142
rect 4102 3106 4134 3142
rect 3760 2932 3794 2948
rect 3856 3024 3890 3040
rect 3856 2882 3890 2948
rect 3952 3024 3986 3106
rect 4060 3094 4120 3106
rect 3952 2932 3986 2948
rect 4048 3024 4082 3040
rect 4048 2882 4082 2948
rect 3748 2864 3774 2882
rect 3612 2848 3774 2864
rect 3808 2848 3842 2882
rect 3876 2848 3910 2882
rect 3944 2848 3978 2882
rect 4012 2848 4046 2882
rect 4080 2848 4104 2882
rect 3612 2812 4104 2848
rect 2248 2750 2446 2790
rect 2484 2776 2896 2810
rect 2932 2776 2948 2810
rect 2982 2776 3574 2810
rect 3612 2796 3774 2812
rect 2248 2714 2390 2750
rect 2426 2714 2446 2750
rect 2248 2676 2446 2714
rect 2862 2742 2896 2776
rect 2862 2708 3082 2742
rect 3116 2708 3132 2742
rect 2248 2640 2390 2676
rect 2426 2640 2446 2676
rect 2248 2626 2446 2640
rect 2136 2430 2170 2480
rect 1368 2394 2170 2430
rect 1142 2374 1334 2384
rect 1142 2368 1284 2374
rect 1142 2334 1226 2368
rect 1268 2340 1284 2368
rect 1318 2340 1334 2374
rect 904 2300 920 2334
rect 980 2300 996 2334
rect 1138 2300 1154 2334
rect 1214 2300 1230 2334
rect 1268 2330 1334 2340
rect 908 2294 992 2300
rect 1142 2294 1226 2300
rect 1368 2296 1402 2394
rect 588 2216 638 2290
rect 712 2216 786 2290
rect 588 2156 786 2216
rect 904 2212 920 2246
rect 980 2212 996 2246
rect 1138 2212 1154 2246
rect 1214 2212 1230 2246
rect 588 2122 604 2156
rect 638 2122 676 2156
rect 710 2122 748 2156
rect 782 2122 786 2156
rect 588 2084 786 2122
rect 908 2146 992 2212
rect 908 2112 932 2146
rect 968 2112 992 2146
rect 908 2106 992 2112
rect 1142 2146 1226 2212
rect 1368 2204 1402 2220
rect 1464 2296 1498 2314
rect 1142 2112 1166 2146
rect 1202 2112 1226 2146
rect 1142 2106 1226 2112
rect 588 2050 604 2084
rect 638 2050 676 2084
rect 710 2050 748 2084
rect 782 2050 786 2084
rect 588 2012 786 2050
rect 1464 2062 1498 2220
rect 1560 2296 1594 2394
rect 1560 2204 1594 2220
rect 1656 2296 1690 2312
rect 1656 2062 1690 2220
rect 1752 2296 1786 2394
rect 1752 2204 1786 2220
rect 1848 2296 1882 2312
rect 1848 2062 1882 2220
rect 1944 2296 1978 2394
rect 1944 2204 1978 2220
rect 2040 2296 2074 2312
rect 2040 2062 2074 2220
rect 2136 2296 2170 2394
rect 2370 2368 2446 2626
rect 2822 2590 2856 2606
rect 2136 2204 2170 2220
rect 2364 2348 2554 2368
rect 2364 2198 2384 2348
rect 2534 2198 2554 2348
rect 2364 2178 2554 2198
rect 2636 2124 2780 2134
rect 2636 2090 2652 2124
rect 2686 2090 2730 2124
rect 2764 2090 2780 2124
rect 2822 2090 2856 2214
rect 2918 2590 2952 2708
rect 3176 2674 3210 2776
rect 3110 2640 3210 2674
rect 3386 2694 3508 2710
rect 3386 2658 3392 2694
rect 3428 2658 3466 2694
rect 3502 2658 3508 2694
rect 3386 2642 3508 2658
rect 2918 2198 2952 2214
rect 3014 2590 3048 2606
rect 3014 2090 3048 2214
rect 3110 2590 3144 2640
rect 3110 2198 3144 2214
rect 3206 2590 3240 2606
rect 3612 2470 3680 2796
rect 3748 2778 3774 2796
rect 3808 2778 3842 2812
rect 3876 2778 3910 2812
rect 3944 2778 3978 2812
rect 4012 2778 4046 2812
rect 4080 2778 4104 2812
rect 3206 2090 3240 2214
rect 3542 2402 3680 2470
rect 3760 2712 3794 2728
rect 3760 2548 3794 2636
rect 3856 2712 3890 2778
rect 3856 2620 3890 2636
rect 3952 2712 3986 2728
rect 3952 2554 3986 2636
rect 4048 2712 4082 2778
rect 4048 2620 4082 2636
rect 4064 2554 4124 2564
rect 3952 2552 4136 2554
rect 3760 2531 3918 2548
rect 3760 2497 3882 2531
rect 3916 2497 3918 2531
rect 3760 2480 3918 2497
rect 3952 2516 4070 2552
rect 4106 2516 4136 2552
rect 2636 2080 2780 2090
rect 1464 2048 2074 2062
rect 2816 2054 2840 2090
rect 2876 2054 2932 2090
rect 2968 2054 3024 2090
rect 3060 2054 3116 2090
rect 3152 2054 3208 2090
rect 3244 2054 3268 2090
rect 2816 2052 3268 2054
rect 3542 2052 3622 2402
rect 3760 2386 3794 2480
rect 3760 2194 3794 2210
rect 3856 2386 3890 2402
rect 3856 2130 3890 2210
rect 3952 2386 3986 2516
rect 4064 2504 4124 2516
rect 3952 2194 3986 2210
rect 4048 2386 4082 2402
rect 4048 2130 4082 2210
rect 4170 2130 4226 3530
rect 4296 3496 4362 3504
rect 4296 3462 4312 3496
rect 4346 3462 4362 3496
rect 4296 3452 4362 3462
rect 4296 3402 4330 3418
rect 4296 3072 4330 3266
rect 4392 3402 4426 3418
rect 4392 3250 4426 3266
rect 4488 3402 4522 3538
rect 4792 3498 4858 3504
rect 4792 3462 4808 3498
rect 4842 3462 4858 3498
rect 4792 3452 4858 3462
rect 4488 3250 4522 3266
rect 4584 3402 4618 3418
rect 4584 3250 4618 3266
rect 4680 3402 4714 3418
rect 4412 3206 4478 3214
rect 4412 3172 4428 3206
rect 4462 3172 4478 3206
rect 4412 3162 4478 3172
rect 4680 3156 4714 3266
rect 4792 3402 4826 3418
rect 4680 3150 4728 3156
rect 4680 3146 4688 3150
rect 4508 3116 4688 3146
rect 4722 3116 4728 3150
rect 4508 3108 4728 3116
rect 4508 3088 4542 3108
rect 4296 2996 4330 3012
rect 4392 3072 4426 3088
rect 4392 2948 4426 3012
rect 4488 3072 4542 3088
rect 4522 3012 4542 3072
rect 4488 2996 4542 3012
rect 4792 3072 4826 3266
rect 4888 3402 4922 3418
rect 4888 3250 4922 3266
rect 4984 3402 5018 3538
rect 4984 3250 5018 3266
rect 5080 3402 5114 3418
rect 5080 3250 5114 3266
rect 5176 3402 5210 3418
rect 4908 3206 4974 3214
rect 4908 3172 4924 3206
rect 4958 3172 4974 3206
rect 4908 3162 4974 3172
rect 5176 3146 5210 3266
rect 5268 3292 5466 3830
rect 5268 3218 5326 3292
rect 5400 3218 5466 3292
rect 5004 3140 5234 3146
rect 5004 3108 5112 3140
rect 5004 3088 5038 3108
rect 5100 3104 5112 3108
rect 5148 3104 5186 3140
rect 5222 3104 5234 3140
rect 5100 3098 5234 3104
rect 4792 2996 4826 3012
rect 4888 3072 4922 3088
rect 4888 2948 4922 3012
rect 4984 3072 5038 3088
rect 5018 3012 5038 3072
rect 4984 2996 5038 3012
rect 5268 2948 5466 3218
rect 4366 2946 5466 2948
rect 4260 2930 4308 2946
rect 4260 2896 4268 2930
rect 4302 2896 4308 2930
rect 4366 2912 4392 2946
rect 4426 2912 4888 2946
rect 4922 2912 5466 2946
rect 4366 2896 5466 2912
rect 4260 2564 4308 2896
rect 4260 2528 4266 2564
rect 4302 2528 4308 2564
rect 4260 2212 4308 2528
rect 4342 2840 4390 2852
rect 4342 2804 4348 2840
rect 4384 2804 4390 2840
rect 4342 2504 4390 2804
rect 4528 2752 4614 2896
rect 4528 2718 4552 2752
rect 4586 2718 4614 2752
rect 5268 2818 5466 2896
rect 5268 2744 5326 2818
rect 5400 2744 5466 2818
rect 4342 2468 4348 2504
rect 4384 2468 4390 2504
rect 4342 2456 4390 2468
rect 4456 2652 4490 2668
rect 4456 2398 4490 2592
rect 4552 2652 4586 2718
rect 4552 2576 4586 2592
rect 4648 2652 4702 2668
rect 4682 2592 4702 2652
rect 4648 2576 4702 2592
rect 4668 2556 4702 2576
rect 4668 2550 5074 2556
rect 4668 2518 4950 2550
rect 4572 2492 4638 2502
rect 4572 2458 4588 2492
rect 4622 2458 4638 2492
rect 4572 2450 4638 2458
rect 4456 2246 4490 2262
rect 4552 2398 4586 2414
rect 4552 2246 4586 2262
rect 4648 2398 4682 2414
rect 4260 2202 4522 2212
rect 4260 2168 4472 2202
rect 4506 2168 4522 2202
rect 4260 2160 4522 2168
rect 3680 2092 3772 2130
rect 3810 2092 3848 2130
rect 3886 2092 3924 2130
rect 3962 2092 4000 2130
rect 4038 2126 4226 2130
rect 4648 2126 4682 2262
rect 4744 2398 4778 2414
rect 4744 2246 4778 2262
rect 4840 2398 4874 2518
rect 4938 2514 4950 2518
rect 4986 2514 5026 2550
rect 5062 2514 5074 2550
rect 4938 2508 5074 2514
rect 4840 2246 4874 2262
rect 5268 2344 5466 2744
rect 5268 2270 5326 2344
rect 5400 2270 5466 2344
rect 5268 2156 5466 2270
rect 4038 2092 4512 2126
rect 4546 2092 4580 2126
rect 4614 2092 4648 2126
rect 4682 2092 4716 2126
rect 4750 2092 4784 2126
rect 4818 2092 4846 2126
rect 5268 2122 5282 2156
rect 5316 2122 5354 2156
rect 5388 2122 5426 2156
rect 5460 2122 5466 2156
rect 5268 2084 5466 2122
rect 588 1978 604 2012
rect 638 1978 676 2012
rect 710 1978 748 2012
rect 782 1978 786 2012
rect 1350 2046 2168 2048
rect 1350 2010 1374 2046
rect 1410 2010 1492 2046
rect 1528 2010 1610 2046
rect 1646 2010 1728 2046
rect 1764 2010 1846 2046
rect 1882 2010 1964 2046
rect 2000 2010 2082 2046
rect 2118 2010 2168 2046
rect 1350 2006 2168 2010
rect 3542 2034 4514 2052
rect 3542 2032 3624 2034
rect 588 1940 786 1978
rect 588 1906 604 1940
rect 638 1906 676 1940
rect 710 1906 748 1940
rect 782 1906 786 1940
rect 588 1868 786 1906
rect 588 1834 602 1868
rect 636 1834 674 1868
rect 708 1834 746 1868
rect 780 1834 786 1868
rect 588 1768 786 1834
rect 588 1338 606 1768
rect 764 1338 786 1768
rect 1474 1708 1934 2006
rect 3542 1996 3550 2032
rect 3586 1998 3624 2032
rect 3660 1998 3704 2034
rect 3740 1998 3784 2034
rect 3820 1998 3864 2034
rect 3900 1998 4514 2034
rect 3586 1996 4514 1998
rect 3542 1982 4514 1996
rect 4054 1708 4514 1982
rect 5268 2050 5282 2084
rect 5316 2050 5354 2084
rect 5388 2050 5426 2084
rect 5460 2050 5466 2084
rect 5268 2012 5466 2050
rect 5268 1978 5282 2012
rect 5316 1978 5354 2012
rect 5388 1978 5426 2012
rect 5460 1978 5466 2012
rect 5268 1940 5466 1978
rect 5268 1906 5282 1940
rect 5316 1906 5354 1940
rect 5388 1906 5426 1940
rect 5460 1906 5466 1940
rect 5268 1868 5466 1906
rect 5268 1834 5282 1868
rect 5316 1834 5354 1868
rect 5388 1834 5426 1868
rect 5460 1834 5466 1868
rect 588 1218 786 1338
rect 588 778 614 1218
rect 744 778 786 1218
rect 588 690 786 778
rect 588 648 652 690
rect 726 648 786 690
rect 588 238 614 648
rect 774 238 786 648
rect 904 1688 5084 1708
rect 904 1638 1504 1688
rect 1904 1638 4084 1688
rect 4484 1638 5084 1688
rect 904 1628 5084 1638
rect 904 368 984 1628
rect 1474 1618 1934 1628
rect 4054 1618 4514 1628
rect 1144 1408 1164 1508
rect 1284 1408 1324 1508
rect 1444 1408 1484 1508
rect 1604 1408 1644 1508
rect 1764 1408 1804 1508
rect 1924 1408 1964 1508
rect 2084 1408 2124 1508
rect 2244 1408 3744 1508
rect 3864 1408 3904 1508
rect 4024 1408 4064 1508
rect 4184 1408 4224 1508
rect 4344 1408 4384 1508
rect 4504 1408 4544 1508
rect 4664 1408 4704 1508
rect 4824 1408 4844 1508
rect 1144 1388 4844 1408
rect 1064 1308 1624 1348
rect 1064 1258 1174 1308
rect 1664 1268 1734 1388
rect 1114 1208 1174 1258
rect 1214 1228 1734 1268
rect 1064 1188 1174 1208
rect 1064 1168 1624 1188
rect 1134 1148 1624 1168
rect 1134 1118 1174 1148
rect 1064 1078 1174 1118
rect 1664 1108 1734 1228
rect 1134 1028 1174 1078
rect 1214 1068 1734 1108
rect 1774 1038 1814 1348
rect 1854 1088 1894 1388
rect 1934 1038 1974 1348
rect 2014 1088 2054 1388
rect 2094 1038 2134 1348
rect 2174 1088 2214 1388
rect 2254 1038 2294 1348
rect 2334 1088 2374 1388
rect 2414 1038 2454 1348
rect 2494 1088 2534 1388
rect 2574 1038 2614 1348
rect 2654 1088 2694 1388
rect 2734 1038 2774 1348
rect 2814 1088 2854 1388
rect 2894 1038 2934 1348
rect 2974 1088 3014 1388
rect 3054 1038 3094 1348
rect 3134 1088 3174 1388
rect 3214 1038 3254 1348
rect 3294 1088 3334 1388
rect 3374 1038 3414 1348
rect 3454 1088 3494 1388
rect 3534 1038 3574 1348
rect 3614 1088 3654 1388
rect 3694 1038 3734 1348
rect 3774 1088 3814 1388
rect 3854 1038 3894 1348
rect 3934 1088 3974 1388
rect 4014 1038 4054 1348
rect 4094 1088 4134 1388
rect 4174 1038 4214 1348
rect 4254 1268 4324 1388
rect 4364 1308 4924 1348
rect 4254 1228 4774 1268
rect 4814 1248 4924 1308
rect 4254 1108 4324 1228
rect 4814 1198 4874 1248
rect 4814 1188 4924 1198
rect 4364 1158 4924 1188
rect 4364 1148 4854 1158
rect 4814 1108 4854 1148
rect 4254 1068 4764 1108
rect 4814 1068 4924 1108
rect 1774 1028 4214 1038
rect 4814 1028 4854 1068
rect 1064 1018 4854 1028
rect 1064 978 4924 1018
rect 1134 968 4924 978
rect 1134 928 1174 968
rect 1774 958 4214 968
rect 1064 888 1174 928
rect 1214 888 1734 928
rect 1134 848 1174 888
rect 1134 838 1624 848
rect 1064 808 1624 838
rect 1064 798 1174 808
rect 1114 748 1174 798
rect 1664 768 1734 888
rect 1064 688 1174 748
rect 1214 728 1734 768
rect 1064 648 1624 688
rect 1664 608 1734 728
rect 1774 648 1814 958
rect 1854 608 1894 908
rect 1934 648 1974 958
rect 2014 608 2054 908
rect 2094 648 2134 958
rect 2174 608 2214 908
rect 2254 648 2294 958
rect 2334 608 2374 908
rect 2414 648 2454 958
rect 2494 608 2534 908
rect 2574 648 2614 958
rect 2654 608 2694 908
rect 2734 648 2774 958
rect 2814 608 2854 908
rect 2894 658 2934 958
rect 2974 608 3014 908
rect 3054 658 3094 958
rect 3134 608 3174 908
rect 3214 648 3254 958
rect 3294 608 3334 908
rect 3374 648 3414 958
rect 3454 608 3494 908
rect 3534 648 3574 958
rect 3614 608 3654 908
rect 3694 648 3734 958
rect 3774 608 3814 908
rect 3854 648 3894 958
rect 3934 608 3974 908
rect 4014 648 4054 958
rect 4094 608 4134 908
rect 4174 648 4214 958
rect 4254 888 4764 928
rect 4814 918 4854 968
rect 4254 768 4324 888
rect 4814 878 4924 918
rect 4814 848 4854 878
rect 4364 828 4854 848
rect 4364 808 4924 828
rect 4814 788 4924 808
rect 4254 728 4774 768
rect 4814 738 4874 788
rect 4254 608 4324 728
rect 4814 688 4924 738
rect 4364 648 4924 688
rect 1144 588 4844 608
rect 1144 488 1164 588
rect 1284 488 1324 588
rect 1444 488 1484 588
rect 1604 488 1644 588
rect 1764 488 1804 588
rect 1924 488 1964 588
rect 2084 488 2124 588
rect 2244 488 3744 588
rect 3864 488 3904 588
rect 4024 488 4064 588
rect 4184 488 4224 588
rect 4344 488 4384 588
rect 4504 488 4544 588
rect 4664 488 4704 588
rect 4824 488 4844 588
rect 1474 368 1934 378
rect 4054 368 4514 378
rect 5004 368 5084 1628
rect 904 358 5084 368
rect 904 308 1504 358
rect 1904 308 4084 358
rect 4484 308 5084 358
rect 904 288 5084 308
rect 5268 1608 5466 1834
rect 5268 1534 5326 1608
rect 5400 1534 5466 1608
rect 5268 1134 5466 1534
rect 5268 1060 5326 1134
rect 5400 1060 5466 1134
rect 5268 660 5466 1060
rect 5268 586 5326 660
rect 5400 586 5466 660
rect 588 198 786 238
rect 1474 198 1934 288
rect 4054 198 4514 288
rect 5268 198 5466 586
rect 588 130 5466 198
rect 588 56 1182 130
rect 1256 56 1730 130
rect 1804 56 2278 130
rect 2352 56 2826 130
rect 2900 56 3374 130
rect 3448 56 3922 130
rect 3996 56 4472 130
rect 4546 56 5466 130
rect 588 0 5466 56
<< viali >>
rect 624 5324 646 5348
rect 646 5324 720 5348
rect 720 5324 754 5348
rect 624 4948 754 5324
rect 608 4450 744 4808
rect 608 4376 646 4450
rect 646 4376 720 4450
rect 720 4376 744 4450
rect 608 4368 744 4376
rect 608 3976 764 4248
rect 608 3902 646 3976
rect 646 3902 720 3976
rect 720 3902 764 3976
rect 608 3818 764 3902
rect 1164 4998 1284 5098
rect 1324 4998 1444 5098
rect 1484 4998 1604 5098
rect 1644 4998 1764 5098
rect 4224 4998 4344 5098
rect 4384 4998 4504 5098
rect 4544 4998 4664 5098
rect 4704 4998 4824 5098
rect 1084 4708 1114 4758
rect 1114 4708 1134 4758
rect 1084 4618 1114 4668
rect 1114 4618 1134 4668
rect 4854 4698 4874 4748
rect 4874 4698 4904 4748
rect 4854 4608 4874 4658
rect 4874 4608 4904 4658
rect 1084 4518 1114 4568
rect 1114 4518 1134 4568
rect 1084 4428 1114 4478
rect 1114 4428 1134 4478
rect 4854 4508 4874 4558
rect 4874 4508 4904 4558
rect 4854 4418 4874 4468
rect 4874 4418 4904 4468
rect 1164 4078 1284 4178
rect 1324 4078 1444 4178
rect 1484 4078 1604 4178
rect 1644 4078 1764 4178
rect 4224 4078 4344 4178
rect 4384 4078 4504 4178
rect 4544 4078 4664 4178
rect 4704 4078 4824 4178
rect 3772 3572 3808 3608
rect 3848 3572 3884 3608
rect 3924 3572 3960 3608
rect 4000 3572 4036 3608
rect 4076 3572 4112 3608
rect 4152 3572 4188 3608
rect 1152 3444 1186 3480
rect 1230 3444 1264 3480
rect 1302 3444 1336 3480
rect 1386 3444 1420 3478
rect 1470 3444 1504 3478
rect 1554 3444 1588 3478
rect 1638 3444 1672 3478
rect 1722 3444 1756 3478
rect 1806 3444 1840 3478
rect 1890 3444 1924 3478
rect 1974 3444 2008 3478
rect 2058 3444 2092 3478
rect 2148 3444 2182 3478
rect 2694 3454 2728 3488
rect 2778 3454 2812 3488
rect 2862 3454 2896 3488
rect 2946 3454 2980 3488
rect 3030 3454 3064 3488
rect 3114 3454 3148 3488
rect 3198 3454 3232 3488
rect 3282 3454 3316 3488
rect 2284 3278 2434 3428
rect 932 2778 968 2812
rect 1166 2778 1202 2812
rect 920 2644 980 2678
rect 1154 2644 1214 2678
rect 920 2462 980 2496
rect 1154 2462 1214 2496
rect 836 2374 870 2408
rect 1070 2374 1104 2408
rect 1550 3004 1590 3044
rect 1648 2978 1684 3014
rect 1942 3054 1982 3094
rect 2390 3048 2426 3084
rect 2390 2974 2426 3010
rect 2390 2900 2426 2936
rect 2390 2790 2426 2826
rect 3684 3140 3720 3174
rect 3684 3068 3720 3102
rect 4066 3106 4102 3142
rect 2390 2714 2426 2750
rect 2390 2640 2426 2676
rect 604 2122 638 2156
rect 676 2122 710 2156
rect 748 2122 782 2156
rect 932 2112 968 2146
rect 1166 2112 1202 2146
rect 604 2050 638 2084
rect 676 2050 710 2084
rect 748 2050 782 2084
rect 2384 2198 2534 2348
rect 2652 2090 2686 2124
rect 2730 2090 2764 2124
rect 3392 2658 3428 2694
rect 3466 2658 3502 2694
rect 4070 2516 4106 2552
rect 2840 2054 2876 2090
rect 2932 2054 2968 2090
rect 3024 2054 3060 2090
rect 3116 2054 3152 2090
rect 3208 2054 3244 2090
rect 4808 3496 4842 3498
rect 4808 3464 4842 3496
rect 4428 3172 4462 3206
rect 4688 3116 4722 3150
rect 4296 3012 4330 3072
rect 4488 3012 4522 3072
rect 4924 3172 4958 3206
rect 5112 3104 5148 3140
rect 5186 3104 5222 3140
rect 4792 3012 4826 3072
rect 4984 3012 5018 3072
rect 4266 2528 4302 2564
rect 4348 2804 4384 2840
rect 4348 2468 4384 2504
rect 4456 2592 4490 2652
rect 4648 2592 4682 2652
rect 4588 2458 4622 2492
rect 4950 2514 4986 2550
rect 5026 2514 5062 2550
rect 5282 2122 5316 2156
rect 5354 2122 5388 2156
rect 5426 2122 5460 2156
rect 604 1978 638 2012
rect 676 1978 710 2012
rect 748 1978 782 2012
rect 1374 2010 1410 2046
rect 1492 2010 1528 2046
rect 1610 2010 1646 2046
rect 1728 2010 1764 2046
rect 1846 2010 1882 2046
rect 1964 2010 2000 2046
rect 2082 2010 2118 2046
rect 604 1906 638 1940
rect 676 1906 710 1940
rect 748 1906 782 1940
rect 602 1834 636 1868
rect 674 1834 708 1868
rect 746 1834 780 1868
rect 606 1638 764 1768
rect 606 1564 652 1638
rect 652 1564 726 1638
rect 726 1564 764 1638
rect 606 1338 764 1564
rect 3550 1996 3586 2032
rect 3624 1998 3660 2034
rect 3704 1998 3740 2034
rect 3784 1998 3820 2034
rect 3864 1998 3900 2034
rect 5282 2050 5316 2084
rect 5354 2050 5388 2084
rect 5426 2050 5460 2084
rect 5282 1978 5316 2012
rect 5354 1978 5388 2012
rect 5426 1978 5460 2012
rect 5282 1906 5316 1940
rect 5354 1906 5388 1940
rect 5426 1906 5460 1940
rect 5282 1834 5316 1868
rect 5354 1834 5388 1868
rect 5426 1834 5460 1868
rect 614 1164 744 1218
rect 614 1090 652 1164
rect 652 1090 726 1164
rect 726 1090 744 1164
rect 614 778 744 1090
rect 614 616 652 648
rect 652 616 726 648
rect 726 616 774 648
rect 614 238 774 616
rect 1164 1408 1284 1508
rect 1324 1408 1444 1508
rect 1484 1408 1604 1508
rect 1644 1408 1764 1508
rect 4224 1408 4344 1508
rect 4384 1408 4504 1508
rect 4544 1408 4664 1508
rect 4704 1408 4824 1508
rect 1084 1118 1114 1168
rect 1114 1118 1134 1168
rect 1084 1028 1114 1078
rect 1114 1028 1134 1078
rect 4854 1108 4874 1158
rect 4874 1108 4904 1158
rect 4854 1018 4874 1068
rect 4874 1018 4904 1068
rect 1084 928 1114 978
rect 1114 928 1134 978
rect 1084 838 1114 888
rect 1114 838 1134 888
rect 4854 918 4874 968
rect 4874 918 4904 968
rect 4854 828 4874 878
rect 4874 828 4904 878
rect 1164 488 1284 588
rect 1324 488 1444 588
rect 1484 488 1604 588
rect 1644 488 1764 588
rect 4224 488 4344 588
rect 4384 488 4504 588
rect 4544 488 4664 588
rect 4704 488 4824 588
<< metal1 >>
rect 588 5358 1464 5378
rect 588 5348 844 5358
rect 588 4948 624 5348
rect 754 5158 844 5348
rect 1044 5158 1244 5358
rect 1444 5158 1464 5358
rect 754 5138 1464 5158
rect 1944 5358 4044 5378
rect 1944 5158 1964 5358
rect 2164 5158 2184 5358
rect 2384 5158 2904 5358
rect 3084 5158 3604 5358
rect 3804 5158 3824 5358
rect 4024 5158 4044 5358
rect 1944 5138 4044 5158
rect 4524 5358 5164 5378
rect 4524 5158 4544 5358
rect 4744 5158 4944 5358
rect 5144 5158 5164 5358
rect 4524 5138 5164 5158
rect 754 5108 1284 5138
rect 754 5098 2904 5108
rect 754 5038 1164 5098
rect 754 4948 844 5038
rect 588 4908 844 4948
rect 824 4838 844 4908
rect 1044 4998 1164 5038
rect 1284 4998 1324 5098
rect 1444 4998 1484 5098
rect 1604 4998 1644 5098
rect 1764 5078 2904 5098
rect 1764 4998 1784 5078
rect 2934 5048 3054 5138
rect 4704 5108 5164 5138
rect 3084 5098 5164 5108
rect 3084 5078 4224 5098
rect 1814 5018 4174 5048
rect 1044 4988 1784 4998
rect 1044 4838 1064 4988
rect 1154 4978 2904 4988
rect 588 4808 764 4828
rect 824 4808 1064 4838
rect 588 4368 608 4808
rect 744 4368 764 4808
rect 824 4758 1154 4778
rect 824 4748 1084 4758
rect 824 4638 844 4748
rect 1044 4708 1084 4748
rect 1134 4708 1154 4758
rect 1184 4708 1214 4978
rect 1044 4668 1154 4708
rect 1044 4638 1084 4668
rect 824 4618 1084 4638
rect 1134 4648 1154 4668
rect 1244 4648 1274 4948
rect 1304 4708 1334 4978
rect 1364 4648 1394 4948
rect 1424 4708 1454 4978
rect 1484 4648 1514 4948
rect 1544 4708 1574 4978
rect 1664 4958 2904 4978
rect 1604 4648 1634 4948
rect 1664 4868 1784 4958
rect 2934 4928 3054 5018
rect 4204 4998 4224 5078
rect 4344 4998 4384 5098
rect 4504 4998 4544 5098
rect 4664 4998 4704 5098
rect 4824 5038 5164 5098
rect 4824 4998 4944 5038
rect 4204 4988 4944 4998
rect 3084 4978 4834 4988
rect 3084 4958 4324 4978
rect 1814 4898 4174 4928
rect 1664 4838 2904 4868
rect 1664 4748 1784 4838
rect 2934 4808 3054 4898
rect 4204 4868 4324 4958
rect 3084 4838 4324 4868
rect 1814 4778 4174 4808
rect 1664 4718 2904 4748
rect 1664 4678 1784 4718
rect 2934 4688 3054 4778
rect 4204 4748 4324 4838
rect 3084 4718 4324 4748
rect 1814 4658 4174 4688
rect 4204 4678 4324 4718
rect 1134 4628 1634 4648
rect 2934 4628 3054 4658
rect 4354 4648 4384 4948
rect 4414 4708 4444 4978
rect 4474 4648 4504 4948
rect 4534 4708 4564 4978
rect 4594 4648 4624 4948
rect 4654 4708 4684 4978
rect 4714 4648 4744 4948
rect 4774 4708 4804 4978
rect 4924 4838 4944 4988
rect 5144 4838 5164 5038
rect 4924 4808 5164 4838
rect 4834 4748 5164 4768
rect 4834 4698 4854 4748
rect 4904 4698 4944 4748
rect 4834 4658 4944 4698
rect 4834 4648 4854 4658
rect 4354 4628 4854 4648
rect 1134 4618 4854 4628
rect 824 4608 4854 4618
rect 4904 4638 4944 4658
rect 5144 4638 5164 4748
rect 4904 4608 5164 4638
rect 824 4568 5164 4608
rect 824 4538 1084 4568
rect 824 4428 844 4538
rect 1044 4518 1084 4538
rect 1134 4558 5164 4568
rect 1134 4518 4854 4558
rect 1044 4508 4854 4518
rect 4904 4538 5164 4558
rect 4904 4508 4944 4538
rect 1044 4488 4944 4508
rect 1044 4478 1154 4488
rect 1044 4428 1084 4478
rect 1134 4428 1154 4478
rect 824 4408 1154 4428
rect 588 4348 764 4368
rect 824 4338 1064 4368
rect 824 4268 844 4338
rect 588 4248 844 4268
rect 588 3818 608 4248
rect 764 4138 844 4248
rect 1044 4188 1064 4338
rect 1184 4198 1214 4458
rect 1244 4228 1274 4488
rect 1304 4198 1334 4458
rect 1364 4228 1394 4488
rect 1424 4198 1454 4458
rect 1484 4228 1514 4488
rect 1544 4198 1574 4458
rect 1604 4228 1634 4488
rect 1664 4428 2904 4458
rect 1664 4338 1784 4428
rect 2934 4398 3054 4488
rect 3084 4428 4324 4458
rect 1814 4368 4174 4398
rect 1664 4308 2904 4338
rect 1664 4218 1784 4308
rect 2934 4278 3054 4368
rect 4204 4338 4324 4428
rect 3084 4308 4324 4338
rect 1814 4248 4174 4278
rect 1664 4198 2904 4218
rect 1154 4188 2904 4198
rect 1044 4178 1784 4188
rect 1044 4138 1164 4178
rect 764 4078 1164 4138
rect 1284 4078 1324 4178
rect 1444 4078 1484 4178
rect 1604 4078 1644 4178
rect 1764 4098 1784 4178
rect 2934 4158 3054 4248
rect 4204 4218 4324 4308
rect 4354 4228 4384 4488
rect 3084 4198 4324 4218
rect 4414 4198 4444 4458
rect 4474 4228 4504 4488
rect 4534 4198 4564 4458
rect 4594 4228 4624 4488
rect 4654 4198 4684 4458
rect 4714 4228 4744 4488
rect 4834 4468 4944 4488
rect 4774 4198 4804 4458
rect 4834 4418 4854 4468
rect 4904 4428 4944 4468
rect 5144 4428 5164 4538
rect 4904 4418 5164 4428
rect 4834 4398 5164 4418
rect 4924 4338 5164 4368
rect 3084 4188 4834 4198
rect 4924 4188 4944 4338
rect 4204 4178 4944 4188
rect 1814 4128 4174 4158
rect 1764 4078 2904 4098
rect 764 4068 2904 4078
rect 764 4038 1284 4068
rect 2934 4038 3054 4128
rect 4204 4098 4224 4178
rect 3084 4078 4224 4098
rect 4344 4078 4384 4178
rect 4504 4078 4544 4178
rect 4664 4078 4704 4178
rect 4824 4138 4944 4178
rect 5144 4138 5164 4338
rect 4824 4078 5164 4138
rect 3084 4068 5164 4078
rect 4704 4038 5164 4068
rect 764 4018 1464 4038
rect 764 3818 844 4018
rect 1044 3818 1244 4018
rect 1444 3818 1464 4018
rect 588 3798 1464 3818
rect 1944 4018 4044 4038
rect 1944 3818 1964 4018
rect 2164 3818 2184 4018
rect 2384 3818 2904 4018
rect 3084 3818 3604 4018
rect 3804 3818 3824 4018
rect 4024 3818 4044 4018
rect 1944 3798 4044 3818
rect 4524 4018 5164 4038
rect 4524 3818 4544 4018
rect 4744 3818 4944 4018
rect 5144 3818 5164 4018
rect 4524 3798 5164 3818
rect 0 3748 5984 3770
rect 0 3558 64 3748
rect 224 3608 5804 3748
rect 224 3572 3772 3608
rect 3808 3572 3848 3608
rect 3884 3572 3924 3608
rect 3960 3572 4000 3608
rect 4036 3572 4076 3608
rect 4112 3572 4152 3608
rect 4188 3572 5804 3608
rect 224 3558 5804 3572
rect 5964 3558 5984 3748
rect 0 3540 5984 3558
rect 1140 3480 2212 3540
rect 1140 3444 1152 3480
rect 1186 3444 1230 3480
rect 1264 3444 1302 3480
rect 1336 3478 2212 3480
rect 1336 3444 1386 3478
rect 1420 3444 1470 3478
rect 1504 3444 1554 3478
rect 1588 3444 1638 3478
rect 1672 3444 1722 3478
rect 1756 3444 1806 3478
rect 1840 3444 1890 3478
rect 1924 3444 1974 3478
rect 2008 3444 2058 3478
rect 2092 3444 2148 3478
rect 2182 3444 2212 3478
rect 2656 3488 3380 3540
rect 2656 3454 2694 3488
rect 2728 3454 2778 3488
rect 2812 3454 2862 3488
rect 2896 3454 2946 3488
rect 2980 3454 3030 3488
rect 3064 3454 3114 3488
rect 3148 3454 3198 3488
rect 3232 3454 3282 3488
rect 3316 3454 3380 3488
rect 2656 3448 3380 3454
rect 4120 3504 4364 3510
rect 4120 3498 4854 3504
rect 4120 3476 4808 3498
rect 1140 3438 2212 3444
rect 2264 3428 2454 3448
rect 2264 3278 2284 3428
rect 2434 3278 2454 3428
rect 2264 3258 2454 3278
rect 3670 3174 3726 3190
rect 3670 3140 3684 3174
rect 3720 3140 3726 3174
rect 4120 3154 4156 3476
rect 4792 3464 4808 3476
rect 4842 3464 4854 3498
rect 4792 3458 4854 3464
rect 4412 3210 4478 3214
rect 4908 3212 4974 3214
rect 4896 3210 5214 3212
rect 4280 3206 4638 3210
rect 4280 3174 4428 3206
rect 4412 3172 4428 3174
rect 4462 3174 4638 3206
rect 4462 3172 4478 3174
rect 4412 3162 4478 3172
rect 0 3094 1998 3110
rect 3670 3102 3726 3140
rect 0 3082 1942 3094
rect 1926 3054 1942 3082
rect 1982 3054 1998 3094
rect 0 3044 1606 3054
rect 1926 3044 1998 3054
rect 2378 3084 2438 3094
rect 2378 3048 2390 3084
rect 2426 3048 2438 3084
rect 3670 3068 3684 3102
rect 3720 3068 3726 3102
rect 4060 3142 4156 3154
rect 4060 3106 4066 3142
rect 4102 3106 4156 3142
rect 4060 3094 4156 3106
rect 3670 3050 3726 3068
rect 0 3026 1550 3044
rect 1534 3004 1550 3026
rect 1590 3004 1606 3044
rect 1534 2994 1606 3004
rect 1636 3016 1690 3020
rect 2378 3016 2438 3048
rect 1636 3014 2438 3016
rect 1636 3002 1648 3014
rect 1634 2978 1648 3002
rect 1684 3010 2438 3014
rect 1684 2978 2390 3010
rect 1634 2974 2390 2978
rect 2426 2974 2438 3010
rect 1634 2964 2438 2974
rect 2378 2936 2438 2964
rect 2378 2900 2390 2936
rect 2426 2900 2438 2936
rect 2378 2894 2438 2900
rect 4120 2852 4156 3094
rect 4290 3072 4336 3084
rect 4290 3012 4296 3072
rect 4330 3056 4336 3072
rect 4482 3072 4528 3084
rect 4482 3056 4488 3072
rect 4330 3028 4488 3056
rect 4330 3012 4336 3028
rect 4290 3000 4336 3012
rect 4482 3012 4488 3028
rect 4522 3012 4528 3072
rect 4602 3062 4638 3174
rect 4692 3206 5214 3210
rect 4692 3174 4924 3206
rect 4692 3162 4728 3174
rect 4908 3172 4924 3174
rect 4958 3204 5214 3206
rect 4958 3176 6010 3204
rect 4958 3172 4974 3176
rect 4908 3162 4974 3172
rect 4680 3150 4728 3162
rect 4680 3116 4688 3150
rect 4722 3116 4728 3150
rect 4680 3104 4728 3116
rect 5100 3140 5234 3146
rect 5100 3104 5112 3140
rect 5148 3104 5186 3140
rect 5222 3136 5234 3140
rect 5222 3108 6010 3136
rect 5222 3104 5234 3108
rect 5100 3098 5234 3104
rect 4786 3072 4832 3084
rect 4786 3062 4792 3072
rect 4602 3026 4792 3062
rect 4482 3000 4528 3012
rect 4786 3012 4792 3026
rect 4826 3056 4832 3072
rect 4978 3072 5024 3084
rect 4978 3056 4984 3072
rect 4826 3028 4984 3056
rect 4826 3012 4832 3028
rect 4786 3000 4832 3012
rect 4978 3012 4984 3028
rect 5018 3012 5024 3072
rect 4978 3000 5024 3012
rect 4120 2840 4390 2852
rect 2378 2826 2438 2832
rect 900 2812 998 2818
rect 900 2778 932 2812
rect 968 2778 998 2812
rect 900 2772 998 2778
rect 1134 2812 1232 2818
rect 1134 2778 1166 2812
rect 1202 2778 1232 2812
rect 1134 2772 1232 2778
rect 2378 2790 2390 2826
rect 2426 2790 2438 2826
rect 4120 2814 4348 2840
rect 4342 2804 4348 2814
rect 4384 2804 4390 2840
rect 4342 2792 4390 2804
rect 2378 2750 2438 2790
rect 2378 2714 2390 2750
rect 2426 2714 2438 2750
rect 912 2678 990 2692
rect 912 2644 920 2678
rect 980 2644 990 2678
rect 912 2496 990 2644
rect 912 2462 920 2496
rect 980 2462 990 2496
rect 912 2450 990 2462
rect 1146 2678 1224 2692
rect 1146 2644 1154 2678
rect 1214 2644 1224 2678
rect 1146 2496 1224 2644
rect 2378 2678 2438 2714
rect 3382 2694 3512 2710
rect 3382 2678 3392 2694
rect 2378 2676 3392 2678
rect 2378 2640 2390 2676
rect 2426 2658 3392 2676
rect 3428 2658 3466 2694
rect 3502 2658 3512 2694
rect 2426 2642 3512 2658
rect 4450 2652 4496 2664
rect 2426 2640 2438 2642
rect 2378 2634 2438 2640
rect 4450 2592 4456 2652
rect 4490 2636 4496 2652
rect 4642 2652 4688 2664
rect 4642 2636 4648 2652
rect 4490 2608 4648 2636
rect 4490 2592 4496 2608
rect 4450 2580 4496 2592
rect 4642 2592 4648 2608
rect 4682 2592 4688 2652
rect 4642 2580 4688 2592
rect 4260 2564 4308 2576
rect 4064 2554 4124 2564
rect 4260 2554 4266 2564
rect 4064 2552 4266 2554
rect 4064 2516 4070 2552
rect 4106 2528 4266 2552
rect 4302 2528 4308 2564
rect 4106 2516 4308 2528
rect 4938 2550 5074 2556
rect 4064 2504 4124 2516
rect 4342 2504 4390 2516
rect 4938 2514 4950 2550
rect 4986 2514 5026 2550
rect 5062 2546 5074 2550
rect 5062 2518 5328 2546
rect 5062 2514 5074 2518
rect 4938 2508 5074 2514
rect 1146 2462 1154 2496
rect 1214 2462 1224 2496
rect 1146 2450 1224 2462
rect 4342 2468 4348 2504
rect 4384 2490 4390 2504
rect 4572 2492 4638 2502
rect 4572 2490 4588 2492
rect 4384 2468 4588 2490
rect 4342 2458 4588 2468
rect 4622 2458 4638 2492
rect 4342 2454 4638 2458
rect 4342 2452 4440 2454
rect 4572 2450 4638 2454
rect 814 2408 876 2424
rect 814 2406 836 2408
rect 672 2378 836 2406
rect 814 2374 836 2378
rect 870 2374 876 2408
rect 814 2358 876 2374
rect 1054 2408 1110 2424
rect 1054 2374 1070 2408
rect 1104 2390 1110 2408
rect 1104 2374 1314 2390
rect 1054 2358 1314 2374
rect 588 2156 788 2176
rect 588 2122 604 2156
rect 638 2122 676 2156
rect 710 2122 748 2156
rect 782 2146 1242 2156
rect 782 2122 932 2146
rect 588 2112 932 2122
rect 968 2112 1166 2146
rect 1202 2112 1242 2146
rect 588 2084 1242 2112
rect 588 2052 604 2084
rect 0 2050 604 2052
rect 638 2050 676 2084
rect 710 2050 748 2084
rect 782 2052 1242 2084
rect 1272 2134 1314 2358
rect 2364 2348 2554 2368
rect 2364 2198 2384 2348
rect 2534 2198 2554 2348
rect 2364 2178 2554 2198
rect 5268 2156 5466 2176
rect 1272 2124 2780 2134
rect 1272 2090 2652 2124
rect 2686 2090 2730 2124
rect 2764 2090 2780 2124
rect 5268 2122 5282 2156
rect 5316 2122 5354 2156
rect 5388 2122 5426 2156
rect 5460 2122 5466 2156
rect 1272 2080 2780 2090
rect 2816 2090 3268 2096
rect 2816 2054 2840 2090
rect 2876 2054 2932 2090
rect 2968 2054 3024 2090
rect 3060 2054 3116 2090
rect 3152 2054 3208 2090
rect 3244 2054 3268 2090
rect 2816 2052 3268 2054
rect 5268 2084 5466 2122
rect 5268 2052 5282 2084
rect 782 2050 5282 2052
rect 5316 2050 5354 2084
rect 5388 2050 5426 2084
rect 5460 2052 5466 2084
rect 5460 2050 5714 2052
rect 0 2046 5714 2050
rect 0 2028 1374 2046
rect 0 1838 344 2028
rect 504 2024 1374 2028
rect 504 2012 844 2024
rect 504 1978 604 2012
rect 638 1978 676 2012
rect 710 1978 748 2012
rect 782 1978 844 2012
rect 1410 2010 1492 2046
rect 1528 2010 1610 2046
rect 1646 2010 1728 2046
rect 1764 2010 1846 2046
rect 1882 2010 1964 2046
rect 2000 2010 2082 2046
rect 2118 2034 5714 2046
rect 2118 2032 3624 2034
rect 2118 2010 3550 2032
rect 504 1940 844 1978
rect 504 1906 604 1940
rect 638 1906 676 1940
rect 710 1906 748 1940
rect 782 1906 844 1940
rect 504 1868 844 1906
rect 504 1838 602 1868
rect 0 1834 602 1838
rect 636 1834 674 1868
rect 708 1834 746 1868
rect 780 1858 844 1868
rect 1400 1996 3550 2010
rect 3586 1998 3624 2032
rect 3660 1998 3704 2034
rect 3740 1998 3784 2034
rect 3820 1998 3864 2034
rect 3900 2028 5714 2034
rect 3900 2012 5534 2028
rect 3900 1998 5282 2012
rect 3586 1996 5282 1998
rect 1400 1978 5282 1996
rect 5316 1978 5354 2012
rect 5388 1978 5426 2012
rect 5460 1978 5534 2012
rect 1400 1940 5534 1978
rect 1400 1906 5282 1940
rect 5316 1906 5354 1940
rect 5388 1906 5426 1940
rect 5460 1906 5534 1940
rect 1400 1868 5534 1906
rect 1400 1858 5282 1868
rect 780 1834 5282 1858
rect 5316 1834 5354 1868
rect 5388 1834 5426 1868
rect 5460 1838 5534 1868
rect 5694 1838 5714 2028
rect 5460 1834 5714 1838
rect 0 1820 5714 1834
rect 586 1768 1464 1788
rect 586 1338 606 1768
rect 764 1568 844 1768
rect 1044 1568 1244 1768
rect 1444 1568 1464 1768
rect 764 1548 1464 1568
rect 1944 1768 4044 1788
rect 1944 1568 1964 1768
rect 2164 1568 2184 1768
rect 2384 1568 2904 1768
rect 3084 1568 3604 1768
rect 3804 1568 3824 1768
rect 4024 1568 4044 1768
rect 1944 1548 4044 1568
rect 4524 1768 5164 1788
rect 4524 1568 4544 1768
rect 4744 1568 4944 1768
rect 5144 1568 5164 1768
rect 4524 1548 5164 1568
rect 764 1518 1284 1548
rect 764 1508 2904 1518
rect 764 1448 1164 1508
rect 764 1338 844 1448
rect 586 1318 844 1338
rect 824 1248 844 1318
rect 1044 1408 1164 1448
rect 1284 1408 1324 1508
rect 1444 1408 1484 1508
rect 1604 1408 1644 1508
rect 1764 1488 2904 1508
rect 1764 1408 1784 1488
rect 2934 1458 3054 1548
rect 4704 1518 5164 1548
rect 3084 1508 5164 1518
rect 3084 1488 4224 1508
rect 1814 1428 4174 1458
rect 1044 1398 1784 1408
rect 1044 1248 1064 1398
rect 1154 1388 2904 1398
rect 588 1218 764 1238
rect 824 1218 1064 1248
rect 588 778 614 1218
rect 744 778 764 1218
rect 824 1168 1154 1188
rect 824 1158 1084 1168
rect 824 1048 844 1158
rect 1044 1118 1084 1158
rect 1134 1118 1154 1168
rect 1184 1118 1214 1388
rect 1044 1078 1154 1118
rect 1044 1048 1084 1078
rect 824 1028 1084 1048
rect 1134 1058 1154 1078
rect 1244 1058 1274 1358
rect 1304 1118 1334 1388
rect 1364 1058 1394 1358
rect 1424 1118 1454 1388
rect 1484 1058 1514 1358
rect 1544 1118 1574 1388
rect 1664 1368 2904 1388
rect 1604 1058 1634 1358
rect 1664 1278 1784 1368
rect 2934 1338 3054 1428
rect 4204 1408 4224 1488
rect 4344 1408 4384 1508
rect 4504 1408 4544 1508
rect 4664 1408 4704 1508
rect 4824 1448 5164 1508
rect 4824 1408 4944 1448
rect 4204 1398 4944 1408
rect 3084 1388 4834 1398
rect 3084 1368 4324 1388
rect 1814 1308 4174 1338
rect 1664 1248 2904 1278
rect 1664 1158 1784 1248
rect 2934 1218 3054 1308
rect 4204 1278 4324 1368
rect 3084 1248 4324 1278
rect 1814 1188 4174 1218
rect 1664 1128 2904 1158
rect 1664 1088 1784 1128
rect 2934 1098 3054 1188
rect 4204 1158 4324 1248
rect 3084 1128 4324 1158
rect 1814 1068 4174 1098
rect 4204 1088 4324 1128
rect 1134 1038 1634 1058
rect 2934 1038 3054 1068
rect 4354 1058 4384 1358
rect 4414 1118 4444 1388
rect 4474 1058 4504 1358
rect 4534 1118 4564 1388
rect 4594 1058 4624 1358
rect 4654 1118 4684 1388
rect 4714 1058 4744 1358
rect 4774 1118 4804 1388
rect 4924 1248 4944 1398
rect 5144 1248 5164 1448
rect 4924 1218 5164 1248
rect 4834 1158 5164 1178
rect 4834 1108 4854 1158
rect 4904 1108 4944 1158
rect 4834 1068 4944 1108
rect 4834 1058 4854 1068
rect 4354 1038 4854 1058
rect 1134 1028 4854 1038
rect 824 1018 4854 1028
rect 4904 1048 4944 1068
rect 5144 1048 5164 1158
rect 4904 1018 5164 1048
rect 824 978 5164 1018
rect 824 948 1084 978
rect 824 838 844 948
rect 1044 928 1084 948
rect 1134 968 5164 978
rect 1134 928 4854 968
rect 1044 918 4854 928
rect 4904 948 5164 968
rect 4904 918 4944 948
rect 1044 898 4944 918
rect 1044 888 1154 898
rect 1044 838 1084 888
rect 1134 838 1154 888
rect 824 818 1154 838
rect 588 758 764 778
rect 824 748 1064 778
rect 824 678 844 748
rect 588 648 844 678
rect 588 238 614 648
rect 774 548 844 648
rect 1044 598 1064 748
rect 1184 608 1214 868
rect 1244 638 1274 898
rect 1304 608 1334 868
rect 1364 638 1394 898
rect 1424 608 1454 868
rect 1484 638 1514 898
rect 1544 608 1574 868
rect 1604 638 1634 898
rect 1664 838 2904 868
rect 1664 748 1784 838
rect 2934 808 3054 898
rect 3084 838 4324 868
rect 1814 778 4174 808
rect 1664 718 2904 748
rect 1664 628 1784 718
rect 2934 688 3054 778
rect 4204 748 4324 838
rect 3084 718 4324 748
rect 1814 658 4174 688
rect 1664 608 2904 628
rect 1154 598 2904 608
rect 1044 588 1784 598
rect 1044 548 1164 588
rect 774 488 1164 548
rect 1284 488 1324 588
rect 1444 488 1484 588
rect 1604 488 1644 588
rect 1764 508 1784 588
rect 2934 568 3054 658
rect 4204 628 4324 718
rect 4354 638 4384 898
rect 3084 608 4324 628
rect 4414 608 4444 868
rect 4474 638 4504 898
rect 4534 608 4564 868
rect 4594 638 4624 898
rect 4654 608 4684 868
rect 4714 638 4744 898
rect 4834 878 4944 898
rect 4774 608 4804 868
rect 4834 828 4854 878
rect 4904 838 4944 878
rect 5144 838 5164 948
rect 4904 828 5164 838
rect 4834 808 5164 828
rect 4924 748 5164 778
rect 3084 598 4834 608
rect 4924 598 4944 748
rect 4204 588 4944 598
rect 1814 538 4174 568
rect 1764 488 2904 508
rect 774 478 2904 488
rect 774 448 1284 478
rect 2934 448 3054 538
rect 4204 508 4224 588
rect 3084 488 4224 508
rect 4344 488 4384 588
rect 4504 488 4544 588
rect 4664 488 4704 588
rect 4824 548 4944 588
rect 5144 548 5164 748
rect 4824 488 5164 548
rect 3084 478 5164 488
rect 4704 448 5164 478
rect 774 428 1464 448
rect 774 238 844 428
rect 588 228 844 238
rect 1044 228 1244 428
rect 1444 228 1464 428
rect 588 208 1464 228
rect 1944 428 4044 448
rect 1944 228 1964 428
rect 2164 228 2184 428
rect 2384 228 2904 428
rect 3084 228 3604 428
rect 3804 228 3824 428
rect 4024 228 4044 428
rect 1944 208 4044 228
rect 4524 428 5164 448
rect 4524 228 4544 428
rect 4744 228 4944 428
rect 5144 228 5164 428
rect 4524 208 5164 228
<< via1 >>
rect 624 4948 754 5348
rect 844 5158 1044 5358
rect 1244 5158 1444 5358
rect 1964 5158 2164 5358
rect 2184 5158 2384 5358
rect 2904 5158 3084 5358
rect 3604 5158 3804 5358
rect 3824 5158 4024 5358
rect 4544 5158 4744 5358
rect 4944 5158 5144 5358
rect 844 4838 1044 5038
rect 608 4368 744 4808
rect 844 4638 1044 4748
rect 4944 4838 5144 5038
rect 4944 4638 5144 4748
rect 844 4428 1044 4538
rect 844 4138 1044 4338
rect 4944 4428 5144 4538
rect 4944 4138 5144 4338
rect 844 3818 1044 4018
rect 1244 3818 1444 4018
rect 1964 3818 2164 4018
rect 2184 3818 2384 4018
rect 2904 3818 3084 4018
rect 3604 3818 3804 4018
rect 3824 3818 4024 4018
rect 4544 3818 4744 4018
rect 4944 3818 5144 4018
rect 64 3558 224 3748
rect 5804 3558 5964 3748
rect 2284 3278 2434 3428
rect 2384 2198 2534 2348
rect 344 1838 504 2028
rect 844 2010 1374 2024
rect 1374 2010 1400 2024
rect 844 1858 1400 2010
rect 5534 1838 5694 2028
rect 844 1568 1044 1768
rect 1244 1568 1444 1768
rect 1964 1568 2164 1768
rect 2184 1568 2384 1768
rect 2904 1568 3084 1768
rect 3604 1568 3804 1768
rect 3824 1568 4024 1768
rect 4544 1568 4744 1768
rect 4944 1568 5144 1768
rect 844 1248 1044 1448
rect 614 778 744 1218
rect 844 1048 1044 1158
rect 4944 1248 5144 1448
rect 4944 1048 5144 1158
rect 844 838 1044 948
rect 614 238 774 648
rect 844 548 1044 748
rect 4944 838 5144 948
rect 4944 548 5144 748
rect 844 228 1044 428
rect 1244 228 1444 428
rect 1964 228 2164 428
rect 2184 228 2384 428
rect 2904 228 3084 428
rect 3604 228 3804 428
rect 3824 228 4024 428
rect 4544 228 4744 428
rect 4944 228 5144 428
<< metal2 >>
rect 588 5358 1464 5378
rect 588 5348 844 5358
rect 588 4948 624 5348
rect 754 5158 844 5348
rect 1044 5158 1244 5358
rect 1444 5158 1464 5358
rect 754 5138 1464 5158
rect 1944 5358 4044 5378
rect 1944 5158 1964 5358
rect 2164 5158 2184 5358
rect 2384 5158 2904 5358
rect 3084 5158 3604 5358
rect 3804 5158 3824 5358
rect 4024 5158 4044 5358
rect 754 5038 1214 5138
rect 1944 5098 4044 5158
rect 4524 5358 5164 5378
rect 4524 5158 4544 5358
rect 4744 5158 4944 5358
rect 5144 5158 5164 5358
rect 4524 5138 5164 5158
rect 754 4948 844 5038
rect 588 4908 844 4948
rect 824 4838 844 4908
rect 1044 4948 1214 5038
rect 1244 4978 4744 5098
rect 4774 5038 5164 5138
rect 1044 4918 1614 4948
rect 1044 4838 1214 4918
rect 1644 4888 1704 4978
rect 1244 4858 1704 4888
rect 824 4828 1214 4838
rect 588 4808 764 4828
rect 824 4808 1614 4828
rect 588 4368 608 4808
rect 744 4368 764 4808
rect 1104 4798 1614 4808
rect 824 4748 1064 4768
rect 824 4638 844 4748
rect 1044 4638 1064 4748
rect 824 4538 1064 4638
rect 824 4428 844 4538
rect 1044 4428 1064 4538
rect 824 4408 1064 4428
rect 1104 4678 1214 4798
rect 1644 4768 1704 4858
rect 1244 4738 1704 4768
rect 1104 4618 1614 4678
rect 1644 4648 1704 4738
rect 1734 4618 1764 4948
rect 1794 4648 1824 4978
rect 1854 4618 1884 4948
rect 1914 4648 1944 4978
rect 1974 4618 2004 4948
rect 2034 4648 2064 4978
rect 2094 4618 2124 4948
rect 2154 4648 2184 4978
rect 2214 4618 2244 4948
rect 2274 4648 2304 4978
rect 2334 4618 2364 4948
rect 2394 4648 2424 4978
rect 2454 4618 2484 4948
rect 2514 4648 2544 4978
rect 2574 4618 2604 4948
rect 2634 4648 2664 4978
rect 2694 4618 2724 4948
rect 2754 4648 2784 4978
rect 2814 4618 2844 4948
rect 2874 4648 2904 4978
rect 2934 4618 3054 4948
rect 3084 4648 3114 4978
rect 3144 4618 3174 4948
rect 3204 4648 3234 4978
rect 3264 4618 3294 4948
rect 3324 4648 3354 4978
rect 3384 4618 3414 4948
rect 3444 4648 3474 4978
rect 3504 4618 3534 4948
rect 3564 4648 3594 4978
rect 3624 4618 3654 4948
rect 3684 4648 3714 4978
rect 3744 4618 3774 4948
rect 3804 4648 3834 4978
rect 3864 4618 3894 4948
rect 3924 4648 3954 4978
rect 3984 4618 4014 4948
rect 4044 4648 4074 4978
rect 4104 4618 4134 4948
rect 4164 4648 4194 4978
rect 4224 4618 4254 4948
rect 4284 4888 4344 4978
rect 4774 4948 4944 5038
rect 4374 4918 4944 4948
rect 4284 4858 4744 4888
rect 4284 4768 4344 4858
rect 4774 4838 4944 4918
rect 5144 4838 5164 5038
rect 4774 4828 5164 4838
rect 4374 4808 5164 4828
rect 4374 4798 4884 4808
rect 4284 4738 4744 4768
rect 4284 4648 4344 4738
rect 4774 4678 4884 4798
rect 4374 4618 4884 4678
rect 1104 4558 4884 4618
rect 1104 4468 1614 4558
rect 1104 4378 1214 4468
rect 1644 4438 1704 4528
rect 1244 4408 1704 4438
rect 1104 4368 1614 4378
rect 588 4348 764 4368
rect 824 4348 1614 4368
rect 824 4338 1214 4348
rect 824 4138 844 4338
rect 1044 4258 1214 4338
rect 1644 4318 1704 4408
rect 1244 4288 1704 4318
rect 1044 4228 1614 4258
rect 1044 4138 1214 4228
rect 1644 4198 1704 4288
rect 1734 4228 1764 4558
rect 1794 4198 1824 4528
rect 1854 4228 1884 4558
rect 1914 4198 1944 4528
rect 1974 4228 2004 4558
rect 2034 4198 2064 4528
rect 2094 4228 2124 4558
rect 2154 4198 2184 4528
rect 2214 4228 2244 4558
rect 2274 4198 2304 4528
rect 2334 4228 2364 4558
rect 2394 4198 2424 4528
rect 2454 4228 2484 4558
rect 2514 4198 2544 4528
rect 2574 4228 2604 4558
rect 2634 4198 2664 4528
rect 2694 4228 2724 4558
rect 2754 4198 2784 4528
rect 2814 4228 2844 4558
rect 2874 4198 2904 4528
rect 2934 4228 3054 4558
rect 3084 4198 3114 4528
rect 3144 4228 3174 4558
rect 3204 4198 3234 4528
rect 3264 4228 3294 4558
rect 3324 4198 3354 4528
rect 3384 4228 3414 4558
rect 3444 4198 3474 4528
rect 3504 4228 3534 4558
rect 3564 4198 3594 4528
rect 3624 4228 3654 4558
rect 3684 4198 3714 4528
rect 3744 4228 3774 4558
rect 3804 4198 3834 4528
rect 3864 4228 3894 4558
rect 3924 4198 3954 4528
rect 3984 4228 4014 4558
rect 4044 4198 4074 4528
rect 4104 4228 4134 4558
rect 4164 4198 4194 4528
rect 4224 4228 4254 4558
rect 4284 4438 4344 4528
rect 4374 4468 4884 4558
rect 4284 4408 4744 4438
rect 4284 4318 4344 4408
rect 4774 4378 4884 4468
rect 4924 4748 5164 4768
rect 4924 4638 4944 4748
rect 5144 4638 5164 4748
rect 4924 4538 5164 4638
rect 4924 4428 4944 4538
rect 5144 4428 5164 4538
rect 4924 4408 5164 4428
rect 4374 4368 4884 4378
rect 4374 4348 5164 4368
rect 4774 4338 5164 4348
rect 4284 4288 4744 4318
rect 4284 4198 4344 4288
rect 4774 4258 4944 4338
rect 4374 4228 4944 4258
rect 824 4038 1214 4138
rect 1244 4078 4744 4198
rect 4774 4138 4944 4228
rect 5144 4138 5164 4338
rect 824 4018 1464 4038
rect 824 3818 844 4018
rect 1044 3818 1244 4018
rect 1444 3818 1464 4018
rect 824 3798 1464 3818
rect 1944 4018 4044 4078
rect 4774 4038 5164 4138
rect 1944 3818 1964 4018
rect 2164 3818 2184 4018
rect 2384 3818 2904 4018
rect 3084 3818 3604 4018
rect 3804 3818 3824 4018
rect 4024 3818 4044 4018
rect 1944 3798 4044 3818
rect 4524 4018 5164 4038
rect 4524 3818 4544 4018
rect 4744 3818 4944 4018
rect 5144 3818 5164 4018
rect 4524 3798 5164 3818
rect 46 3748 246 3770
rect 46 3558 64 3748
rect 224 3558 246 3748
rect 46 3540 246 3558
rect 2264 3428 2454 3798
rect 5784 3748 5984 3770
rect 5784 3558 5804 3748
rect 5964 3558 5984 3748
rect 5784 3540 5984 3558
rect 2264 3278 2284 3428
rect 2434 3278 2454 3428
rect 2264 3258 2454 3278
rect 2364 2348 2554 2368
rect 2364 2198 2384 2348
rect 2534 2198 2554 2348
rect 322 2028 522 2052
rect 322 1838 344 2028
rect 504 1838 522 2028
rect 816 2024 1446 2052
rect 816 1858 844 2024
rect 1400 1858 1446 2024
rect 816 1852 1446 1858
rect 322 1820 522 1838
rect 824 1788 1454 1852
rect 2364 1788 2554 2198
rect 5514 2028 5714 2052
rect 5514 1838 5534 2028
rect 5694 1838 5714 2028
rect 5514 1820 5714 1838
rect 824 1768 1464 1788
rect 824 1568 844 1768
rect 1044 1568 1244 1768
rect 1444 1568 1464 1768
rect 824 1548 1464 1568
rect 1944 1768 4044 1788
rect 1944 1568 1964 1768
rect 2164 1568 2184 1768
rect 2384 1568 2904 1768
rect 3084 1568 3604 1768
rect 3804 1568 3824 1768
rect 4024 1568 4044 1768
rect 824 1448 1214 1548
rect 1944 1508 4044 1568
rect 4524 1768 5164 1788
rect 4524 1568 4544 1768
rect 4744 1568 4944 1768
rect 5144 1568 5164 1768
rect 4524 1548 5164 1568
rect 824 1248 844 1448
rect 1044 1358 1214 1448
rect 1244 1388 4744 1508
rect 4774 1448 5164 1548
rect 1044 1328 1614 1358
rect 1044 1248 1214 1328
rect 1644 1298 1704 1388
rect 1244 1268 1704 1298
rect 824 1238 1214 1248
rect 588 1218 764 1238
rect 824 1218 1614 1238
rect 588 778 614 1218
rect 744 778 764 1218
rect 1104 1208 1614 1218
rect 824 1158 1064 1178
rect 824 1048 844 1158
rect 1044 1048 1064 1158
rect 824 948 1064 1048
rect 824 838 844 948
rect 1044 838 1064 948
rect 824 818 1064 838
rect 1104 1088 1214 1208
rect 1644 1178 1704 1268
rect 1244 1148 1704 1178
rect 1104 1028 1614 1088
rect 1644 1058 1704 1148
rect 1734 1028 1764 1358
rect 1794 1058 1824 1388
rect 1854 1028 1884 1358
rect 1914 1058 1944 1388
rect 1974 1028 2004 1358
rect 2034 1058 2064 1388
rect 2094 1028 2124 1358
rect 2154 1058 2184 1388
rect 2214 1028 2244 1358
rect 2274 1058 2304 1388
rect 2334 1028 2364 1358
rect 2394 1058 2424 1388
rect 2454 1028 2484 1358
rect 2514 1058 2544 1388
rect 2574 1028 2604 1358
rect 2634 1058 2664 1388
rect 2694 1028 2724 1358
rect 2754 1058 2784 1388
rect 2814 1028 2844 1358
rect 2874 1058 2904 1388
rect 2934 1028 3054 1358
rect 3084 1058 3114 1388
rect 3144 1028 3174 1358
rect 3204 1058 3234 1388
rect 3264 1028 3294 1358
rect 3324 1058 3354 1388
rect 3384 1028 3414 1358
rect 3444 1058 3474 1388
rect 3504 1028 3534 1358
rect 3564 1058 3594 1388
rect 3624 1028 3654 1358
rect 3684 1058 3714 1388
rect 3744 1028 3774 1358
rect 3804 1058 3834 1388
rect 3864 1028 3894 1358
rect 3924 1058 3954 1388
rect 3984 1028 4014 1358
rect 4044 1058 4074 1388
rect 4104 1028 4134 1358
rect 4164 1058 4194 1388
rect 4224 1028 4254 1358
rect 4284 1298 4344 1388
rect 4774 1358 4944 1448
rect 4374 1328 4944 1358
rect 4284 1268 4744 1298
rect 4284 1178 4344 1268
rect 4774 1248 4944 1328
rect 5144 1248 5164 1448
rect 4774 1238 5164 1248
rect 4374 1218 5164 1238
rect 4374 1208 4884 1218
rect 4284 1148 4744 1178
rect 4284 1058 4344 1148
rect 4774 1088 4884 1208
rect 4374 1028 4884 1088
rect 1104 968 4884 1028
rect 1104 878 1614 968
rect 1104 788 1214 878
rect 1644 848 1704 938
rect 1244 818 1704 848
rect 1104 778 1614 788
rect 588 758 764 778
rect 824 758 1614 778
rect 824 748 1214 758
rect 824 678 844 748
rect 588 648 844 678
rect 588 238 614 648
rect 774 548 844 648
rect 1044 668 1214 748
rect 1644 728 1704 818
rect 1244 698 1704 728
rect 1044 638 1614 668
rect 1044 548 1214 638
rect 1644 608 1704 698
rect 1734 638 1764 968
rect 1794 608 1824 938
rect 1854 638 1884 968
rect 1914 608 1944 938
rect 1974 638 2004 968
rect 2034 608 2064 938
rect 2094 638 2124 968
rect 2154 608 2184 938
rect 2214 638 2244 968
rect 2274 608 2304 938
rect 2334 638 2364 968
rect 2394 608 2424 938
rect 2454 638 2484 968
rect 2514 608 2544 938
rect 2574 638 2604 968
rect 2634 608 2664 938
rect 2694 638 2724 968
rect 2754 608 2784 938
rect 2814 638 2844 968
rect 2874 608 2904 938
rect 2934 638 3054 968
rect 3084 608 3114 938
rect 3144 638 3174 968
rect 3204 608 3234 938
rect 3264 638 3294 968
rect 3324 608 3354 938
rect 3384 638 3414 968
rect 3444 608 3474 938
rect 3504 638 3534 968
rect 3564 608 3594 938
rect 3624 638 3654 968
rect 3684 608 3714 938
rect 3744 638 3774 968
rect 3804 608 3834 938
rect 3864 638 3894 968
rect 3924 608 3954 938
rect 3984 638 4014 968
rect 4044 608 4074 938
rect 4104 638 4134 968
rect 4164 608 4194 938
rect 4224 638 4254 968
rect 4284 848 4344 938
rect 4374 878 4884 968
rect 4284 818 4744 848
rect 4284 728 4344 818
rect 4774 788 4884 878
rect 4924 1158 5164 1178
rect 4924 1048 4944 1158
rect 5144 1048 5164 1158
rect 4924 948 5164 1048
rect 4924 838 4944 948
rect 5144 838 5164 948
rect 4924 818 5164 838
rect 4374 778 4884 788
rect 4374 758 5164 778
rect 4774 748 5164 758
rect 4284 698 4744 728
rect 4284 608 4344 698
rect 4774 668 4944 748
rect 4374 638 4944 668
rect 774 448 1214 548
rect 1244 488 4744 608
rect 4774 548 4944 638
rect 5144 548 5164 748
rect 774 428 1464 448
rect 774 238 844 428
rect 588 228 844 238
rect 1044 228 1244 428
rect 1444 228 1464 428
rect 588 208 1464 228
rect 1944 428 4044 488
rect 4774 448 5164 548
rect 1944 228 1964 428
rect 2164 228 2184 428
rect 2384 228 2904 428
rect 3084 228 3604 428
rect 3804 228 3824 428
rect 4024 228 4044 428
rect 1944 208 4044 228
rect 4524 428 5164 448
rect 4524 228 4544 428
rect 4744 228 4944 428
rect 5144 228 5164 428
rect 4524 208 5164 228
<< via2 >>
rect 624 4948 754 5348
rect 608 4368 744 4808
rect 64 3558 224 3748
rect 5804 3558 5964 3748
rect 344 1838 504 2028
rect 844 1858 1400 2024
rect 5534 1838 5694 2028
rect 614 778 744 1218
rect 614 238 774 648
<< metal3 >>
rect 588 5358 1464 5378
rect 588 5348 844 5358
rect 588 4948 624 5348
rect 754 5188 844 5348
rect 1014 5188 1264 5358
rect 1434 5188 1464 5358
rect 1944 5358 4044 5378
rect 1944 5228 1964 5358
rect 2094 5228 2124 5358
rect 2254 5228 3734 5358
rect 3864 5228 3894 5358
rect 4024 5228 4044 5358
rect 1944 5208 4044 5228
rect 4524 5358 5164 5378
rect 754 5128 1464 5188
rect 4524 5188 4554 5358
rect 4724 5188 4974 5358
rect 5144 5188 5164 5358
rect 4524 5128 5164 5188
rect 754 5098 5164 5128
rect 754 4948 844 5098
rect 588 4928 844 4948
rect 1014 4928 4974 5098
rect 5144 4928 5164 5098
rect 588 4908 5164 4928
rect 824 4898 5164 4908
rect 588 4808 764 4828
rect 588 4368 608 4808
rect 744 4368 764 4808
rect 588 4348 764 4368
rect 824 4808 994 4828
rect 824 4608 844 4808
rect 974 4608 994 4808
rect 824 4568 994 4608
rect 824 4368 844 4568
rect 974 4368 994 4568
rect 824 4348 994 4368
rect 1074 4278 4914 4898
rect 4994 4808 5164 4828
rect 4994 4608 5014 4808
rect 5144 4608 5164 4808
rect 4994 4568 5164 4608
rect 4994 4368 5014 4568
rect 5144 4368 5164 4568
rect 4994 4348 5164 4368
rect 824 4248 5164 4278
rect 824 4078 844 4248
rect 1014 4078 4974 4248
rect 5144 4078 5164 4248
rect 824 4048 5164 4078
rect 824 3988 1464 4048
rect 824 3818 844 3988
rect 1014 3818 1264 3988
rect 1434 3818 1464 3988
rect 4524 3988 5164 4048
rect 824 3798 1464 3818
rect 1944 3948 4044 3968
rect 1944 3818 1964 3948
rect 2094 3818 2124 3948
rect 2254 3818 3734 3948
rect 3864 3818 3894 3948
rect 4024 3818 4044 3948
rect 1944 3798 4044 3818
rect 4524 3818 4554 3988
rect 4724 3818 4974 3988
rect 5144 3818 5164 3988
rect 4524 3798 5164 3818
rect 46 3748 246 3770
rect 46 3558 64 3748
rect 224 3558 246 3748
rect 46 3540 246 3558
rect 5784 3748 5984 3770
rect 5784 3558 5804 3748
rect 5964 3558 5984 3748
rect 5784 3540 5984 3558
rect 322 2028 522 2052
rect 322 1838 344 2028
rect 504 1838 522 2028
rect 816 2024 1446 2052
rect 816 1858 844 2024
rect 1400 1858 1446 2024
rect 816 1852 1446 1858
rect 5514 2028 5714 2052
rect 322 1820 522 1838
rect 5514 1838 5534 2028
rect 5694 1838 5714 2028
rect 5514 1820 5714 1838
rect 824 1768 1464 1788
rect 824 1598 844 1768
rect 1014 1598 1264 1768
rect 1434 1598 1464 1768
rect 1944 1768 4044 1788
rect 1944 1638 1964 1768
rect 2094 1638 2124 1768
rect 2254 1638 3734 1768
rect 3864 1638 3894 1768
rect 4024 1638 4044 1768
rect 1944 1618 4044 1638
rect 4524 1768 5164 1788
rect 824 1538 1464 1598
rect 4524 1598 4554 1768
rect 4724 1598 4974 1768
rect 5144 1598 5164 1768
rect 4524 1538 5164 1598
rect 824 1508 5164 1538
rect 824 1338 844 1508
rect 1014 1338 4974 1508
rect 5144 1338 5164 1508
rect 824 1308 5164 1338
rect 588 1218 764 1238
rect 588 778 614 1218
rect 744 778 764 1218
rect 588 758 764 778
rect 824 1218 994 1238
rect 824 1018 844 1218
rect 974 1018 994 1218
rect 824 978 994 1018
rect 824 778 844 978
rect 974 778 994 978
rect 824 758 994 778
rect 1074 688 4914 1308
rect 4994 1218 5164 1238
rect 4994 1018 5014 1218
rect 5144 1018 5164 1218
rect 4994 978 5164 1018
rect 4994 778 5014 978
rect 5144 778 5164 978
rect 4994 758 5164 778
rect 824 678 5164 688
rect 588 658 5164 678
rect 588 648 844 658
rect 588 238 614 648
rect 774 488 844 648
rect 1014 488 4974 658
rect 5144 488 5164 658
rect 774 458 5164 488
rect 774 398 1464 458
rect 774 238 844 398
rect 588 228 844 238
rect 1014 228 1264 398
rect 1434 228 1464 398
rect 4524 398 5164 458
rect 588 208 1464 228
rect 1944 358 4044 378
rect 1944 228 1964 358
rect 2094 228 2124 358
rect 2254 228 3734 358
rect 3864 228 3894 358
rect 4024 228 4044 358
rect 1944 208 4044 228
rect 4524 228 4554 398
rect 4724 228 4974 398
rect 5144 228 5164 398
rect 4524 208 5164 228
<< via3 >>
rect 624 4948 754 5348
rect 844 5188 1014 5358
rect 1264 5188 1434 5358
rect 1964 5228 2094 5358
rect 2124 5228 2254 5358
rect 3734 5228 3864 5358
rect 3894 5228 4024 5358
rect 4554 5188 4724 5358
rect 4974 5188 5144 5358
rect 844 4928 1014 5098
rect 4974 4928 5144 5098
rect 608 4368 744 4808
rect 844 4608 974 4808
rect 844 4368 974 4568
rect 5014 4608 5144 4808
rect 5014 4368 5144 4568
rect 844 4078 1014 4248
rect 4974 4078 5144 4248
rect 844 3818 1014 3988
rect 1264 3818 1434 3988
rect 1964 3818 2094 3948
rect 2124 3818 2254 3948
rect 3734 3818 3864 3948
rect 3894 3818 4024 3948
rect 4554 3818 4724 3988
rect 4974 3818 5144 3988
rect 64 3558 224 3748
rect 5804 3558 5964 3748
rect 344 1838 504 2028
rect 5534 1838 5694 2028
rect 844 1598 1014 1768
rect 1264 1598 1434 1768
rect 1964 1638 2094 1768
rect 2124 1638 2254 1768
rect 3734 1638 3864 1768
rect 3894 1638 4024 1768
rect 4554 1598 4724 1768
rect 4974 1598 5144 1768
rect 844 1338 1014 1508
rect 4974 1338 5144 1508
rect 614 778 744 1218
rect 844 1018 974 1218
rect 844 778 974 978
rect 5014 1018 5144 1218
rect 5014 778 5144 978
rect 614 238 774 648
rect 844 488 1014 658
rect 4974 488 5144 658
rect 844 228 1014 398
rect 1264 228 1434 398
rect 1964 228 2094 358
rect 2124 228 2254 358
rect 3734 228 3864 358
rect 3894 228 4024 358
rect 4554 228 4724 398
rect 4974 228 5144 398
<< mimcap >>
rect 1104 5068 4884 5098
rect 1104 4108 1134 5068
rect 4854 4108 4884 5068
rect 1104 4078 4884 4108
rect 1104 1478 4884 1508
rect 1104 518 1134 1478
rect 4854 518 4884 1478
rect 1104 488 4884 518
<< mimcapcontact >>
rect 1134 4108 4854 5068
rect 1134 518 4854 1478
<< metal4 >>
rect 46 3748 246 5596
rect 46 3558 64 3748
rect 224 3558 246 3748
rect 46 0 246 3558
rect 322 2028 522 5596
rect 588 5358 1454 5378
rect 588 5348 844 5358
rect 588 4948 624 5348
rect 754 5188 844 5348
rect 1014 5188 1264 5358
rect 1434 5188 1454 5358
rect 754 5168 1454 5188
rect 1944 5358 4044 5378
rect 1944 5228 1964 5358
rect 2094 5228 2124 5358
rect 2254 5228 3734 5358
rect 3864 5228 3894 5358
rect 4024 5228 4044 5358
rect 754 5098 1034 5168
rect 754 4948 844 5098
rect 588 4928 844 4948
rect 1014 4928 1034 5098
rect 1944 5088 4044 5228
rect 4534 5358 5164 5378
rect 4534 5188 4554 5358
rect 4724 5188 4974 5358
rect 5144 5188 5164 5358
rect 4534 5168 5164 5188
rect 4954 5098 5164 5168
rect 588 4908 1034 4928
rect 1114 5068 4874 5088
rect 1114 4828 1134 5068
rect 588 4808 1134 4828
rect 588 4368 608 4808
rect 744 4608 844 4808
rect 974 4608 1134 4808
rect 744 4568 1134 4608
rect 744 4368 844 4568
rect 974 4368 1134 4568
rect 588 4348 1134 4368
rect 824 4248 1034 4268
rect 824 4078 844 4248
rect 1014 4078 1034 4248
rect 1114 4108 1134 4348
rect 4854 4828 4874 5068
rect 4954 4928 4974 5098
rect 5144 4928 5164 5098
rect 4954 4908 5164 4928
rect 4854 4808 5164 4828
rect 4854 4608 5014 4808
rect 5144 4608 5164 4808
rect 4854 4568 5164 4608
rect 4854 4368 5014 4568
rect 5144 4368 5164 4568
rect 4854 4348 5164 4368
rect 4854 4108 4874 4348
rect 1114 4088 4874 4108
rect 4954 4248 5164 4268
rect 824 4008 1034 4078
rect 824 3988 1454 4008
rect 824 3818 844 3988
rect 1014 3818 1264 3988
rect 1434 3818 1454 3988
rect 824 3798 1454 3818
rect 1944 3948 4044 4088
rect 4954 4078 4974 4248
rect 5144 4078 5164 4248
rect 4954 4008 5164 4078
rect 1944 3818 1964 3948
rect 2094 3818 2124 3948
rect 2254 3818 3734 3948
rect 3864 3818 3894 3948
rect 4024 3818 4044 3948
rect 1944 3798 4044 3818
rect 4534 3988 5164 4008
rect 4534 3818 4554 3988
rect 4724 3818 4974 3988
rect 5144 3818 5164 3988
rect 4534 3798 5164 3818
rect 322 1838 344 2028
rect 504 1838 522 2028
rect 322 0 522 1838
rect 5514 2028 5714 5596
rect 5514 1838 5534 2028
rect 5694 1838 5714 2028
rect 824 1768 1454 1788
rect 824 1598 844 1768
rect 1014 1598 1264 1768
rect 1434 1598 1454 1768
rect 824 1578 1454 1598
rect 1944 1768 4044 1788
rect 1944 1638 1964 1768
rect 2094 1638 2124 1768
rect 2254 1638 3734 1768
rect 3864 1638 3894 1768
rect 4024 1638 4044 1768
rect 824 1508 1034 1578
rect 824 1338 844 1508
rect 1014 1338 1034 1508
rect 1944 1498 4044 1638
rect 4534 1768 5164 1788
rect 4534 1598 4554 1768
rect 4724 1598 4974 1768
rect 5144 1598 5164 1768
rect 4534 1578 5164 1598
rect 4954 1508 5164 1578
rect 824 1318 1034 1338
rect 1114 1478 4874 1498
rect 1114 1238 1134 1478
rect 588 1218 1134 1238
rect 588 778 614 1218
rect 744 1018 844 1218
rect 974 1018 1134 1218
rect 744 978 1134 1018
rect 744 778 844 978
rect 974 778 1134 978
rect 588 758 1134 778
rect 588 658 1034 678
rect 588 648 844 658
rect 588 238 614 648
rect 774 488 844 648
rect 1014 488 1034 658
rect 1114 518 1134 758
rect 4854 1238 4874 1478
rect 4954 1338 4974 1508
rect 5144 1338 5164 1508
rect 4954 1318 5164 1338
rect 4854 1218 5164 1238
rect 4854 1018 5014 1218
rect 5144 1018 5164 1218
rect 4854 978 5164 1018
rect 4854 778 5014 978
rect 5144 778 5164 978
rect 4854 758 5164 778
rect 4854 518 4874 758
rect 1114 498 4874 518
rect 4954 658 5164 678
rect 774 418 1034 488
rect 774 398 1454 418
rect 774 238 844 398
rect 588 228 844 238
rect 1014 228 1264 398
rect 1434 228 1454 398
rect 588 208 1454 228
rect 1944 358 4044 498
rect 4954 488 4974 658
rect 5144 488 5164 658
rect 4954 418 5164 488
rect 1944 228 1964 358
rect 2094 228 2124 358
rect 2254 228 3734 358
rect 3864 228 3894 358
rect 4024 228 4044 358
rect 1944 208 4044 228
rect 4534 398 5164 418
rect 4534 228 4554 398
rect 4724 228 4974 398
rect 5144 228 5164 398
rect 4534 208 5164 228
rect 5514 0 5714 1838
rect 5784 3748 5984 5596
rect 5784 3558 5804 3748
rect 5964 3558 5984 3748
rect 5784 0 5984 3558
<< comment >>
rect 1368 3320 1400 3362
rect 1564 3316 1596 3358
rect 1754 3314 1786 3356
rect 1946 3314 1978 3356
rect 2138 3316 2170 3358
rect 2606 3028 2624 3232
rect 2828 3040 2848 3260
rect 3022 3012 3042 3232
rect 3216 3070 3236 3290
rect 4378 3264 4398 3412
rect 4486 3264 4524 3400
rect 4612 3258 4632 3406
rect 4874 3264 4894 3412
rect 4982 3264 5020 3400
rect 5108 3258 5128 3406
rect 3856 3240 3890 3254
rect 4048 3242 4082 3256
rect 3442 3028 3460 3232
rect 3856 3044 3890 3056
rect 4048 3044 4082 3056
rect 4394 3018 4422 3066
rect 4890 3018 4918 3066
rect 1374 2626 1406 2668
rect 1562 2640 1594 2682
rect 1750 2642 1782 2684
rect 1954 2646 1986 2688
rect 2142 2654 2174 2696
rect 3856 2604 3890 2616
rect 4048 2604 4082 2616
rect 4554 2598 4582 2646
rect 2822 2322 2850 2490
rect 3016 2320 3044 2488
rect 3208 2306 3236 2474
rect 3856 2406 3890 2420
rect 4048 2404 4082 2418
rect 1466 2238 1498 2280
rect 1664 2236 1696 2278
rect 1852 2238 1884 2280
rect 2040 2238 2072 2280
rect 4538 2252 4558 2400
rect 4646 2264 4684 2400
rect 4772 2258 4792 2406
<< labels >>
flabel metal1 s 0 3026 14 3054 7 FreeSans 160 0 0 0 inn
port 30 w analog input
flabel metal1 s 0 3082 14 3110 7 FreeSans 160 0 0 0 inp
port 31 w analog input
flabel metal1 s 0 3540 28 3770 7 FreeSans 160 0 0 0 VDD
port 27 w power bidirectional
flabel metal1 s 0 1820 22 2052 7 FreeSans 160 0 0 0 VSS
port 26 w power bidirectional
flabel metal1 s 5848 3176 6010 3204 3 FreeSans 160 0 0 0 latch_q
port 21 e signal output
flabel metal1 s 5848 3108 6010 3136 3 FreeSans 160 0 0 0 latch_qn
port 22 e signal output
flabel metal1 s 5166 2518 5328 2546 3 FreeSans 160 0 0 0 comp_trig
port 23 e signal output
flabel metal1 s 672 2378 686 2406 7 FreeSans 160 0 0 0 clk
port 32 w signal input
rlabel poly 4248 3108 4248 3140 7 NOR-Latch_0/R
rlabel metal1 4242 3478 4242 3510 7 NOR-Latch_0/S
rlabel locali 4336 3538 4336 3572 7 NOR-Latch_0/VDD
rlabel locali 5210 3108 5210 3148 3 NOR-Latch_0/QN
rlabel metal1 5214 3176 5214 3212 3 NOR-Latch_0/Q
rlabel locali 4366 2912 4366 2946 7 NOR-Latch_0/VSS
rlabel locali 4832 3538 4832 3572 7 NOR-Latch_0/NOR_1/VDD
rlabel locali 5210 3108 5210 3146 3 NOR-Latch_0/NOR_1/Q
rlabel metal1 4776 3174 4776 3210 7 NOR-Latch_0/NOR_1/B
rlabel locali 4792 3452 4792 3504 7 NOR-Latch_0/NOR_1/A
rlabel locali 4864 2912 4864 2946 7 NOR-Latch_0/NOR_1/VSS
rlabel locali 4336 3538 4336 3572 7 NOR-Latch_0/NOR_0/VDD
rlabel locali 4714 3108 4714 3146 3 NOR-Latch_0/NOR_0/Q
rlabel metal1 4280 3174 4280 3210 7 NOR-Latch_0/NOR_0/B
rlabel locali 4296 3452 4296 3504 7 NOR-Latch_0/NOR_0/A
rlabel locali 4368 2912 4368 2946 7 NOR-Latch_0/NOR_0/VSS
rlabel locali 4496 2092 4496 2126 7 NOR_0/VDD
rlabel locali 4874 2518 4874 2556 3 NOR_0/Q
rlabel metal1 4440 2454 4440 2490 7 NOR_0/B
rlabel locali 4456 2160 4456 2212 7 NOR_0/A
rlabel locali 4528 2718 4528 2752 7 NOR_0/VSS
rlabel locali 2484 2776 2484 2810 7 adc_comp_circuit_0/bn
rlabel locali 3574 2776 3574 2810 3 adc_comp_circuit_0/bp
rlabel locali 4136 2516 4136 2554 3 adc_comp_circuit_0/outn
rlabel locali 4134 3106 4134 3144 3 adc_comp_circuit_0/outp
rlabel locali 1848 2928 1848 2960 7 adc_comp_circuit_0/on
rlabel locali 1464 2928 1464 2960 7 adc_comp_circuit_0/op
rlabel locali 2714 2080 2714 2134 7 adc_comp_circuit_0/nclk
rlabel locali 1268 2334 1268 2364 7 adc_comp_circuit_0/clk
flabel metal4 5514 0 5714 5596 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VSS
flabel metal4 5784 0 5984 5596 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VDD
flabel metal4 322 0 522 5596 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VSS
flabel metal4 46 0 246 5596 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VDD
rlabel metal1 0 3082 0 3110 7 adc_comp_circuit_0/inp
rlabel metal1 0 3026 0 3054 7 adc_comp_circuit_0/inn
rlabel metal1 0 1894 0 2052 7 adc_comp_circuit_0/VSS
rlabel metal1 0 3540 0 3678 7 adc_comp_circuit_0/VDD
flabel metal1 824 3798 1464 4038 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 824 5138 1464 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 4524 3798 5164 4038 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 4524 5138 5164 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 824 4808 1064 5378 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 824 3798 1064 4368 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 4924 3798 5164 4368 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 4924 4808 5164 5378 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 1944 3798 4044 4038 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel metal1 1944 5138 4044 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel metal1 824 4408 1064 4778 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel metal1 4924 4398 5164 4768 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel locali 1474 3798 1934 3878 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel locali 4054 3798 4514 3878 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel locali 1474 5298 1934 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel locali 4054 5298 4514 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel metal3 824 3798 1464 4038 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 4524 3798 5164 4038 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 824 5138 1464 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 4524 5138 5164 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 824 4898 1074 5378 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 824 3798 1074 4278 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 4914 3798 5164 4278 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 4914 4898 5164 5378 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 1944 3798 4044 3968 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal3 1944 5208 4044 5378 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal3 4994 4348 5164 4828 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal3 824 4348 994 4828 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal1 824 208 1464 448 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 824 1548 1464 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 4524 208 5164 448 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 4524 1548 5164 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 824 1218 1064 1788 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 824 208 1064 778 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 4924 208 5164 778 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 4924 1218 5164 1788 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 1944 208 4044 448 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel metal1 1944 1548 4044 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel metal1 824 818 1064 1188 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel metal1 4924 808 5164 1178 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel locali 1474 208 1934 288 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel locali 4054 208 4514 288 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel locali 1474 1708 1934 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel locali 4054 1708 4514 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel metal3 824 208 1464 448 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 4524 208 5164 448 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 824 1548 1464 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 4524 1548 5164 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 824 1308 1074 1788 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 824 208 1074 688 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 4914 208 5164 688 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 4914 1308 5164 1788 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 1944 208 4044 378 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
flabel metal3 1944 1618 4044 1788 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
flabel metal3 4994 758 5164 1238 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
flabel metal3 824 758 994 1238 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
rlabel locali 3680 2796 3680 2834 7 adc_comp_circuit_0/adc_comp_buffer_1/VSS
rlabel locali 3680 2092 3680 2130 7 adc_comp_circuit_0/adc_comp_buffer_1/VDD
rlabel locali 4130 2516 4130 2554 3 adc_comp_circuit_0/adc_comp_buffer_1/out
rlabel poly 3680 2526 3680 2582 7 adc_comp_circuit_0/adc_comp_buffer_1/in
rlabel locali 3680 2826 3680 2864 7 adc_comp_circuit_0/adc_comp_buffer_0/VSS
rlabel locali 3680 3530 3680 3568 7 adc_comp_circuit_0/adc_comp_buffer_0/VDD
rlabel locali 4130 3106 4130 3144 3 adc_comp_circuit_0/adc_comp_buffer_0/out
rlabel poly 3680 3078 3680 3134 7 adc_comp_circuit_0/adc_comp_buffer_0/in
rlabel locali 820 2368 820 2414 7 inverter_0/in
rlabel locali 1054 2368 1054 2414 3 inverter_0/out
rlabel metal1 902 2106 902 2152 7 inverter_0/VSS
rlabel metal1 900 2772 900 2818 7 inverter_0/VDD
rlabel locali 1054 2368 1054 2414 7 inverter_1/in
rlabel locali 1288 2368 1288 2414 3 inverter_1/out
rlabel metal1 1136 2106 1136 2152 7 inverter_1/VSS
rlabel metal1 1134 2772 1134 2818 7 inverter_1/VDD
<< end >>
