magic
tech sky130A
magscale 1 2
timestamp 1665691632
<< nwell >>
rect 111 880 1004 1004
rect 0 506 1004 880
rect 141 499 859 506
<< nmos >>
rect 227 51 271 431
rect 329 51 373 431
rect 431 51 475 431
rect 533 51 577 431
rect 635 51 679 431
rect 737 51 781 431
<< pmos >>
rect 223 588 267 968
rect 325 588 369 968
rect 427 588 471 968
rect 529 588 573 968
rect 631 588 675 968
rect 733 588 777 968
<< ndiff >>
rect 169 419 227 431
rect 169 100 181 419
rect 215 100 227 419
rect 169 51 227 100
rect 271 419 329 431
rect 271 63 283 419
rect 317 63 329 419
rect 271 51 329 63
rect 373 419 431 431
rect 373 63 385 419
rect 419 63 431 419
rect 373 51 431 63
rect 475 419 533 431
rect 475 63 487 419
rect 521 63 533 419
rect 475 51 533 63
rect 577 419 635 431
rect 577 63 589 419
rect 623 63 635 419
rect 577 51 635 63
rect 679 419 737 431
rect 679 63 691 419
rect 725 63 737 419
rect 679 51 737 63
rect 781 419 840 431
rect 781 103 793 419
rect 827 103 840 419
rect 781 51 840 103
<< pdiff >>
rect 170 928 223 968
rect 170 600 178 928
rect 212 600 223 928
rect 170 588 223 600
rect 267 956 325 968
rect 267 600 279 956
rect 313 600 325 956
rect 267 588 325 600
rect 369 956 427 968
rect 369 600 381 956
rect 415 600 427 956
rect 369 588 427 600
rect 471 956 529 968
rect 471 607 483 956
rect 517 607 529 956
rect 471 588 529 607
rect 573 956 631 968
rect 573 600 585 956
rect 619 600 631 956
rect 573 588 631 600
rect 675 956 733 968
rect 675 600 687 956
rect 721 600 733 956
rect 675 588 733 600
rect 777 930 835 968
rect 777 600 789 930
rect 823 600 835 930
rect 777 588 835 600
<< ndiffc >>
rect 181 100 215 419
rect 283 63 317 419
rect 385 63 419 419
rect 487 63 521 419
rect 589 63 623 419
rect 691 63 725 419
rect 793 103 827 419
<< pdiffc >>
rect 178 600 212 928
rect 279 600 313 956
rect 381 600 415 956
rect 483 607 517 956
rect 585 600 619 956
rect 687 600 721 956
rect 789 600 823 930
<< psubdiff >>
rect 895 192 970 216
rect 895 136 903 192
rect 963 136 970 192
rect 895 112 970 136
<< nsubdiff >>
rect 898 832 967 876
rect 898 776 907 832
rect 958 776 967 832
rect 898 720 967 776
<< psubdiffcont >>
rect 903 136 963 192
<< nsubdiffcont >>
rect 907 776 958 832
<< poly >>
rect 223 968 267 994
rect 325 968 369 994
rect 427 968 471 994
rect 529 968 573 994
rect 631 968 675 994
rect 733 968 777 994
rect 223 572 267 588
rect 325 572 369 588
rect 223 528 369 572
rect 427 573 471 588
rect 529 573 573 588
rect 631 573 675 588
rect 733 573 777 588
rect 427 569 777 573
rect 427 543 781 569
rect 223 493 268 528
rect 335 493 369 528
rect 223 476 369 493
rect 631 532 781 543
rect 631 497 683 532
rect 737 497 781 532
rect 223 450 577 476
rect 227 446 577 450
rect 631 447 781 497
rect 227 431 271 446
rect 329 431 373 446
rect 431 431 475 446
rect 533 431 577 446
rect 635 446 781 447
rect 635 431 679 446
rect 737 431 781 446
rect 227 4 271 51
rect 329 4 373 51
rect 431 4 475 51
rect 533 4 577 51
rect 635 4 679 51
rect 737 4 781 51
<< polycont >>
rect 268 493 335 528
rect 683 497 737 532
<< locali >>
rect 34 970 148 1004
rect 34 924 142 970
rect 267 956 323 972
rect 267 953 279 956
rect 34 888 46 924
rect 136 888 142 924
rect 34 706 142 888
rect 34 670 46 706
rect 121 670 142 706
rect 34 610 142 670
rect 34 574 46 610
rect 121 574 142 610
rect 34 266 142 574
rect 178 928 279 953
rect 212 600 279 928
rect 313 709 323 956
rect 370 956 426 972
rect 370 709 381 956
rect 313 647 381 709
rect 313 600 323 647
rect 178 572 323 600
rect 370 600 381 647
rect 415 600 426 956
rect 370 584 426 600
rect 483 956 517 972
rect 483 591 517 607
rect 585 956 619 972
rect 585 584 619 600
rect 687 956 721 972
rect 854 970 970 1004
rect 687 584 721 600
rect 789 930 823 946
rect 857 924 970 970
rect 857 888 866 924
rect 958 888 970 924
rect 857 882 970 888
rect 907 847 958 848
rect 907 760 958 776
rect 789 584 823 600
rect 857 706 970 715
rect 857 670 879 706
rect 958 670 970 706
rect 857 610 970 670
rect 857 574 879 610
rect 958 574 970 610
rect 178 536 218 572
rect 34 232 82 266
rect 116 232 142 266
rect 34 129 142 232
rect 177 419 217 536
rect 252 493 268 528
rect 335 493 351 528
rect 667 497 683 532
rect 737 497 753 532
rect 857 531 970 574
rect 34 102 141 129
rect 34 66 46 102
rect 136 66 141 102
rect 177 100 181 419
rect 215 100 217 419
rect 177 76 217 100
rect 272 419 327 435
rect 34 34 141 66
rect 272 56 283 419
rect 317 56 327 419
rect 272 47 327 56
rect 374 419 430 435
rect 374 63 385 419
rect 419 63 430 419
rect 374 47 430 63
rect 487 419 521 437
rect 487 47 521 56
rect 589 419 623 437
rect 691 419 827 435
rect 623 283 691 345
rect 725 338 793 419
rect 725 300 792 338
rect 589 47 623 63
rect 725 103 793 300
rect 862 340 970 531
rect 862 282 878 340
rect 958 282 970 340
rect 862 230 970 282
rect 887 136 903 192
rect 963 136 979 192
rect 725 86 827 103
rect 691 47 725 63
rect 34 0 148 34
rect 854 0 970 51
<< viali >>
rect 46 888 136 924
rect 46 670 121 706
rect 46 574 121 610
rect 381 657 415 700
rect 483 889 517 927
rect 585 658 619 701
rect 687 888 721 926
rect 866 888 958 924
rect 907 832 958 847
rect 907 804 958 832
rect 789 657 823 700
rect 879 670 958 706
rect 879 574 958 610
rect 82 232 116 266
rect 268 493 335 528
rect 683 497 737 532
rect 46 66 136 102
rect 181 300 215 337
rect 283 63 317 98
rect 283 56 317 63
rect 385 300 419 337
rect 487 63 521 98
rect 487 56 521 63
rect 589 283 623 339
rect 691 300 725 338
rect 792 300 793 338
rect 793 300 826 338
rect 878 282 958 340
rect 903 143 963 185
<< metal1 >>
rect 34 924 148 1004
rect 854 963 970 1004
rect 34 888 46 924
rect 136 888 148 924
rect 34 882 148 888
rect 266 882 272 934
rect 324 927 733 934
rect 324 889 483 927
rect 517 926 733 927
rect 517 889 687 926
rect 324 888 687 889
rect 721 888 733 926
rect 324 882 733 888
rect 854 924 879 963
rect 854 888 866 924
rect 961 888 970 963
rect 854 882 970 888
rect 0 847 1004 854
rect 0 804 907 847
rect 958 804 1004 847
rect 0 798 1004 804
rect 0 740 1004 770
rect 34 706 133 712
rect 34 670 46 706
rect 121 670 133 706
rect 34 610 133 670
rect 347 700 574 707
rect 347 657 381 700
rect 415 657 574 700
rect 630 700 835 707
rect 347 651 574 657
rect 630 657 789 700
rect 823 657 835 700
rect 630 651 835 657
rect 865 706 970 712
rect 865 670 879 706
rect 958 670 970 706
rect 34 574 46 610
rect 121 574 133 610
rect 865 650 970 670
rect 34 568 133 574
rect 161 568 821 600
rect 865 575 876 650
rect 865 574 879 575
rect 958 574 970 650
rect 865 568 970 574
rect 161 540 189 568
rect 790 540 821 568
rect 0 512 189 540
rect 252 528 353 540
rect 252 493 268 528
rect 335 493 353 528
rect 252 487 353 493
rect 405 487 411 540
rect 667 532 701 540
rect 667 497 683 532
rect 667 491 701 497
rect 695 488 701 491
rect 753 488 759 540
rect 790 512 1004 540
rect 0 430 1004 458
rect 0 374 1004 402
rect 169 339 838 345
rect 169 337 578 339
rect 169 300 181 337
rect 215 300 385 337
rect 419 300 578 337
rect 169 294 578 300
rect 572 283 578 294
rect 630 338 838 339
rect 630 300 691 338
rect 725 300 792 338
rect 826 300 838 338
rect 630 294 838 300
rect 866 340 970 346
rect 866 334 878 340
rect 958 334 970 340
rect 630 283 643 294
rect 76 266 122 278
rect 572 277 643 283
rect 866 282 872 334
rect 964 282 970 334
rect 866 276 970 282
rect 76 248 82 266
rect 0 232 82 248
rect 116 248 122 266
rect 116 232 1004 248
rect 0 220 1004 232
rect 0 185 1004 192
rect 0 143 903 185
rect 963 143 1004 185
rect 0 136 1004 143
rect 34 102 148 108
rect 34 66 46 102
rect 136 66 148 102
rect 34 0 148 66
rect 258 56 272 108
rect 324 104 330 108
rect 854 107 970 108
rect 324 98 533 104
rect 324 56 487 98
rect 521 56 533 98
rect 258 47 533 56
rect 854 55 866 107
rect 958 55 970 107
rect 277 0 317 47
rect 854 0 970 55
<< via1 >>
rect 272 882 324 934
rect 879 924 961 963
rect 879 888 958 924
rect 958 888 961 924
rect 574 701 630 707
rect 574 658 585 701
rect 585 658 619 701
rect 619 658 630 701
rect 574 651 630 658
rect 876 610 958 650
rect 876 575 879 610
rect 879 575 958 610
rect 353 487 405 540
rect 701 532 753 540
rect 701 497 737 532
rect 737 497 753 532
rect 701 488 753 497
rect 578 283 589 339
rect 589 283 623 339
rect 623 283 630 339
rect 872 282 878 334
rect 878 282 958 334
rect 958 282 964 334
rect 272 98 324 108
rect 272 56 283 98
rect 283 56 317 98
rect 317 56 324 98
rect 866 55 958 107
<< metal2 >>
rect 32 962 244 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 244 962
rect 352 962 832 972
rect 32 866 244 906
rect 32 810 42 866
rect 98 810 244 866
rect 32 770 244 810
rect 32 714 42 770
rect 98 714 244 770
rect 32 674 244 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 244 674
rect 32 578 244 618
rect 32 522 42 578
rect 98 522 244 578
rect 32 482 244 522
rect 32 426 42 482
rect 98 426 244 482
rect 32 386 244 426
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 244 386
rect 32 290 244 330
rect 32 234 42 290
rect 98 234 244 290
rect 32 194 244 234
rect 32 138 42 194
rect 98 138 244 194
rect 32 98 244 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 244 98
rect 272 934 324 940
rect 272 108 324 882
rect 352 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 832 962
rect 352 866 832 906
rect 352 810 618 866
rect 674 810 832 866
rect 352 745 832 810
rect 352 608 537 745
rect 573 707 631 716
rect 573 642 631 651
rect 665 608 832 745
rect 352 576 832 608
rect 434 572 832 576
rect 272 50 324 56
rect 352 540 406 546
rect 352 487 353 540
rect 405 487 406 540
rect 352 481 406 487
rect 32 32 244 42
rect 352 0 391 481
rect 434 439 664 572
rect 695 488 701 540
rect 753 488 765 540
rect 695 472 765 488
rect 434 379 698 439
rect 434 242 540 379
rect 568 339 639 348
rect 568 283 578 339
rect 634 283 639 339
rect 568 273 639 283
rect 667 242 698 379
rect 434 49 698 242
rect 726 0 765 472
rect 804 513 832 572
rect 865 963 972 972
rect 865 888 879 963
rect 961 888 972 963
rect 865 650 972 888
rect 865 575 876 650
rect 958 575 972 650
rect 865 552 972 575
rect 804 512 833 513
rect 804 482 972 512
rect 804 426 906 482
rect 962 426 972 482
rect 804 416 972 426
rect 861 334 972 359
rect 861 282 872 334
rect 964 282 972 334
rect 861 107 972 282
rect 861 55 866 107
rect 958 55 972 107
rect 861 32 972 55
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 42 810 98 866
rect 42 714 98 770
rect 42 618 98 674
rect 138 618 194 674
rect 42 522 98 578
rect 42 426 98 482
rect 42 330 98 386
rect 138 330 194 386
rect 42 234 98 290
rect 42 138 98 194
rect 42 42 98 98
rect 138 42 194 98
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 618 810 674 866
rect 573 651 574 707
rect 574 651 630 707
rect 630 651 631 707
rect 578 283 630 339
rect 630 283 634 339
rect 906 426 962 482
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 36 680 104 714
rect 324 680 392 900
rect 612 866 680 900
rect 612 810 618 866
rect 674 810 680 866
rect 612 784 680 810
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 36 674 392 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 392 674
rect 558 707 657 724
rect 558 698 573 707
rect 631 698 657 707
rect 558 633 570 698
rect 634 633 657 698
rect 900 680 968 900
rect 558 627 657 633
rect 36 612 392 618
rect 772 612 968 680
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 482 968 612
rect 36 392 104 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 324 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 324 386
rect 36 324 324 330
rect 558 342 645 366
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 558 278 570 342
rect 634 278 645 342
rect 776 324 968 392
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 558 254 645 278
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 36 104 104 138
rect 900 104 968 324
rect 36 98 324 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 324 98
rect 36 36 324 42
rect 692 36 968 104
<< via3 >>
rect 180 756 248 824
rect 756 756 824 824
rect 570 651 573 698
rect 573 651 631 698
rect 631 651 634 698
rect 570 633 634 651
rect 180 468 248 536
rect 756 468 824 536
rect 570 339 634 342
rect 570 283 578 339
rect 578 283 634 339
rect 570 278 634 283
rect 180 180 248 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 248 760 360 820
rect 248 756 264 760
rect 164 740 264 756
rect 184 552 244 740
rect 472 699 532 934
rect 760 840 820 934
rect 740 824 840 840
rect 740 820 756 824
rect 646 760 756 820
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 472 698 635 699
rect 472 633 570 698
rect 634 633 635 698
rect 472 632 635 633
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 468 264 536
rect 164 452 264 468
rect 184 264 244 452
rect 472 344 532 632
rect 760 552 820 740
rect 740 536 840 552
rect 740 468 756 536
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 472 342 635 344
rect 472 278 570 342
rect 634 278 635 342
rect 472 276 635 278
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 180 264 248
rect 164 164 264 180
rect 184 70 244 164
rect 472 48 532 276
rect 760 264 820 452
rect 740 248 840 264
rect 740 180 756 248
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
rlabel metal1 0 740 0 770 7 sample_n
port 2 w
rlabel metal1 0 512 0 540 7 colon_n
port 3 w
rlabel metal1 0 430 0 458 7 col_n
port 4 w
rlabel metal1 0 374 0 402 7 sample
port 5 w
rlabel metal1 0 220 0 248 7 vcom
port 6 w
rlabel metal1 0 136 0 192 7 VSS
port 7 w
rlabel locali 854 0 970 0 5 row_n
port 8 s
rlabel metal1 0 798 0 854 7 VDD
port 13 w
flabel metal1 277 0 317 22 0 FreeSans 64 0 0 0 analog_in
port 16 nsew
flabel metal2 352 0 391 23 0 FreeSans 80 0 0 0 sw
port 17 nsew
flabel metal2 726 0 765 23 0 FreeSans 80 0 0 0 sw_n
port 19 nsew
<< end >>
