* NGSPICE file created from sky130_mm_sc_hd_dlyPoly5ns.ext - technology: sky130A

.subckt sky130_mm_sc_hd_dlyPoly5ns VPWR in out VGND VNB VPB
X0 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.0453e+12p ps=9.52e+06u w=420000u l=3.83e+06u
X1 a_1724_71# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2 VPWR out a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND out a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4 a_1783_329# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 a_1724_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7 a_1783_329# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X8 out cap_top a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10 out cap_top a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
C0 a_1724_71# VGND 0.48fF
C1 cap_top out 0.05fF
C2 cap_top a_1783_329# 0.03fF
C3 cap_top VPB 0.17fF
C4 cap_top in 0.15fF
C5 a_1724_71# VPWR 0.05fF
C6 cap_top VGND 1.77fF
C7 a_1783_329# out 0.04fF
C8 VPB out 0.05fF
C9 out in 0.00fF
C10 VPB a_1783_329# 0.02fF
C11 a_1783_329# in 0.00fF
C12 out VGND 0.09fF
C13 VPB in 0.23fF
C14 a_1783_329# VGND 0.29fF
C15 cap_top VPWR 0.42fF
C16 VPB VGND 0.15fF
C17 VGND in 0.33fF
C18 cap_top a_1724_71# 0.07fF
C19 out VPWR 0.17fF
C20 a_1724_71# out 0.08fF
C21 a_1783_329# VPWR 0.52fF
C22 a_1724_71# a_1783_329# 0.00fF
C23 VPB VPWR 0.28fF
C24 VPWR in 0.20fF
C25 a_1724_71# VPB 0.00fF
C26 a_1724_71# in 0.00fF
C27 VGND VPWR 0.31fF
.ends

