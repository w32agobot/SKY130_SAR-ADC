* SPICE3 file created from adc_array_wafflecap_8(2)x557aF_25um2.ext - technology: sky130A

.subckt adc_array_wafflecap_8(2)x557aF_25um2 cbot ctop
C0 ctop nc 0.26fF
C1 nc cbot 3.26fF
C2 ctop cbot 1.13fF
C3 cbot VSUBS 2.01fF
C4 nc VSUBS 0.41fF
.ends
