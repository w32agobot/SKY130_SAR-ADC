* SPICE3 file created from Extract.ext - technology: sky130A

C0 cbot_2 ctop_dummy 2.54fF
C1 cbot_1 ctop_1_floating 8.18fF
C2 ctop_dummy ctop_16 4.22fF
C3 cbot_2 ctop_2 56.42fF
C4 ctop_2 ctop_dummy 3.77fF
C5 cdummy_bot ctop_1 2.20fF
C6 cbot_8 ctop_8_floating 4.27fF
C7 ctop_dummy cbot_4 2.55fF
C8 cbot_8 ctop_dummy 2.55fF
C9 cdummy_bot cbot_1 23.53fF
C10 cbot_1 ctop_1 55.85fF
C11 ctop_4 cdummy_bot 2.29fF
C12 ctop_8 ctop_dummy 4.17fF
C13 cbot_8 ctop_8 59.74fF
C14 cbot_16 ctop_16 54.98fF
C15 cdummy_bot cbot_2 23.52fF
C16 cdummy_bot ctop_16 2.41fF
C17 cbot_16 ctop_dummy 2.38fF
C18 cdummy_bot ctop_dummy 600.79fF
C19 cdummy_bot ctop_2 2.23fF
C20 cbot_2 ctop_2_floating 7.62fF
C21 cdummy_bot cbot_4 23.53fF
C22 ctop_dummy ctop_1 3.77fF
C23 cdummy_bot cbot_8 23.53fF
C24 cbot_1 ctop_dummy 2.54fF
C25 cbot_4 ctop_4_floating 6.52fF
C26 ctop_4 ctop_dummy 3.97fF
C27 cdummy_bot ctop_8 2.41fF
C28 ctop_4 cbot_4 57.53fF
C29 cdummy_bot cbot_16 21.48fF
C30 cbot_2 VSUBS 5.62fF
C31 cbot_4 VSUBS 5.62fF
C32 cbot_8 VSUBS 5.62fF
C33 cdummy_bot VSUBS 76.82fF
C34 cbot_16 VSUBS 4.36fF
C35 cbot_1 VSUBS 5.62fF
