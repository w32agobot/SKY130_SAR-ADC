magic
tech sky130A
magscale 1 2
timestamp 1666970908
<< psubdiff >>
rect 35396 19655 35810 19862
rect 36540 19692 36954 19900
rect 1046 18357 1460 19462
rect 1046 18356 1169 18357
rect 1046 18298 1074 18356
rect 1130 18299 1169 18356
rect 1225 18356 1460 18357
rect 1225 18299 1278 18356
rect 1130 18298 1278 18299
rect 1334 18298 1373 18356
rect 1429 18298 1460 18356
rect 1046 18147 1460 18298
rect 1046 18146 1169 18147
rect 1046 18088 1074 18146
rect 1130 18089 1169 18146
rect 1225 18146 1460 18147
rect 1225 18089 1278 18146
rect 1130 18088 1278 18089
rect 1334 18088 1373 18146
rect 1429 18088 1460 18146
rect 1046 17144 1460 18088
rect 1046 17143 1169 17144
rect 1046 17085 1074 17143
rect 1130 17086 1169 17143
rect 1225 17143 1460 17144
rect 1225 17086 1278 17143
rect 1130 17085 1278 17086
rect 1334 17085 1373 17143
rect 1429 17085 1460 17143
rect 1046 16139 1460 17085
rect 1046 16138 1169 16139
rect 1046 16080 1074 16138
rect 1130 16081 1169 16138
rect 1225 16138 1460 16139
rect 1225 16081 1278 16138
rect 1130 16080 1278 16081
rect 1334 16080 1373 16138
rect 1429 16080 1460 16138
rect 1046 15136 1460 16080
rect 1046 15135 1169 15136
rect 1046 15077 1074 15135
rect 1130 15078 1169 15135
rect 1225 15135 1460 15136
rect 1225 15078 1278 15135
rect 1130 15077 1278 15078
rect 1334 15077 1373 15135
rect 1429 15077 1460 15135
rect 1046 14132 1460 15077
rect 1046 14131 1169 14132
rect 1046 14073 1074 14131
rect 1130 14074 1169 14131
rect 1225 14131 1460 14132
rect 1225 14074 1278 14131
rect 1130 14073 1278 14074
rect 1334 14073 1373 14131
rect 1429 14073 1460 14131
rect 1046 13128 1460 14073
rect 1046 13127 1169 13128
rect 1046 13069 1074 13127
rect 1130 13070 1169 13127
rect 1225 13127 1460 13128
rect 1225 13070 1278 13127
rect 1130 13069 1278 13070
rect 1334 13069 1373 13127
rect 1429 13069 1460 13127
rect 1046 12124 1460 13069
rect 1046 12123 1169 12124
rect 1046 12065 1074 12123
rect 1130 12066 1169 12123
rect 1225 12123 1460 12124
rect 1225 12066 1278 12123
rect 1130 12065 1278 12066
rect 1334 12065 1373 12123
rect 1429 12065 1460 12123
rect 1046 11120 1460 12065
rect 1046 11119 1169 11120
rect 1046 11061 1074 11119
rect 1130 11062 1169 11119
rect 1225 11119 1460 11120
rect 1225 11062 1278 11119
rect 1130 11061 1278 11062
rect 1334 11061 1373 11119
rect 1429 11061 1460 11119
rect 1046 10116 1460 11061
rect 1046 10115 1169 10116
rect 1046 10057 1074 10115
rect 1130 10058 1169 10115
rect 1225 10115 1460 10116
rect 1225 10058 1278 10115
rect 1130 10057 1278 10058
rect 1334 10057 1373 10115
rect 1429 10057 1460 10115
rect 1046 9112 1460 10057
rect 1046 9111 1169 9112
rect 1046 9053 1074 9111
rect 1130 9054 1169 9111
rect 1225 9111 1460 9112
rect 1225 9054 1278 9111
rect 1130 9053 1278 9054
rect 1334 9053 1373 9111
rect 1429 9053 1460 9111
rect 1046 8108 1460 9053
rect 1046 8107 1169 8108
rect 1046 8049 1074 8107
rect 1130 8050 1169 8107
rect 1225 8107 1460 8108
rect 1225 8050 1278 8107
rect 1130 8049 1278 8050
rect 1334 8049 1373 8107
rect 1429 8049 1460 8107
rect 1046 7104 1460 8049
rect 1046 7103 1169 7104
rect 1046 7045 1074 7103
rect 1130 7046 1169 7103
rect 1225 7103 1460 7104
rect 1225 7046 1278 7103
rect 1130 7045 1278 7046
rect 1334 7045 1373 7103
rect 1429 7045 1460 7103
rect 1046 6100 1460 7045
rect 1046 6099 1169 6100
rect 1046 6041 1074 6099
rect 1130 6042 1169 6099
rect 1225 6099 1460 6100
rect 1225 6042 1278 6099
rect 1130 6041 1278 6042
rect 1334 6041 1373 6099
rect 1429 6041 1460 6099
rect 1046 5096 1460 6041
rect 1046 5095 1169 5096
rect 1046 5037 1074 5095
rect 1130 5038 1169 5095
rect 1225 5095 1460 5096
rect 1225 5038 1278 5095
rect 1130 5037 1278 5038
rect 1334 5037 1373 5095
rect 1429 5037 1460 5095
rect 1046 4092 1460 5037
rect 1046 4091 1169 4092
rect 1046 4033 1074 4091
rect 1130 4034 1169 4091
rect 1225 4091 1460 4092
rect 1225 4034 1278 4091
rect 1130 4033 1278 4034
rect 1334 4033 1373 4091
rect 1429 4033 1460 4091
rect 1046 3086 1460 4033
rect 1046 3085 1169 3086
rect 1046 3027 1074 3085
rect 1130 3028 1169 3085
rect 1225 3085 1460 3086
rect 1225 3028 1278 3085
rect 1130 3027 1278 3028
rect 1334 3027 1373 3085
rect 1429 3027 1460 3085
rect 1046 2083 1460 3027
rect 1046 2082 1169 2083
rect 1046 2024 1074 2082
rect 1130 2025 1169 2082
rect 1225 2082 1460 2083
rect 1225 2025 1278 2082
rect 1130 2024 1278 2025
rect 1334 2024 1373 2082
rect 1429 2024 1460 2082
rect 1046 1428 1460 2024
rect 1046 1427 1169 1428
rect 1046 1369 1074 1427
rect 1130 1370 1169 1427
rect 1225 1427 1460 1428
rect 1225 1370 1278 1427
rect 1130 1369 1278 1370
rect 1334 1369 1373 1427
rect 1429 1369 1460 1427
rect 1046 1318 1460 1369
rect 1046 1317 1169 1318
rect 1046 1259 1074 1317
rect 1130 1260 1169 1317
rect 1225 1317 1460 1318
rect 1225 1260 1278 1317
rect 1130 1259 1278 1260
rect 1334 1259 1373 1317
rect 1429 1259 1460 1317
rect 1046 1079 1460 1259
rect 1046 1078 1169 1079
rect 1046 1020 1074 1078
rect 1130 1021 1169 1078
rect 1225 1078 1460 1079
rect 1225 1021 1278 1078
rect 1130 1020 1278 1021
rect 1334 1020 1373 1078
rect 1429 1020 1460 1078
rect 1046 480 1460 1020
rect 36064 18662 36478 19585
rect 36064 18380 36480 18662
rect 36064 18148 36478 18380
rect 36064 18147 36187 18148
rect 36064 18089 36092 18147
rect 36148 18090 36187 18147
rect 36243 18147 36478 18148
rect 36243 18090 36296 18147
rect 36148 18089 36296 18090
rect 36352 18089 36391 18147
rect 36447 18089 36478 18147
rect 36064 17144 36478 18089
rect 36064 17143 36187 17144
rect 36064 17085 36092 17143
rect 36148 17086 36187 17143
rect 36243 17143 36478 17144
rect 36243 17086 36296 17143
rect 36148 17085 36296 17086
rect 36352 17085 36391 17143
rect 36447 17085 36478 17143
rect 36064 16140 36478 17085
rect 36064 16139 36187 16140
rect 36064 16081 36092 16139
rect 36148 16082 36187 16139
rect 36243 16139 36478 16140
rect 36243 16082 36296 16139
rect 36148 16081 36296 16082
rect 36352 16081 36391 16139
rect 36447 16081 36478 16139
rect 36064 15136 36478 16081
rect 36064 15135 36187 15136
rect 36064 15077 36092 15135
rect 36148 15078 36187 15135
rect 36243 15135 36478 15136
rect 36243 15078 36296 15135
rect 36148 15077 36296 15078
rect 36352 15077 36391 15135
rect 36447 15077 36478 15135
rect 36064 14132 36478 15077
rect 36064 14131 36187 14132
rect 36064 14073 36092 14131
rect 36148 14074 36187 14131
rect 36243 14131 36478 14132
rect 36243 14074 36296 14131
rect 36148 14073 36296 14074
rect 36352 14073 36391 14131
rect 36447 14073 36478 14131
rect 36064 13128 36478 14073
rect 36064 13127 36187 13128
rect 36064 13069 36092 13127
rect 36148 13070 36187 13127
rect 36243 13127 36478 13128
rect 36243 13070 36296 13127
rect 36148 13069 36296 13070
rect 36352 13069 36391 13127
rect 36447 13069 36478 13127
rect 36064 12124 36478 13069
rect 36064 12123 36187 12124
rect 36064 12065 36092 12123
rect 36148 12066 36187 12123
rect 36243 12123 36478 12124
rect 36243 12066 36296 12123
rect 36148 12065 36296 12066
rect 36352 12065 36391 12123
rect 36447 12065 36478 12123
rect 36064 11120 36478 12065
rect 36064 11119 36187 11120
rect 36064 11061 36092 11119
rect 36148 11062 36187 11119
rect 36243 11119 36478 11120
rect 36243 11062 36296 11119
rect 36148 11061 36296 11062
rect 36352 11061 36391 11119
rect 36447 11061 36478 11119
rect 36064 10116 36478 11061
rect 36064 10115 36187 10116
rect 36064 10057 36092 10115
rect 36148 10058 36187 10115
rect 36243 10115 36478 10116
rect 36243 10058 36296 10115
rect 36148 10057 36296 10058
rect 36352 10057 36391 10115
rect 36447 10057 36478 10115
rect 36064 9112 36478 10057
rect 36064 9111 36187 9112
rect 36064 9053 36092 9111
rect 36148 9054 36187 9111
rect 36243 9111 36478 9112
rect 36243 9054 36296 9111
rect 36148 9053 36296 9054
rect 36352 9053 36391 9111
rect 36447 9053 36478 9111
rect 36064 8108 36478 9053
rect 36064 8107 36187 8108
rect 36064 8049 36092 8107
rect 36148 8050 36187 8107
rect 36243 8107 36478 8108
rect 36243 8050 36296 8107
rect 36148 8049 36296 8050
rect 36352 8049 36391 8107
rect 36447 8049 36478 8107
rect 36064 7104 36478 8049
rect 36064 7103 36187 7104
rect 36064 7045 36092 7103
rect 36148 7046 36187 7103
rect 36243 7103 36478 7104
rect 36243 7046 36296 7103
rect 36148 7045 36296 7046
rect 36352 7045 36391 7103
rect 36447 7045 36478 7103
rect 36064 6576 36478 7045
rect 36064 6294 36480 6576
rect 36064 6100 36478 6294
rect 36064 6099 36187 6100
rect 36064 6041 36092 6099
rect 36148 6042 36187 6099
rect 36243 6099 36478 6100
rect 36243 6042 36296 6099
rect 36148 6041 36296 6042
rect 36352 6041 36391 6099
rect 36447 6041 36478 6099
rect 36064 5096 36478 6041
rect 36064 5095 36187 5096
rect 36064 5037 36092 5095
rect 36148 5038 36187 5095
rect 36243 5095 36478 5096
rect 36243 5038 36296 5095
rect 36148 5037 36296 5038
rect 36352 5037 36391 5095
rect 36447 5037 36478 5095
rect 36064 4092 36478 5037
rect 36064 4091 36187 4092
rect 36064 4033 36092 4091
rect 36148 4034 36187 4091
rect 36243 4091 36478 4092
rect 36243 4034 36296 4091
rect 36148 4033 36296 4034
rect 36352 4033 36391 4091
rect 36447 4033 36478 4091
rect 36064 3088 36478 4033
rect 36064 3087 36187 3088
rect 36064 3029 36092 3087
rect 36148 3030 36187 3087
rect 36243 3087 36478 3088
rect 36243 3030 36296 3087
rect 36148 3029 36296 3030
rect 36352 3029 36391 3087
rect 36447 3029 36478 3087
rect 36064 2084 36478 3029
rect 36064 2083 36187 2084
rect 36064 2025 36092 2083
rect 36148 2026 36187 2083
rect 36243 2083 36478 2084
rect 36243 2026 36296 2083
rect 36148 2025 36296 2026
rect 36352 2025 36391 2083
rect 36447 2025 36478 2083
rect 36064 1080 36478 2025
rect 36064 1079 36187 1080
rect 36064 1021 36092 1079
rect 36148 1022 36187 1079
rect 36243 1079 36478 1080
rect 36243 1022 36296 1079
rect 36148 1021 36296 1022
rect 36352 1021 36391 1079
rect 36447 1021 36478 1079
rect 36064 610 36478 1021
<< psubdiffcont >>
rect 1074 18298 1130 18356
rect 1169 18299 1225 18357
rect 1278 18298 1334 18356
rect 1373 18298 1429 18356
rect 1074 18088 1130 18146
rect 1169 18089 1225 18147
rect 1278 18088 1334 18146
rect 1373 18088 1429 18146
rect 1074 17085 1130 17143
rect 1169 17086 1225 17144
rect 1278 17085 1334 17143
rect 1373 17085 1429 17143
rect 1074 16080 1130 16138
rect 1169 16081 1225 16139
rect 1278 16080 1334 16138
rect 1373 16080 1429 16138
rect 1074 15077 1130 15135
rect 1169 15078 1225 15136
rect 1278 15077 1334 15135
rect 1373 15077 1429 15135
rect 1074 14073 1130 14131
rect 1169 14074 1225 14132
rect 1278 14073 1334 14131
rect 1373 14073 1429 14131
rect 1074 13069 1130 13127
rect 1169 13070 1225 13128
rect 1278 13069 1334 13127
rect 1373 13069 1429 13127
rect 1074 12065 1130 12123
rect 1169 12066 1225 12124
rect 1278 12065 1334 12123
rect 1373 12065 1429 12123
rect 1074 11061 1130 11119
rect 1169 11062 1225 11120
rect 1278 11061 1334 11119
rect 1373 11061 1429 11119
rect 1074 10057 1130 10115
rect 1169 10058 1225 10116
rect 1278 10057 1334 10115
rect 1373 10057 1429 10115
rect 1074 9053 1130 9111
rect 1169 9054 1225 9112
rect 1278 9053 1334 9111
rect 1373 9053 1429 9111
rect 1074 8049 1130 8107
rect 1169 8050 1225 8108
rect 1278 8049 1334 8107
rect 1373 8049 1429 8107
rect 1074 7045 1130 7103
rect 1169 7046 1225 7104
rect 1278 7045 1334 7103
rect 1373 7045 1429 7103
rect 1074 6041 1130 6099
rect 1169 6042 1225 6100
rect 1278 6041 1334 6099
rect 1373 6041 1429 6099
rect 1074 5037 1130 5095
rect 1169 5038 1225 5096
rect 1278 5037 1334 5095
rect 1373 5037 1429 5095
rect 1074 4033 1130 4091
rect 1169 4034 1225 4092
rect 1278 4033 1334 4091
rect 1373 4033 1429 4091
rect 1074 3027 1130 3085
rect 1169 3028 1225 3086
rect 1278 3027 1334 3085
rect 1373 3027 1429 3085
rect 1074 2024 1130 2082
rect 1169 2025 1225 2083
rect 1278 2024 1334 2082
rect 1373 2024 1429 2082
rect 1074 1369 1130 1427
rect 1169 1370 1225 1428
rect 1278 1369 1334 1427
rect 1373 1369 1429 1427
rect 1074 1259 1130 1317
rect 1169 1260 1225 1318
rect 1278 1259 1334 1317
rect 1373 1259 1429 1317
rect 1074 1020 1130 1078
rect 1169 1021 1225 1079
rect 1278 1020 1334 1078
rect 1373 1020 1429 1078
rect 36092 18089 36148 18147
rect 36187 18090 36243 18148
rect 36296 18089 36352 18147
rect 36391 18089 36447 18147
rect 36092 17085 36148 17143
rect 36187 17086 36243 17144
rect 36296 17085 36352 17143
rect 36391 17085 36447 17143
rect 36092 16081 36148 16139
rect 36187 16082 36243 16140
rect 36296 16081 36352 16139
rect 36391 16081 36447 16139
rect 36092 15077 36148 15135
rect 36187 15078 36243 15136
rect 36296 15077 36352 15135
rect 36391 15077 36447 15135
rect 36092 14073 36148 14131
rect 36187 14074 36243 14132
rect 36296 14073 36352 14131
rect 36391 14073 36447 14131
rect 36092 13069 36148 13127
rect 36187 13070 36243 13128
rect 36296 13069 36352 13127
rect 36391 13069 36447 13127
rect 36092 12065 36148 12123
rect 36187 12066 36243 12124
rect 36296 12065 36352 12123
rect 36391 12065 36447 12123
rect 36092 11061 36148 11119
rect 36187 11062 36243 11120
rect 36296 11061 36352 11119
rect 36391 11061 36447 11119
rect 36092 10057 36148 10115
rect 36187 10058 36243 10116
rect 36296 10057 36352 10115
rect 36391 10057 36447 10115
rect 36092 9053 36148 9111
rect 36187 9054 36243 9112
rect 36296 9053 36352 9111
rect 36391 9053 36447 9111
rect 36092 8049 36148 8107
rect 36187 8050 36243 8108
rect 36296 8049 36352 8107
rect 36391 8049 36447 8107
rect 36092 7045 36148 7103
rect 36187 7046 36243 7104
rect 36296 7045 36352 7103
rect 36391 7045 36447 7103
rect 36092 6041 36148 6099
rect 36187 6042 36243 6100
rect 36296 6041 36352 6099
rect 36391 6041 36447 6099
rect 36092 5037 36148 5095
rect 36187 5038 36243 5096
rect 36296 5037 36352 5095
rect 36391 5037 36447 5095
rect 36092 4033 36148 4091
rect 36187 4034 36243 4092
rect 36296 4033 36352 4091
rect 36391 4033 36447 4091
rect 36092 3029 36148 3087
rect 36187 3030 36243 3088
rect 36296 3029 36352 3087
rect 36391 3029 36447 3087
rect 36092 2025 36148 2083
rect 36187 2026 36243 2084
rect 36296 2025 36352 2083
rect 36391 2025 36447 2083
rect 36092 1021 36148 1079
rect 36187 1022 36243 1080
rect 36296 1021 36352 1079
rect 36391 1021 36447 1079
<< locali >>
rect 41602 23250 42660 23276
rect 41602 22838 42422 23250
rect 42634 22838 42660 23250
rect 41602 22814 42660 22838
rect 41602 21492 42660 21518
rect 41602 21080 42422 21492
rect 42634 21080 42660 21492
rect 41602 21056 42660 21080
rect 1884 20104 2176 20120
rect 1884 19946 1898 20104
rect 2160 19946 2176 20104
rect 1884 19442 2176 19946
rect 1884 19386 1904 19442
rect 1960 19386 1998 19442
rect 2054 19386 2092 19442
rect 2148 19386 2176 19442
rect 1884 19348 2176 19386
rect 1884 19292 1904 19348
rect 1960 19292 1998 19348
rect 2054 19292 2092 19348
rect 2148 19292 2176 19348
rect 1884 19254 2176 19292
rect 1884 19198 1904 19254
rect 1960 19198 1998 19254
rect 2054 19198 2092 19254
rect 2148 19198 2176 19254
rect 1884 19182 2176 19198
rect 2584 19442 2876 20166
rect 2584 19386 2604 19442
rect 2660 19386 2698 19442
rect 2754 19386 2792 19442
rect 2848 19386 2876 19442
rect 2584 19348 2876 19386
rect 2584 19292 2604 19348
rect 2660 19292 2698 19348
rect 2754 19292 2792 19348
rect 2848 19292 2876 19348
rect 2584 19254 2876 19292
rect 2584 19198 2604 19254
rect 2660 19198 2698 19254
rect 2754 19198 2792 19254
rect 2848 19198 2876 19254
rect 2584 19182 2876 19198
rect 5012 20104 5304 20120
rect 5012 19946 5026 20104
rect 5288 19946 5304 20104
rect 5012 19442 5304 19946
rect 5012 19386 5032 19442
rect 5088 19386 5126 19442
rect 5182 19386 5220 19442
rect 5276 19386 5304 19442
rect 5012 19348 5304 19386
rect 5012 19292 5032 19348
rect 5088 19292 5126 19348
rect 5182 19292 5220 19348
rect 5276 19292 5304 19348
rect 5012 19254 5304 19292
rect 5012 19198 5032 19254
rect 5088 19198 5126 19254
rect 5182 19198 5220 19254
rect 5276 19198 5304 19254
rect 5012 19182 5304 19198
rect 5884 20104 6176 20120
rect 5884 19946 5898 20104
rect 6160 19946 6176 20104
rect 5884 19442 6176 19946
rect 5884 19386 5904 19442
rect 5960 19386 5998 19442
rect 6054 19386 6092 19442
rect 6148 19386 6176 19442
rect 5884 19348 6176 19386
rect 5884 19292 5904 19348
rect 5960 19292 5998 19348
rect 6054 19292 6092 19348
rect 6148 19292 6176 19348
rect 5884 19254 6176 19292
rect 5884 19198 5904 19254
rect 5960 19198 5998 19254
rect 6054 19198 6092 19254
rect 6148 19198 6176 19254
rect 5884 19182 6176 19198
rect 6584 19442 6876 20166
rect 6584 19386 6604 19442
rect 6660 19386 6698 19442
rect 6754 19386 6792 19442
rect 6848 19386 6876 19442
rect 6584 19348 6876 19386
rect 6584 19292 6604 19348
rect 6660 19292 6698 19348
rect 6754 19292 6792 19348
rect 6848 19292 6876 19348
rect 6584 19254 6876 19292
rect 6584 19198 6604 19254
rect 6660 19198 6698 19254
rect 6754 19198 6792 19254
rect 6848 19198 6876 19254
rect 6584 19182 6876 19198
rect 9012 20104 9304 20120
rect 9012 19946 9026 20104
rect 9288 19946 9304 20104
rect 9012 19442 9304 19946
rect 9012 19386 9032 19442
rect 9088 19386 9126 19442
rect 9182 19386 9220 19442
rect 9276 19386 9304 19442
rect 9012 19348 9304 19386
rect 9012 19292 9032 19348
rect 9088 19292 9126 19348
rect 9182 19292 9220 19348
rect 9276 19292 9304 19348
rect 9012 19254 9304 19292
rect 9012 19198 9032 19254
rect 9088 19198 9126 19254
rect 9182 19198 9220 19254
rect 9276 19198 9304 19254
rect 9012 19182 9304 19198
rect 9884 20104 10176 20120
rect 9884 19946 9898 20104
rect 10160 19946 10176 20104
rect 9884 19442 10176 19946
rect 9884 19386 9904 19442
rect 9960 19386 9998 19442
rect 10054 19386 10092 19442
rect 10148 19386 10176 19442
rect 9884 19348 10176 19386
rect 9884 19292 9904 19348
rect 9960 19292 9998 19348
rect 10054 19292 10092 19348
rect 10148 19292 10176 19348
rect 9884 19254 10176 19292
rect 9884 19198 9904 19254
rect 9960 19198 9998 19254
rect 10054 19198 10092 19254
rect 10148 19198 10176 19254
rect 9884 19182 10176 19198
rect 10584 19442 10876 20166
rect 10584 19386 10604 19442
rect 10660 19386 10698 19442
rect 10754 19386 10792 19442
rect 10848 19386 10876 19442
rect 10584 19348 10876 19386
rect 10584 19292 10604 19348
rect 10660 19292 10698 19348
rect 10754 19292 10792 19348
rect 10848 19292 10876 19348
rect 10584 19254 10876 19292
rect 10584 19198 10604 19254
rect 10660 19198 10698 19254
rect 10754 19198 10792 19254
rect 10848 19198 10876 19254
rect 10584 19182 10876 19198
rect 13012 20104 13304 20120
rect 13012 19946 13026 20104
rect 13288 19946 13304 20104
rect 13012 19442 13304 19946
rect 13012 19386 13032 19442
rect 13088 19386 13126 19442
rect 13182 19386 13220 19442
rect 13276 19386 13304 19442
rect 13012 19348 13304 19386
rect 13012 19292 13032 19348
rect 13088 19292 13126 19348
rect 13182 19292 13220 19348
rect 13276 19292 13304 19348
rect 13012 19254 13304 19292
rect 13012 19198 13032 19254
rect 13088 19198 13126 19254
rect 13182 19198 13220 19254
rect 13276 19198 13304 19254
rect 13012 19182 13304 19198
rect 13884 20104 14176 20120
rect 13884 19946 13898 20104
rect 14160 19946 14176 20104
rect 13884 19442 14176 19946
rect 13884 19386 13904 19442
rect 13960 19386 13998 19442
rect 14054 19386 14092 19442
rect 14148 19386 14176 19442
rect 13884 19348 14176 19386
rect 13884 19292 13904 19348
rect 13960 19292 13998 19348
rect 14054 19292 14092 19348
rect 14148 19292 14176 19348
rect 13884 19254 14176 19292
rect 13884 19198 13904 19254
rect 13960 19198 13998 19254
rect 14054 19198 14092 19254
rect 14148 19198 14176 19254
rect 13884 19182 14176 19198
rect 14584 19442 14876 20166
rect 14584 19386 14604 19442
rect 14660 19386 14698 19442
rect 14754 19386 14792 19442
rect 14848 19386 14876 19442
rect 14584 19348 14876 19386
rect 14584 19292 14604 19348
rect 14660 19292 14698 19348
rect 14754 19292 14792 19348
rect 14848 19292 14876 19348
rect 14584 19254 14876 19292
rect 14584 19198 14604 19254
rect 14660 19198 14698 19254
rect 14754 19198 14792 19254
rect 14848 19198 14876 19254
rect 14584 19182 14876 19198
rect 17012 20104 17304 20120
rect 17012 19946 17026 20104
rect 17288 19946 17304 20104
rect 17012 19442 17304 19946
rect 17012 19386 17032 19442
rect 17088 19386 17126 19442
rect 17182 19386 17220 19442
rect 17276 19386 17304 19442
rect 17012 19348 17304 19386
rect 17012 19292 17032 19348
rect 17088 19292 17126 19348
rect 17182 19292 17220 19348
rect 17276 19292 17304 19348
rect 17012 19254 17304 19292
rect 17012 19198 17032 19254
rect 17088 19198 17126 19254
rect 17182 19198 17220 19254
rect 17276 19198 17304 19254
rect 17012 19182 17304 19198
rect 17884 20104 18176 20120
rect 17884 19946 17898 20104
rect 18160 19946 18176 20104
rect 17884 19442 18176 19946
rect 17884 19386 17904 19442
rect 17960 19386 17998 19442
rect 18054 19386 18092 19442
rect 18148 19386 18176 19442
rect 17884 19348 18176 19386
rect 17884 19292 17904 19348
rect 17960 19292 17998 19348
rect 18054 19292 18092 19348
rect 18148 19292 18176 19348
rect 17884 19254 18176 19292
rect 17884 19198 17904 19254
rect 17960 19198 17998 19254
rect 18054 19198 18092 19254
rect 18148 19198 18176 19254
rect 17884 19182 18176 19198
rect 18584 19442 18876 20166
rect 18584 19386 18604 19442
rect 18660 19386 18698 19442
rect 18754 19386 18792 19442
rect 18848 19386 18876 19442
rect 18584 19348 18876 19386
rect 18584 19292 18604 19348
rect 18660 19292 18698 19348
rect 18754 19292 18792 19348
rect 18848 19292 18876 19348
rect 18584 19254 18876 19292
rect 18584 19198 18604 19254
rect 18660 19198 18698 19254
rect 18754 19198 18792 19254
rect 18848 19198 18876 19254
rect 18584 19182 18876 19198
rect 21012 20104 21304 20120
rect 21012 19946 21026 20104
rect 21288 19946 21304 20104
rect 21012 19442 21304 19946
rect 21012 19386 21032 19442
rect 21088 19386 21126 19442
rect 21182 19386 21220 19442
rect 21276 19386 21304 19442
rect 21012 19348 21304 19386
rect 21012 19292 21032 19348
rect 21088 19292 21126 19348
rect 21182 19292 21220 19348
rect 21276 19292 21304 19348
rect 21012 19254 21304 19292
rect 21012 19198 21032 19254
rect 21088 19198 21126 19254
rect 21182 19198 21220 19254
rect 21276 19198 21304 19254
rect 21012 19182 21304 19198
rect 21884 20104 22176 20120
rect 21884 19946 21898 20104
rect 22160 19946 22176 20104
rect 21884 19442 22176 19946
rect 21884 19386 21904 19442
rect 21960 19386 21998 19442
rect 22054 19386 22092 19442
rect 22148 19386 22176 19442
rect 21884 19348 22176 19386
rect 21884 19292 21904 19348
rect 21960 19292 21998 19348
rect 22054 19292 22092 19348
rect 22148 19292 22176 19348
rect 21884 19254 22176 19292
rect 21884 19198 21904 19254
rect 21960 19198 21998 19254
rect 22054 19198 22092 19254
rect 22148 19198 22176 19254
rect 21884 19182 22176 19198
rect 22584 19442 22876 20166
rect 22584 19386 22604 19442
rect 22660 19386 22698 19442
rect 22754 19386 22792 19442
rect 22848 19386 22876 19442
rect 22584 19348 22876 19386
rect 22584 19292 22604 19348
rect 22660 19292 22698 19348
rect 22754 19292 22792 19348
rect 22848 19292 22876 19348
rect 22584 19254 22876 19292
rect 22584 19198 22604 19254
rect 22660 19198 22698 19254
rect 22754 19198 22792 19254
rect 22848 19198 22876 19254
rect 22584 19182 22876 19198
rect 25012 20104 25304 20120
rect 25012 19946 25026 20104
rect 25288 19946 25304 20104
rect 25012 19442 25304 19946
rect 25012 19386 25032 19442
rect 25088 19386 25126 19442
rect 25182 19386 25220 19442
rect 25276 19386 25304 19442
rect 25012 19348 25304 19386
rect 25012 19292 25032 19348
rect 25088 19292 25126 19348
rect 25182 19292 25220 19348
rect 25276 19292 25304 19348
rect 25012 19254 25304 19292
rect 25012 19198 25032 19254
rect 25088 19198 25126 19254
rect 25182 19198 25220 19254
rect 25276 19198 25304 19254
rect 25012 19182 25304 19198
rect 25884 20104 26176 20120
rect 25884 19946 25898 20104
rect 26160 19946 26176 20104
rect 25884 19442 26176 19946
rect 25884 19386 25904 19442
rect 25960 19386 25998 19442
rect 26054 19386 26092 19442
rect 26148 19386 26176 19442
rect 25884 19348 26176 19386
rect 25884 19292 25904 19348
rect 25960 19292 25998 19348
rect 26054 19292 26092 19348
rect 26148 19292 26176 19348
rect 25884 19254 26176 19292
rect 25884 19198 25904 19254
rect 25960 19198 25998 19254
rect 26054 19198 26092 19254
rect 26148 19198 26176 19254
rect 25884 19182 26176 19198
rect 26584 19442 26876 20166
rect 26584 19386 26604 19442
rect 26660 19386 26698 19442
rect 26754 19386 26792 19442
rect 26848 19386 26876 19442
rect 26584 19348 26876 19386
rect 26584 19292 26604 19348
rect 26660 19292 26698 19348
rect 26754 19292 26792 19348
rect 26848 19292 26876 19348
rect 26584 19254 26876 19292
rect 26584 19198 26604 19254
rect 26660 19198 26698 19254
rect 26754 19198 26792 19254
rect 26848 19198 26876 19254
rect 26584 19182 26876 19198
rect 29012 20104 29304 20120
rect 29012 19946 29026 20104
rect 29288 19946 29304 20104
rect 29012 19442 29304 19946
rect 29012 19386 29032 19442
rect 29088 19386 29126 19442
rect 29182 19386 29220 19442
rect 29276 19386 29304 19442
rect 29012 19348 29304 19386
rect 29012 19292 29032 19348
rect 29088 19292 29126 19348
rect 29182 19292 29220 19348
rect 29276 19292 29304 19348
rect 29012 19254 29304 19292
rect 29012 19198 29032 19254
rect 29088 19198 29126 19254
rect 29182 19198 29220 19254
rect 29276 19198 29304 19254
rect 29012 19182 29304 19198
rect 29884 20104 30176 20120
rect 29884 19946 29898 20104
rect 30160 19946 30176 20104
rect 29884 19442 30176 19946
rect 29884 19386 29904 19442
rect 29960 19386 29998 19442
rect 30054 19386 30092 19442
rect 30148 19386 30176 19442
rect 29884 19348 30176 19386
rect 29884 19292 29904 19348
rect 29960 19292 29998 19348
rect 30054 19292 30092 19348
rect 30148 19292 30176 19348
rect 29884 19254 30176 19292
rect 29884 19198 29904 19254
rect 29960 19198 29998 19254
rect 30054 19198 30092 19254
rect 30148 19198 30176 19254
rect 29884 19182 30176 19198
rect 30584 19442 30876 20166
rect 30584 19386 30604 19442
rect 30660 19386 30698 19442
rect 30754 19386 30792 19442
rect 30848 19386 30876 19442
rect 30584 19348 30876 19386
rect 30584 19292 30604 19348
rect 30660 19292 30698 19348
rect 30754 19292 30792 19348
rect 30848 19292 30876 19348
rect 30584 19254 30876 19292
rect 30584 19198 30604 19254
rect 30660 19198 30698 19254
rect 30754 19198 30792 19254
rect 30848 19198 30876 19254
rect 30584 19182 30876 19198
rect 33012 20104 33304 20120
rect 33012 19946 33026 20104
rect 33288 19946 33304 20104
rect 33012 19442 33304 19946
rect 33012 19386 33032 19442
rect 33088 19386 33126 19442
rect 33182 19386 33220 19442
rect 33276 19386 33304 19442
rect 33012 19348 33304 19386
rect 33012 19292 33032 19348
rect 33088 19292 33126 19348
rect 33182 19292 33220 19348
rect 33276 19292 33304 19348
rect 33012 19254 33304 19292
rect 33012 19198 33032 19254
rect 33088 19198 33126 19254
rect 33182 19198 33220 19254
rect 33276 19198 33304 19254
rect 33012 19182 33304 19198
rect 33884 20104 34176 20120
rect 33884 19946 33898 20104
rect 34160 19946 34176 20104
rect 33884 19442 34176 19946
rect 33884 19386 33904 19442
rect 33960 19386 33998 19442
rect 34054 19386 34092 19442
rect 34148 19386 34176 19442
rect 33884 19348 34176 19386
rect 33884 19292 33904 19348
rect 33960 19292 33998 19348
rect 34054 19292 34092 19348
rect 34148 19292 34176 19348
rect 33884 19254 34176 19292
rect 33884 19198 33904 19254
rect 33960 19198 33998 19254
rect 34054 19198 34092 19254
rect 34148 19198 34176 19254
rect 33884 19182 34176 19198
rect 34584 19442 34876 20166
rect 34584 19386 34604 19442
rect 34660 19386 34698 19442
rect 34754 19386 34792 19442
rect 34848 19386 34876 19442
rect 34584 19348 34876 19386
rect 34584 19292 34604 19348
rect 34660 19292 34698 19348
rect 34754 19292 34792 19348
rect 34848 19292 34876 19348
rect 34584 19254 34876 19292
rect 34584 19198 34604 19254
rect 34660 19198 34698 19254
rect 34754 19198 34792 19254
rect 34848 19198 34876 19254
rect 34584 19182 34876 19198
rect 37444 19212 37602 19276
rect 37444 19160 37451 19212
rect 37503 19160 37542 19212
rect 37594 19160 37602 19212
rect 37444 19110 37602 19160
rect 37444 19058 37451 19110
rect 37503 19058 37542 19110
rect 37594 19058 37602 19110
rect 37444 19007 37602 19058
rect 37444 18955 37452 19007
rect 37504 18955 37543 19007
rect 37595 18955 37602 19007
rect 37444 18914 37602 18955
rect 37444 18862 37452 18914
rect 37504 18862 37543 18914
rect 37595 18862 37602 18914
rect 37444 18816 37602 18862
rect 41602 19250 42660 19276
rect 41602 18838 42422 19250
rect 42634 18838 42660 19250
rect 41602 18814 42660 18838
rect 1046 18357 1460 18383
rect 1046 18356 1169 18357
rect 1046 18298 1074 18356
rect 1130 18299 1169 18356
rect 1225 18356 1460 18357
rect 1225 18299 1278 18356
rect 1130 18298 1278 18299
rect 1334 18298 1373 18356
rect 1429 18298 1460 18356
rect 1046 18273 1460 18298
rect 1046 18147 1460 18173
rect 1046 18146 1169 18147
rect 1046 18088 1074 18146
rect 1130 18089 1169 18146
rect 1225 18146 1460 18147
rect 1225 18089 1278 18146
rect 1130 18088 1278 18089
rect 1334 18088 1373 18146
rect 1429 18088 1460 18146
rect 1046 18063 1460 18088
rect 36064 18148 36478 18174
rect 36064 18147 36187 18148
rect 36064 18089 36092 18147
rect 36148 18090 36187 18147
rect 36243 18147 36478 18148
rect 36243 18090 36296 18147
rect 36148 18089 36296 18090
rect 36352 18089 36391 18147
rect 36447 18089 36478 18147
rect 36064 18064 36478 18089
rect 37444 17452 37602 17516
rect 37444 17400 37451 17452
rect 37503 17400 37542 17452
rect 37594 17400 37602 17452
rect 37444 17350 37602 17400
rect 37444 17298 37451 17350
rect 37503 17298 37542 17350
rect 37594 17298 37602 17350
rect 37444 17247 37602 17298
rect 37444 17195 37452 17247
rect 37504 17195 37543 17247
rect 37595 17195 37602 17247
rect 1046 17144 1460 17170
rect 1046 17143 1169 17144
rect 1046 17085 1074 17143
rect 1130 17086 1169 17143
rect 1225 17143 1460 17144
rect 1225 17086 1278 17143
rect 1130 17085 1278 17086
rect 1334 17085 1373 17143
rect 1429 17085 1460 17143
rect 1046 17060 1460 17085
rect 36064 17144 36478 17170
rect 36064 17143 36187 17144
rect 36064 17085 36092 17143
rect 36148 17086 36187 17143
rect 36243 17143 36478 17144
rect 36243 17086 36296 17143
rect 36148 17085 36296 17086
rect 36352 17085 36391 17143
rect 36447 17085 36478 17143
rect 36064 17060 36478 17085
rect 37444 17154 37602 17195
rect 37444 17102 37452 17154
rect 37504 17102 37543 17154
rect 37595 17102 37602 17154
rect 37444 17056 37602 17102
rect 41602 17492 42660 17518
rect 41602 17080 42422 17492
rect 42634 17080 42660 17492
rect 41602 17056 42660 17080
rect 1046 16139 1460 16165
rect 1046 16138 1169 16139
rect 1046 16080 1074 16138
rect 1130 16081 1169 16138
rect 1225 16138 1460 16139
rect 1225 16081 1278 16138
rect 1130 16080 1278 16081
rect 1334 16080 1373 16138
rect 1429 16080 1460 16138
rect 1046 16055 1460 16080
rect 36064 16140 36478 16166
rect 36064 16139 36187 16140
rect 36064 16081 36092 16139
rect 36148 16082 36187 16139
rect 36243 16139 36478 16140
rect 36243 16082 36296 16139
rect 36148 16081 36296 16082
rect 36352 16081 36391 16139
rect 36447 16081 36478 16139
rect 36064 16056 36478 16081
rect 37444 15212 37602 15276
rect 1046 15136 1460 15162
rect 1046 15135 1169 15136
rect 1046 15077 1074 15135
rect 1130 15078 1169 15135
rect 1225 15135 1460 15136
rect 1225 15078 1278 15135
rect 1130 15077 1278 15078
rect 1334 15077 1373 15135
rect 1429 15077 1460 15135
rect 1046 15052 1460 15077
rect 36064 15136 36478 15162
rect 36064 15135 36187 15136
rect 36064 15077 36092 15135
rect 36148 15078 36187 15135
rect 36243 15135 36478 15136
rect 36243 15078 36296 15135
rect 36148 15077 36296 15078
rect 36352 15077 36391 15135
rect 36447 15077 36478 15135
rect 36064 15052 36478 15077
rect 37444 15160 37451 15212
rect 37503 15160 37542 15212
rect 37594 15160 37602 15212
rect 37444 15110 37602 15160
rect 37444 15058 37451 15110
rect 37503 15058 37542 15110
rect 37594 15058 37602 15110
rect 37444 15007 37602 15058
rect 37444 14955 37452 15007
rect 37504 14955 37543 15007
rect 37595 14955 37602 15007
rect 37444 14914 37602 14955
rect 37444 14862 37452 14914
rect 37504 14862 37543 14914
rect 37595 14862 37602 14914
rect 37444 14816 37602 14862
rect 41602 15250 42660 15276
rect 41602 14838 42422 15250
rect 42634 14838 42660 15250
rect 41602 14814 42660 14838
rect 1046 14132 1460 14158
rect 1046 14131 1169 14132
rect 1046 14073 1074 14131
rect 1130 14074 1169 14131
rect 1225 14131 1460 14132
rect 1225 14074 1278 14131
rect 1130 14073 1278 14074
rect 1334 14073 1373 14131
rect 1429 14073 1460 14131
rect 1046 14048 1460 14073
rect 36064 14132 36478 14158
rect 36064 14131 36187 14132
rect 36064 14073 36092 14131
rect 36148 14074 36187 14131
rect 36243 14131 36478 14132
rect 36243 14074 36296 14131
rect 36148 14073 36296 14074
rect 36352 14073 36391 14131
rect 36447 14073 36478 14131
rect 36064 14048 36478 14073
rect 37444 13452 37602 13516
rect 37444 13400 37451 13452
rect 37503 13400 37542 13452
rect 37594 13400 37602 13452
rect 37444 13350 37602 13400
rect 37444 13298 37451 13350
rect 37503 13298 37542 13350
rect 37594 13298 37602 13350
rect 37444 13247 37602 13298
rect 37444 13195 37452 13247
rect 37504 13195 37543 13247
rect 37595 13195 37602 13247
rect 37444 13154 37602 13195
rect 1046 13128 1460 13154
rect 1046 13127 1169 13128
rect 1046 13069 1074 13127
rect 1130 13070 1169 13127
rect 1225 13127 1460 13128
rect 1225 13070 1278 13127
rect 1130 13069 1278 13070
rect 1334 13069 1373 13127
rect 1429 13069 1460 13127
rect 1046 13044 1460 13069
rect 36064 13128 36478 13154
rect 36064 13127 36187 13128
rect 36064 13069 36092 13127
rect 36148 13070 36187 13127
rect 36243 13127 36478 13128
rect 36243 13070 36296 13127
rect 36148 13069 36296 13070
rect 36352 13069 36391 13127
rect 36447 13069 36478 13127
rect 36064 13044 36478 13069
rect 37444 13102 37452 13154
rect 37504 13102 37543 13154
rect 37595 13102 37602 13154
rect 37444 13056 37602 13102
rect 41602 13492 42660 13518
rect 41602 13080 42422 13492
rect 42634 13080 42660 13492
rect 41602 13056 42660 13080
rect 1046 12124 1460 12150
rect 1046 12123 1169 12124
rect 1046 12065 1074 12123
rect 1130 12066 1169 12123
rect 1225 12123 1460 12124
rect 1225 12066 1278 12123
rect 1130 12065 1278 12066
rect 1334 12065 1373 12123
rect 1429 12065 1460 12123
rect 1046 12040 1460 12065
rect 36064 12124 36478 12150
rect 36064 12123 36187 12124
rect 36064 12065 36092 12123
rect 36148 12066 36187 12123
rect 36243 12123 36478 12124
rect 36243 12066 36296 12123
rect 36148 12065 36296 12066
rect 36352 12065 36391 12123
rect 36447 12065 36478 12123
rect 36064 12040 36478 12065
rect 37444 11212 37602 11276
rect 37444 11160 37451 11212
rect 37503 11160 37542 11212
rect 37594 11160 37602 11212
rect 1046 11120 1460 11146
rect 1046 11119 1169 11120
rect 1046 11061 1074 11119
rect 1130 11062 1169 11119
rect 1225 11119 1460 11120
rect 1225 11062 1278 11119
rect 1130 11061 1278 11062
rect 1334 11061 1373 11119
rect 1429 11061 1460 11119
rect 1046 11036 1460 11061
rect 36064 11120 36478 11146
rect 36064 11119 36187 11120
rect 36064 11061 36092 11119
rect 36148 11062 36187 11119
rect 36243 11119 36478 11120
rect 36243 11062 36296 11119
rect 36148 11061 36296 11062
rect 36352 11061 36391 11119
rect 36447 11061 36478 11119
rect 36064 11036 36478 11061
rect 37444 11110 37602 11160
rect 37444 11058 37451 11110
rect 37503 11058 37542 11110
rect 37594 11058 37602 11110
rect 37444 11007 37602 11058
rect 37444 10955 37452 11007
rect 37504 10955 37543 11007
rect 37595 10955 37602 11007
rect 37444 10914 37602 10955
rect 37444 10862 37452 10914
rect 37504 10862 37543 10914
rect 37595 10862 37602 10914
rect 37444 10816 37602 10862
rect 41602 11250 42660 11276
rect 41602 10838 42422 11250
rect 42634 10838 42660 11250
rect 41602 10814 42660 10838
rect 1046 10116 1460 10142
rect 1046 10115 1169 10116
rect 1046 10057 1074 10115
rect 1130 10058 1169 10115
rect 1225 10115 1460 10116
rect 1225 10058 1278 10115
rect 1130 10057 1278 10058
rect 1334 10057 1373 10115
rect 1429 10057 1460 10115
rect 1046 10032 1460 10057
rect 36064 10116 36478 10142
rect 36064 10115 36187 10116
rect 36064 10057 36092 10115
rect 36148 10058 36187 10115
rect 36243 10115 36478 10116
rect 36243 10058 36296 10115
rect 36148 10057 36296 10058
rect 36352 10057 36391 10115
rect 36447 10057 36478 10115
rect 36064 10032 36478 10057
rect 37444 9452 37602 9516
rect 37444 9400 37451 9452
rect 37503 9400 37542 9452
rect 37594 9400 37602 9452
rect 37444 9350 37602 9400
rect 37444 9298 37451 9350
rect 37503 9298 37542 9350
rect 37594 9298 37602 9350
rect 37444 9247 37602 9298
rect 37444 9195 37452 9247
rect 37504 9195 37543 9247
rect 37595 9195 37602 9247
rect 37444 9154 37602 9195
rect 1046 9112 1460 9138
rect 1046 9111 1169 9112
rect 1046 9053 1074 9111
rect 1130 9054 1169 9111
rect 1225 9111 1460 9112
rect 1225 9054 1278 9111
rect 1130 9053 1278 9054
rect 1334 9053 1373 9111
rect 1429 9053 1460 9111
rect 1046 9028 1460 9053
rect 36064 9112 36478 9138
rect 36064 9111 36187 9112
rect 36064 9053 36092 9111
rect 36148 9054 36187 9111
rect 36243 9111 36478 9112
rect 36243 9054 36296 9111
rect 36148 9053 36296 9054
rect 36352 9053 36391 9111
rect 36447 9053 36478 9111
rect 37444 9102 37452 9154
rect 37504 9102 37543 9154
rect 37595 9102 37602 9154
rect 37444 9056 37602 9102
rect 41602 9492 42660 9518
rect 41602 9080 42422 9492
rect 42634 9080 42660 9492
rect 41602 9056 42660 9080
rect 36064 9028 36478 9053
rect 1046 8108 1460 8134
rect 1046 8107 1169 8108
rect 1046 8049 1074 8107
rect 1130 8050 1169 8107
rect 1225 8107 1460 8108
rect 1225 8050 1278 8107
rect 1130 8049 1278 8050
rect 1334 8049 1373 8107
rect 1429 8049 1460 8107
rect 1046 8024 1460 8049
rect 36064 8108 36478 8134
rect 36064 8107 36187 8108
rect 36064 8049 36092 8107
rect 36148 8050 36187 8107
rect 36243 8107 36478 8108
rect 36243 8050 36296 8107
rect 36148 8049 36296 8050
rect 36352 8049 36391 8107
rect 36447 8049 36478 8107
rect 36064 8024 36478 8049
rect 37444 7212 37602 7276
rect 37444 7160 37451 7212
rect 37503 7160 37542 7212
rect 37594 7160 37602 7212
rect 1046 7104 1460 7130
rect 1046 7103 1169 7104
rect 1046 7045 1074 7103
rect 1130 7046 1169 7103
rect 1225 7103 1460 7104
rect 1225 7046 1278 7103
rect 1130 7045 1278 7046
rect 1334 7045 1373 7103
rect 1429 7045 1460 7103
rect 1046 7020 1460 7045
rect 36064 7104 36478 7130
rect 36064 7103 36187 7104
rect 36064 7045 36092 7103
rect 36148 7046 36187 7103
rect 36243 7103 36478 7104
rect 36243 7046 36296 7103
rect 36148 7045 36296 7046
rect 36352 7045 36391 7103
rect 36447 7045 36478 7103
rect 36064 7020 36478 7045
rect 37444 7110 37602 7160
rect 37444 7058 37451 7110
rect 37503 7058 37542 7110
rect 37594 7058 37602 7110
rect 37444 7007 37602 7058
rect 37444 6955 37452 7007
rect 37504 6955 37543 7007
rect 37595 6955 37602 7007
rect 37444 6914 37602 6955
rect 37444 6862 37452 6914
rect 37504 6862 37543 6914
rect 37595 6862 37602 6914
rect 37444 6816 37602 6862
rect 41602 7250 42660 7276
rect 41602 6838 42422 7250
rect 42634 6838 42660 7250
rect 41602 6814 42660 6838
rect 1046 6100 1460 6126
rect 1046 6099 1169 6100
rect 1046 6041 1074 6099
rect 1130 6042 1169 6099
rect 1225 6099 1460 6100
rect 1225 6042 1278 6099
rect 1130 6041 1278 6042
rect 1334 6041 1373 6099
rect 1429 6041 1460 6099
rect 1046 6016 1460 6041
rect 36064 6100 36478 6126
rect 36064 6099 36187 6100
rect 36064 6041 36092 6099
rect 36148 6042 36187 6099
rect 36243 6099 36478 6100
rect 36243 6042 36296 6099
rect 36148 6041 36296 6042
rect 36352 6041 36391 6099
rect 36447 6041 36478 6099
rect 36064 6016 36478 6041
rect 37444 5452 37602 5516
rect 37444 5400 37451 5452
rect 37503 5400 37542 5452
rect 37594 5400 37602 5452
rect 37444 5350 37602 5400
rect 37444 5298 37451 5350
rect 37503 5298 37542 5350
rect 37594 5298 37602 5350
rect 37444 5247 37602 5298
rect 37444 5195 37452 5247
rect 37504 5195 37543 5247
rect 37595 5195 37602 5247
rect 37444 5154 37602 5195
rect 1046 5096 1460 5122
rect 1046 5095 1169 5096
rect 1046 5037 1074 5095
rect 1130 5038 1169 5095
rect 1225 5095 1460 5096
rect 1225 5038 1278 5095
rect 1130 5037 1278 5038
rect 1334 5037 1373 5095
rect 1429 5037 1460 5095
rect 1046 5012 1460 5037
rect 36064 5096 36478 5122
rect 36064 5095 36187 5096
rect 36064 5037 36092 5095
rect 36148 5038 36187 5095
rect 36243 5095 36478 5096
rect 36243 5038 36296 5095
rect 36148 5037 36296 5038
rect 36352 5037 36391 5095
rect 36447 5037 36478 5095
rect 37444 5102 37452 5154
rect 37504 5102 37543 5154
rect 37595 5102 37602 5154
rect 37444 5056 37602 5102
rect 41602 5492 42660 5518
rect 41602 5080 42422 5492
rect 42634 5080 42660 5492
rect 41602 5056 42660 5080
rect 36064 5012 36478 5037
rect 1046 4092 1460 4118
rect 1046 4091 1169 4092
rect 1046 4033 1074 4091
rect 1130 4034 1169 4091
rect 1225 4091 1460 4092
rect 1225 4034 1278 4091
rect 1130 4033 1278 4034
rect 1334 4033 1373 4091
rect 1429 4033 1460 4091
rect 1046 4008 1460 4033
rect 36064 4092 36478 4118
rect 36064 4091 36187 4092
rect 36064 4033 36092 4091
rect 36148 4034 36187 4091
rect 36243 4091 36478 4092
rect 36243 4034 36296 4091
rect 36148 4033 36296 4034
rect 36352 4033 36391 4091
rect 36447 4033 36478 4091
rect 36064 4008 36478 4033
rect 37444 3222 37602 3276
rect 37444 3170 37451 3222
rect 37503 3170 37542 3222
rect 37594 3170 37602 3222
rect 37444 3120 37602 3170
rect 1046 3086 1460 3112
rect 1046 3085 1169 3086
rect 1046 3027 1074 3085
rect 1130 3028 1169 3085
rect 1225 3085 1460 3086
rect 1225 3028 1278 3085
rect 1130 3027 1278 3028
rect 1334 3027 1373 3085
rect 1429 3027 1460 3085
rect 1046 3002 1460 3027
rect 36064 3088 36478 3114
rect 36064 3087 36187 3088
rect 36064 3029 36092 3087
rect 36148 3030 36187 3087
rect 36243 3087 36478 3088
rect 36243 3030 36296 3087
rect 36148 3029 36296 3030
rect 36352 3029 36391 3087
rect 36447 3029 36478 3087
rect 36064 3004 36478 3029
rect 37444 3068 37451 3120
rect 37503 3068 37542 3120
rect 37594 3068 37602 3120
rect 37444 3017 37602 3068
rect 37444 2965 37452 3017
rect 37504 2965 37543 3017
rect 37595 2965 37602 3017
rect 37444 2924 37602 2965
rect 37444 2872 37452 2924
rect 37504 2872 37543 2924
rect 37595 2872 37602 2924
rect 37444 2816 37602 2872
rect 41602 3250 42660 3276
rect 41602 2838 42422 3250
rect 42634 2838 42660 3250
rect 41602 2814 42660 2838
rect 1046 2083 1460 2109
rect 1046 2082 1169 2083
rect 1046 2024 1074 2082
rect 1130 2025 1169 2082
rect 1225 2082 1460 2083
rect 1225 2025 1278 2082
rect 1130 2024 1278 2025
rect 1334 2024 1373 2082
rect 1429 2024 1460 2082
rect 1046 1999 1460 2024
rect 36064 2084 36478 2110
rect 36064 2083 36187 2084
rect 36064 2025 36092 2083
rect 36148 2026 36187 2083
rect 36243 2083 36478 2084
rect 36243 2026 36296 2083
rect 36148 2025 36296 2026
rect 36352 2025 36391 2083
rect 36447 2025 36478 2083
rect 36064 2000 36478 2025
rect 1046 1428 1460 1454
rect 1046 1427 1169 1428
rect 1046 1369 1074 1427
rect 1130 1370 1169 1427
rect 1225 1427 1460 1428
rect 1225 1370 1278 1427
rect 1130 1369 1278 1370
rect 1334 1369 1373 1427
rect 1429 1369 1460 1427
rect 1046 1318 1460 1369
rect 1046 1317 1169 1318
rect 1046 1259 1074 1317
rect 1130 1260 1169 1317
rect 1225 1317 1460 1318
rect 1225 1260 1278 1317
rect 1130 1259 1278 1260
rect 1334 1259 1373 1317
rect 1429 1259 1460 1317
rect 1046 1234 1460 1259
rect 37444 1452 37602 1516
rect 37444 1400 37451 1452
rect 37503 1400 37542 1452
rect 37594 1400 37602 1452
rect 37444 1350 37602 1400
rect 37444 1298 37451 1350
rect 37503 1298 37542 1350
rect 37594 1298 37602 1350
rect 37444 1247 37602 1298
rect 37444 1195 37452 1247
rect 37504 1195 37543 1247
rect 37595 1195 37602 1247
rect 37444 1154 37602 1195
rect 1046 1079 1460 1105
rect 1046 1078 1169 1079
rect 1046 1020 1074 1078
rect 1130 1021 1169 1078
rect 1225 1078 1460 1079
rect 1225 1021 1278 1078
rect 1130 1020 1278 1021
rect 1334 1020 1373 1078
rect 1429 1020 1460 1078
rect 1046 995 1460 1020
rect 36064 1080 36478 1106
rect 36064 1079 36187 1080
rect 36064 1021 36092 1079
rect 36148 1022 36187 1079
rect 36243 1079 36478 1080
rect 36243 1022 36296 1079
rect 36148 1021 36296 1022
rect 36352 1021 36391 1079
rect 36447 1021 36478 1079
rect 37444 1102 37452 1154
rect 37504 1102 37543 1154
rect 37595 1102 37602 1154
rect 37444 1056 37602 1102
rect 41602 1492 42660 1518
rect 41602 1080 42422 1492
rect 42634 1080 42660 1492
rect 41602 1056 42660 1080
rect 36064 996 36478 1021
rect 2554 893 2670 914
rect 2554 859 2565 893
rect 2662 859 2670 893
rect 2554 847 2670 859
rect 3558 891 3674 914
rect 3558 857 3569 891
rect 3666 857 3674 891
rect 3558 846 3674 857
rect 4194 893 4310 914
rect 4194 859 4205 893
rect 4302 859 4310 893
rect 4194 847 4310 859
rect 4562 892 4678 914
rect 4562 858 4573 892
rect 4670 858 4678 892
rect 4230 846 4264 847
rect 4562 846 4678 858
rect 5566 892 5682 914
rect 5566 858 5577 892
rect 5674 858 5682 892
rect 5566 846 5682 858
rect 6570 892 6686 914
rect 6570 858 6581 892
rect 6678 858 6686 892
rect 6570 846 6686 858
rect 7574 892 7690 914
rect 7574 858 7585 892
rect 7682 858 7690 892
rect 7574 846 7690 858
rect 8578 892 8694 914
rect 8578 858 8589 892
rect 8686 858 8694 892
rect 8578 846 8694 858
rect 9582 892 9698 914
rect 9582 858 9593 892
rect 9690 858 9698 892
rect 9582 846 9698 858
rect 10586 892 10702 914
rect 10586 858 10597 892
rect 10694 858 10702 892
rect 10586 846 10702 858
rect 11590 892 11706 914
rect 11590 858 11601 892
rect 11698 858 11706 892
rect 11590 846 11706 858
rect 12594 892 12710 914
rect 12594 858 12605 892
rect 12702 858 12710 892
rect 12594 846 12710 858
rect 13598 892 13714 914
rect 13598 858 13609 892
rect 13706 858 13714 892
rect 13598 846 13714 858
rect 14602 892 14718 914
rect 14602 858 14613 892
rect 14710 858 14718 892
rect 14602 846 14718 858
rect 15606 892 15722 914
rect 15606 858 15617 892
rect 15714 858 15722 892
rect 15606 846 15722 858
rect 16610 892 16726 914
rect 16610 858 16621 892
rect 16718 858 16726 892
rect 16610 846 16726 858
rect 17614 892 17730 914
rect 17614 858 17625 892
rect 17722 858 17730 892
rect 17614 846 17730 858
rect 18244 893 18360 914
rect 18244 859 18255 893
rect 18352 859 18360 893
rect 18244 847 18360 859
rect 18618 892 18734 914
rect 18618 858 18629 892
rect 18726 858 18734 892
rect 18286 846 18320 847
rect 18618 846 18734 858
rect 19250 893 19366 914
rect 19250 859 19261 893
rect 19358 859 19366 893
rect 19250 847 19366 859
rect 19622 892 19738 914
rect 19622 858 19633 892
rect 19730 858 19738 892
rect 19290 846 19324 847
rect 19622 846 19738 858
rect 20246 893 20362 914
rect 20246 859 20257 893
rect 20354 859 20362 893
rect 20246 847 20362 859
rect 20626 892 20742 914
rect 20626 858 20637 892
rect 20734 858 20742 892
rect 20294 846 20328 847
rect 20626 846 20742 858
rect 21630 892 21746 914
rect 21630 858 21641 892
rect 21738 858 21746 892
rect 21630 846 21746 858
rect 22634 892 22750 914
rect 22634 858 22645 892
rect 22742 858 22750 892
rect 22634 846 22750 858
rect 23638 892 23754 914
rect 23638 858 23649 892
rect 23746 858 23754 892
rect 23638 846 23754 858
rect 24642 892 24758 914
rect 24642 858 24653 892
rect 24750 858 24758 892
rect 24642 846 24758 858
rect 25646 892 25762 914
rect 25646 858 25657 892
rect 25754 858 25762 892
rect 25646 846 25762 858
rect 26650 892 26766 914
rect 26650 858 26661 892
rect 26758 858 26766 892
rect 26650 846 26766 858
rect 27654 892 27770 914
rect 27654 858 27665 892
rect 27762 858 27770 892
rect 27654 846 27770 858
rect 28658 892 28774 914
rect 28658 858 28669 892
rect 28766 858 28774 892
rect 28658 846 28774 858
rect 29662 892 29778 914
rect 29662 858 29673 892
rect 29770 858 29778 892
rect 29662 846 29778 858
rect 30666 893 30782 914
rect 30666 858 30677 893
rect 30774 858 30782 893
rect 30666 846 30782 858
rect 31670 893 31786 914
rect 31670 858 31681 893
rect 31778 858 31786 893
rect 31670 846 31786 858
rect 32674 893 32790 914
rect 32674 858 32685 893
rect 32782 858 32790 893
rect 32674 846 32790 858
rect 33600 893 33716 914
rect 33600 858 33611 893
rect 33708 858 33716 893
rect 33600 846 33716 858
rect 34682 893 34798 914
rect 34682 858 34693 893
rect 34790 858 34798 893
rect 34682 846 34798 858
rect 35686 493 35720 914
rect 35686 487 35728 493
rect 35686 453 35690 487
rect 35724 453 35728 487
rect 35686 447 35728 453
<< viali >>
rect 42422 22838 42634 23250
rect 42422 21080 42634 21492
rect 1898 19946 2160 20104
rect 1904 19386 1960 19442
rect 1998 19386 2054 19442
rect 2092 19386 2148 19442
rect 1904 19292 1960 19348
rect 1998 19292 2054 19348
rect 2092 19292 2148 19348
rect 1904 19198 1960 19254
rect 1998 19198 2054 19254
rect 2092 19198 2148 19254
rect 2604 19386 2660 19442
rect 2698 19386 2754 19442
rect 2792 19386 2848 19442
rect 2604 19292 2660 19348
rect 2698 19292 2754 19348
rect 2792 19292 2848 19348
rect 2604 19198 2660 19254
rect 2698 19198 2754 19254
rect 2792 19198 2848 19254
rect 5026 19946 5288 20104
rect 5032 19386 5088 19442
rect 5126 19386 5182 19442
rect 5220 19386 5276 19442
rect 5032 19292 5088 19348
rect 5126 19292 5182 19348
rect 5220 19292 5276 19348
rect 5032 19198 5088 19254
rect 5126 19198 5182 19254
rect 5220 19198 5276 19254
rect 5898 19946 6160 20104
rect 5904 19386 5960 19442
rect 5998 19386 6054 19442
rect 6092 19386 6148 19442
rect 5904 19292 5960 19348
rect 5998 19292 6054 19348
rect 6092 19292 6148 19348
rect 5904 19198 5960 19254
rect 5998 19198 6054 19254
rect 6092 19198 6148 19254
rect 6604 19386 6660 19442
rect 6698 19386 6754 19442
rect 6792 19386 6848 19442
rect 6604 19292 6660 19348
rect 6698 19292 6754 19348
rect 6792 19292 6848 19348
rect 6604 19198 6660 19254
rect 6698 19198 6754 19254
rect 6792 19198 6848 19254
rect 9026 19946 9288 20104
rect 9032 19386 9088 19442
rect 9126 19386 9182 19442
rect 9220 19386 9276 19442
rect 9032 19292 9088 19348
rect 9126 19292 9182 19348
rect 9220 19292 9276 19348
rect 9032 19198 9088 19254
rect 9126 19198 9182 19254
rect 9220 19198 9276 19254
rect 9898 19946 10160 20104
rect 9904 19386 9960 19442
rect 9998 19386 10054 19442
rect 10092 19386 10148 19442
rect 9904 19292 9960 19348
rect 9998 19292 10054 19348
rect 10092 19292 10148 19348
rect 9904 19198 9960 19254
rect 9998 19198 10054 19254
rect 10092 19198 10148 19254
rect 10604 19386 10660 19442
rect 10698 19386 10754 19442
rect 10792 19386 10848 19442
rect 10604 19292 10660 19348
rect 10698 19292 10754 19348
rect 10792 19292 10848 19348
rect 10604 19198 10660 19254
rect 10698 19198 10754 19254
rect 10792 19198 10848 19254
rect 13026 19946 13288 20104
rect 13032 19386 13088 19442
rect 13126 19386 13182 19442
rect 13220 19386 13276 19442
rect 13032 19292 13088 19348
rect 13126 19292 13182 19348
rect 13220 19292 13276 19348
rect 13032 19198 13088 19254
rect 13126 19198 13182 19254
rect 13220 19198 13276 19254
rect 13898 19946 14160 20104
rect 13904 19386 13960 19442
rect 13998 19386 14054 19442
rect 14092 19386 14148 19442
rect 13904 19292 13960 19348
rect 13998 19292 14054 19348
rect 14092 19292 14148 19348
rect 13904 19198 13960 19254
rect 13998 19198 14054 19254
rect 14092 19198 14148 19254
rect 14604 19386 14660 19442
rect 14698 19386 14754 19442
rect 14792 19386 14848 19442
rect 14604 19292 14660 19348
rect 14698 19292 14754 19348
rect 14792 19292 14848 19348
rect 14604 19198 14660 19254
rect 14698 19198 14754 19254
rect 14792 19198 14848 19254
rect 17026 19946 17288 20104
rect 17032 19386 17088 19442
rect 17126 19386 17182 19442
rect 17220 19386 17276 19442
rect 17032 19292 17088 19348
rect 17126 19292 17182 19348
rect 17220 19292 17276 19348
rect 17032 19198 17088 19254
rect 17126 19198 17182 19254
rect 17220 19198 17276 19254
rect 17898 19946 18160 20104
rect 17904 19386 17960 19442
rect 17998 19386 18054 19442
rect 18092 19386 18148 19442
rect 17904 19292 17960 19348
rect 17998 19292 18054 19348
rect 18092 19292 18148 19348
rect 17904 19198 17960 19254
rect 17998 19198 18054 19254
rect 18092 19198 18148 19254
rect 18604 19386 18660 19442
rect 18698 19386 18754 19442
rect 18792 19386 18848 19442
rect 18604 19292 18660 19348
rect 18698 19292 18754 19348
rect 18792 19292 18848 19348
rect 18604 19198 18660 19254
rect 18698 19198 18754 19254
rect 18792 19198 18848 19254
rect 21026 19946 21288 20104
rect 21032 19386 21088 19442
rect 21126 19386 21182 19442
rect 21220 19386 21276 19442
rect 21032 19292 21088 19348
rect 21126 19292 21182 19348
rect 21220 19292 21276 19348
rect 21032 19198 21088 19254
rect 21126 19198 21182 19254
rect 21220 19198 21276 19254
rect 21898 19946 22160 20104
rect 21904 19386 21960 19442
rect 21998 19386 22054 19442
rect 22092 19386 22148 19442
rect 21904 19292 21960 19348
rect 21998 19292 22054 19348
rect 22092 19292 22148 19348
rect 21904 19198 21960 19254
rect 21998 19198 22054 19254
rect 22092 19198 22148 19254
rect 22604 19386 22660 19442
rect 22698 19386 22754 19442
rect 22792 19386 22848 19442
rect 22604 19292 22660 19348
rect 22698 19292 22754 19348
rect 22792 19292 22848 19348
rect 22604 19198 22660 19254
rect 22698 19198 22754 19254
rect 22792 19198 22848 19254
rect 25026 19946 25288 20104
rect 25032 19386 25088 19442
rect 25126 19386 25182 19442
rect 25220 19386 25276 19442
rect 25032 19292 25088 19348
rect 25126 19292 25182 19348
rect 25220 19292 25276 19348
rect 25032 19198 25088 19254
rect 25126 19198 25182 19254
rect 25220 19198 25276 19254
rect 25898 19946 26160 20104
rect 25904 19386 25960 19442
rect 25998 19386 26054 19442
rect 26092 19386 26148 19442
rect 25904 19292 25960 19348
rect 25998 19292 26054 19348
rect 26092 19292 26148 19348
rect 25904 19198 25960 19254
rect 25998 19198 26054 19254
rect 26092 19198 26148 19254
rect 26604 19386 26660 19442
rect 26698 19386 26754 19442
rect 26792 19386 26848 19442
rect 26604 19292 26660 19348
rect 26698 19292 26754 19348
rect 26792 19292 26848 19348
rect 26604 19198 26660 19254
rect 26698 19198 26754 19254
rect 26792 19198 26848 19254
rect 29026 19946 29288 20104
rect 29032 19386 29088 19442
rect 29126 19386 29182 19442
rect 29220 19386 29276 19442
rect 29032 19292 29088 19348
rect 29126 19292 29182 19348
rect 29220 19292 29276 19348
rect 29032 19198 29088 19254
rect 29126 19198 29182 19254
rect 29220 19198 29276 19254
rect 29898 19946 30160 20104
rect 29904 19386 29960 19442
rect 29998 19386 30054 19442
rect 30092 19386 30148 19442
rect 29904 19292 29960 19348
rect 29998 19292 30054 19348
rect 30092 19292 30148 19348
rect 29904 19198 29960 19254
rect 29998 19198 30054 19254
rect 30092 19198 30148 19254
rect 30604 19386 30660 19442
rect 30698 19386 30754 19442
rect 30792 19386 30848 19442
rect 30604 19292 30660 19348
rect 30698 19292 30754 19348
rect 30792 19292 30848 19348
rect 30604 19198 30660 19254
rect 30698 19198 30754 19254
rect 30792 19198 30848 19254
rect 33026 19946 33288 20104
rect 33032 19386 33088 19442
rect 33126 19386 33182 19442
rect 33220 19386 33276 19442
rect 33032 19292 33088 19348
rect 33126 19292 33182 19348
rect 33220 19292 33276 19348
rect 33032 19198 33088 19254
rect 33126 19198 33182 19254
rect 33220 19198 33276 19254
rect 33898 19946 34160 20104
rect 33904 19386 33960 19442
rect 33998 19386 34054 19442
rect 34092 19386 34148 19442
rect 33904 19292 33960 19348
rect 33998 19292 34054 19348
rect 34092 19292 34148 19348
rect 33904 19198 33960 19254
rect 33998 19198 34054 19254
rect 34092 19198 34148 19254
rect 34604 19386 34660 19442
rect 34698 19386 34754 19442
rect 34792 19386 34848 19442
rect 34604 19292 34660 19348
rect 34698 19292 34754 19348
rect 34792 19292 34848 19348
rect 34604 19198 34660 19254
rect 34698 19198 34754 19254
rect 34792 19198 34848 19254
rect 37451 19160 37503 19212
rect 37542 19160 37594 19212
rect 37451 19058 37503 19110
rect 37542 19058 37594 19110
rect 37452 18955 37504 19007
rect 37543 18955 37595 19007
rect 37452 18862 37504 18914
rect 37543 18862 37595 18914
rect 42422 18838 42634 19250
rect 37451 17400 37503 17452
rect 37542 17400 37594 17452
rect 37451 17298 37503 17350
rect 37542 17298 37594 17350
rect 37452 17195 37504 17247
rect 37543 17195 37595 17247
rect 37452 17102 37504 17154
rect 37543 17102 37595 17154
rect 42422 17080 42634 17492
rect 37451 15160 37503 15212
rect 37542 15160 37594 15212
rect 37451 15058 37503 15110
rect 37542 15058 37594 15110
rect 37452 14955 37504 15007
rect 37543 14955 37595 15007
rect 37452 14862 37504 14914
rect 37543 14862 37595 14914
rect 42422 14838 42634 15250
rect 37451 13400 37503 13452
rect 37542 13400 37594 13452
rect 37451 13298 37503 13350
rect 37542 13298 37594 13350
rect 37452 13195 37504 13247
rect 37543 13195 37595 13247
rect 37452 13102 37504 13154
rect 37543 13102 37595 13154
rect 42422 13080 42634 13492
rect 37451 11160 37503 11212
rect 37542 11160 37594 11212
rect 37451 11058 37503 11110
rect 37542 11058 37594 11110
rect 37452 10955 37504 11007
rect 37543 10955 37595 11007
rect 37452 10862 37504 10914
rect 37543 10862 37595 10914
rect 42422 10838 42634 11250
rect 37451 9400 37503 9452
rect 37542 9400 37594 9452
rect 37451 9298 37503 9350
rect 37542 9298 37594 9350
rect 37452 9195 37504 9247
rect 37543 9195 37595 9247
rect 37452 9102 37504 9154
rect 37543 9102 37595 9154
rect 42422 9080 42634 9492
rect 37451 7160 37503 7212
rect 37542 7160 37594 7212
rect 37451 7058 37503 7110
rect 37542 7058 37594 7110
rect 37452 6955 37504 7007
rect 37543 6955 37595 7007
rect 37452 6862 37504 6914
rect 37543 6862 37595 6914
rect 42422 6838 42634 7250
rect 37451 5400 37503 5452
rect 37542 5400 37594 5452
rect 37451 5298 37503 5350
rect 37542 5298 37594 5350
rect 37452 5195 37504 5247
rect 37543 5195 37595 5247
rect 37452 5102 37504 5154
rect 37543 5102 37595 5154
rect 42422 5080 42634 5492
rect 37451 3170 37503 3222
rect 37542 3170 37594 3222
rect 37451 3068 37503 3120
rect 37542 3068 37594 3120
rect 37452 2965 37504 3017
rect 37543 2965 37595 3017
rect 37452 2872 37504 2924
rect 37543 2872 37595 2924
rect 42422 2838 42634 3250
rect 37451 1400 37503 1452
rect 37542 1400 37594 1452
rect 37451 1298 37503 1350
rect 37542 1298 37594 1350
rect 37452 1195 37504 1247
rect 37543 1195 37595 1247
rect 37452 1102 37504 1154
rect 37543 1102 37595 1154
rect 42422 1080 42634 1492
rect 2565 859 2662 893
rect 3569 857 3666 891
rect 4205 859 4302 893
rect 4573 858 4670 892
rect 5577 858 5674 892
rect 6581 858 6678 892
rect 7585 858 7682 892
rect 8589 858 8686 892
rect 9593 858 9690 892
rect 10597 858 10694 892
rect 11601 858 11698 892
rect 12605 858 12702 892
rect 13609 858 13706 892
rect 14613 858 14710 892
rect 15617 858 15714 892
rect 16621 858 16718 892
rect 17625 858 17722 892
rect 18255 859 18352 893
rect 18629 858 18726 892
rect 19261 859 19358 893
rect 19633 858 19730 892
rect 20257 859 20354 893
rect 20637 858 20734 892
rect 21641 858 21738 892
rect 22645 858 22742 892
rect 23649 858 23746 892
rect 24653 858 24750 892
rect 25657 858 25754 892
rect 26661 858 26758 892
rect 27665 858 27762 892
rect 28669 858 28766 892
rect 29673 858 29770 892
rect 30677 858 30774 893
rect 31681 858 31778 893
rect 32685 858 32782 893
rect 33611 858 33708 893
rect 34693 858 34790 893
rect 35690 453 35724 487
<< metal1 >>
rect 41602 23656 42660 23668
rect 41602 23494 42410 23656
rect 42648 23494 42660 23656
rect 41602 23484 42660 23494
rect 42396 23250 42660 23276
rect 42396 22838 42422 23250
rect 42634 22838 42660 23250
rect 42396 22814 42660 22838
rect 41602 22788 42164 22806
rect 41602 22638 41930 22788
rect 42142 22638 42164 22788
rect 41602 22624 42164 22638
rect 41602 22246 42164 22264
rect 41602 22096 41930 22246
rect 42142 22096 42164 22246
rect 41602 22082 42164 22096
rect 41602 21690 42164 21708
rect 41602 21540 41930 21690
rect 42142 21540 42164 21690
rect 41602 21526 42164 21540
rect 42396 21492 42660 21518
rect 42396 21080 42422 21492
rect 42634 21080 42660 21492
rect 42396 21056 42660 21080
rect 41602 20546 42660 20558
rect 41602 20384 42410 20546
rect 42648 20384 42660 20546
rect 41602 20374 42660 20384
rect 1884 20104 2176 20166
rect 1884 19946 1898 20104
rect 2160 19946 2176 20104
rect 1884 19934 2176 19946
rect 3420 19900 3790 20166
rect 5012 20104 5304 20166
rect 5012 19946 5026 20104
rect 5288 19946 5304 20104
rect 5012 19934 5304 19946
rect 5884 20104 6176 20166
rect 5884 19946 5898 20104
rect 6160 19946 6176 20104
rect 5884 19934 6176 19946
rect 7420 19900 7790 20166
rect 9012 20104 9304 20166
rect 9012 19946 9026 20104
rect 9288 19946 9304 20104
rect 9012 19934 9304 19946
rect 9884 20104 10176 20166
rect 9884 19946 9898 20104
rect 10160 19946 10176 20104
rect 9884 19934 10176 19946
rect 11420 19900 11790 20166
rect 13012 20104 13304 20166
rect 13012 19946 13026 20104
rect 13288 19946 13304 20104
rect 13012 19934 13304 19946
rect 13884 20104 14176 20166
rect 13884 19946 13898 20104
rect 14160 19946 14176 20104
rect 13884 19934 14176 19946
rect 15420 19900 15790 20166
rect 17012 20104 17304 20166
rect 17012 19946 17026 20104
rect 17288 19946 17304 20104
rect 17012 19934 17304 19946
rect 17884 20104 18176 20166
rect 17884 19946 17898 20104
rect 18160 19946 18176 20104
rect 17884 19934 18176 19946
rect 19420 19900 19790 20166
rect 21012 20104 21304 20166
rect 21012 19946 21026 20104
rect 21288 19946 21304 20104
rect 21012 19934 21304 19946
rect 21884 20104 22176 20166
rect 21884 19946 21898 20104
rect 22160 19946 22176 20104
rect 21884 19934 22176 19946
rect 23420 19900 23790 20166
rect 25012 20104 25304 20166
rect 25012 19946 25026 20104
rect 25288 19946 25304 20104
rect 25012 19934 25304 19946
rect 25884 20104 26176 20166
rect 25884 19946 25898 20104
rect 26160 19946 26176 20104
rect 25884 19934 26176 19946
rect 27420 19900 27790 20166
rect 29012 20104 29304 20166
rect 29012 19946 29026 20104
rect 29288 19946 29304 20104
rect 29012 19934 29304 19946
rect 29884 20104 30176 20166
rect 29884 19946 29898 20104
rect 30160 19946 30176 20104
rect 29884 19934 30176 19946
rect 31420 19900 31790 20166
rect 33012 20104 33304 20166
rect 33012 19946 33026 20104
rect 33288 19946 33304 20104
rect 33012 19934 33304 19946
rect 33884 20104 34176 20166
rect 33884 19946 33898 20104
rect 34160 19946 34176 20104
rect 35412 19974 35782 20166
rect 37012 20104 37304 20166
rect 37012 19980 37026 20104
rect 37288 19980 37304 20104
rect 37012 19968 37304 19980
rect 33884 19934 34176 19946
rect 0 19889 36954 19900
rect 0 19634 587 19889
rect 969 19885 36954 19889
rect 969 19882 36570 19885
rect 969 19638 3444 19882
rect 3770 19638 7444 19882
rect 7770 19638 11444 19882
rect 11770 19638 15444 19882
rect 15770 19638 19444 19882
rect 19770 19638 23444 19882
rect 23770 19638 27444 19882
rect 27770 19638 31444 19882
rect 31770 19847 36570 19882
rect 31770 19783 35426 19847
rect 35490 19783 35522 19847
rect 35586 19783 35618 19847
rect 35682 19783 35714 19847
rect 35778 19821 36570 19847
rect 36634 19821 36666 19885
rect 36730 19821 36762 19885
rect 36826 19821 36858 19885
rect 36922 19821 36954 19885
rect 35778 19791 36954 19821
rect 35778 19783 36570 19791
rect 31770 19753 36570 19783
rect 31770 19689 35426 19753
rect 35490 19689 35522 19753
rect 35586 19689 35618 19753
rect 35682 19689 35714 19753
rect 35778 19727 36570 19753
rect 36634 19727 36666 19791
rect 36730 19727 36762 19791
rect 36826 19727 36858 19791
rect 36922 19727 36954 19791
rect 35778 19689 36954 19727
rect 31770 19638 36954 19689
rect 969 19634 36954 19638
rect 0 19620 36954 19634
rect 36064 19577 36954 19620
rect 41602 19656 42660 19668
rect 37394 19551 37602 19585
rect 37394 19495 37427 19551
rect 37483 19495 37516 19551
rect 37572 19495 37602 19551
rect 36064 19462 36478 19485
rect 0 19451 36478 19462
rect 0 19196 1063 19451
rect 1445 19442 36478 19451
rect 1445 19386 1904 19442
rect 1960 19386 1998 19442
rect 2054 19386 2092 19442
rect 2148 19386 2604 19442
rect 2660 19386 2698 19442
rect 2754 19386 2792 19442
rect 2848 19386 5032 19442
rect 5088 19386 5126 19442
rect 5182 19386 5220 19442
rect 5276 19386 5904 19442
rect 5960 19386 5998 19442
rect 6054 19386 6092 19442
rect 6148 19386 6604 19442
rect 6660 19386 6698 19442
rect 6754 19386 6792 19442
rect 6848 19386 9032 19442
rect 9088 19386 9126 19442
rect 9182 19386 9220 19442
rect 9276 19386 9904 19442
rect 9960 19386 9998 19442
rect 10054 19386 10092 19442
rect 10148 19386 10604 19442
rect 10660 19386 10698 19442
rect 10754 19386 10792 19442
rect 10848 19386 13032 19442
rect 13088 19386 13126 19442
rect 13182 19386 13220 19442
rect 13276 19386 13904 19442
rect 13960 19386 13998 19442
rect 14054 19386 14092 19442
rect 14148 19386 14604 19442
rect 14660 19386 14698 19442
rect 14754 19386 14792 19442
rect 14848 19386 17032 19442
rect 17088 19386 17126 19442
rect 17182 19386 17220 19442
rect 17276 19386 17904 19442
rect 17960 19386 17998 19442
rect 18054 19386 18092 19442
rect 18148 19386 18604 19442
rect 18660 19386 18698 19442
rect 18754 19386 18792 19442
rect 18848 19386 21032 19442
rect 21088 19386 21126 19442
rect 21182 19386 21220 19442
rect 21276 19386 21904 19442
rect 21960 19386 21998 19442
rect 22054 19386 22092 19442
rect 22148 19386 22604 19442
rect 22660 19386 22698 19442
rect 22754 19386 22792 19442
rect 22848 19386 25032 19442
rect 25088 19386 25126 19442
rect 25182 19386 25220 19442
rect 25276 19386 25904 19442
rect 25960 19386 25998 19442
rect 26054 19386 26092 19442
rect 26148 19386 26604 19442
rect 26660 19386 26698 19442
rect 26754 19386 26792 19442
rect 26848 19386 29032 19442
rect 29088 19386 29126 19442
rect 29182 19386 29220 19442
rect 29276 19386 29904 19442
rect 29960 19386 29998 19442
rect 30054 19386 30092 19442
rect 30148 19386 30604 19442
rect 30660 19386 30698 19442
rect 30754 19386 30792 19442
rect 30848 19386 33032 19442
rect 33088 19386 33126 19442
rect 33182 19386 33220 19442
rect 33276 19386 33904 19442
rect 33960 19386 33998 19442
rect 34054 19386 34092 19442
rect 34148 19386 34604 19442
rect 34660 19386 34698 19442
rect 34754 19386 34792 19442
rect 34848 19386 36478 19442
rect 1445 19375 36478 19386
rect 1445 19348 36094 19375
rect 1445 19292 1904 19348
rect 1960 19292 1998 19348
rect 2054 19292 2092 19348
rect 2148 19292 2604 19348
rect 2660 19292 2698 19348
rect 2754 19292 2792 19348
rect 2848 19292 5032 19348
rect 5088 19292 5126 19348
rect 5182 19292 5220 19348
rect 5276 19292 5904 19348
rect 5960 19292 5998 19348
rect 6054 19292 6092 19348
rect 6148 19292 6604 19348
rect 6660 19292 6698 19348
rect 6754 19292 6792 19348
rect 6848 19292 9032 19348
rect 9088 19292 9126 19348
rect 9182 19292 9220 19348
rect 9276 19292 9904 19348
rect 9960 19292 9998 19348
rect 10054 19292 10092 19348
rect 10148 19292 10604 19348
rect 10660 19292 10698 19348
rect 10754 19292 10792 19348
rect 10848 19292 13032 19348
rect 13088 19292 13126 19348
rect 13182 19292 13220 19348
rect 13276 19292 13904 19348
rect 13960 19292 13998 19348
rect 14054 19292 14092 19348
rect 14148 19292 14604 19348
rect 14660 19292 14698 19348
rect 14754 19292 14792 19348
rect 14848 19292 17032 19348
rect 17088 19292 17126 19348
rect 17182 19292 17220 19348
rect 17276 19292 17904 19348
rect 17960 19292 17998 19348
rect 18054 19292 18092 19348
rect 18148 19292 18604 19348
rect 18660 19292 18698 19348
rect 18754 19292 18792 19348
rect 18848 19292 21032 19348
rect 21088 19292 21126 19348
rect 21182 19292 21220 19348
rect 21276 19292 21904 19348
rect 21960 19292 21998 19348
rect 22054 19292 22092 19348
rect 22148 19292 22604 19348
rect 22660 19292 22698 19348
rect 22754 19292 22792 19348
rect 22848 19292 25032 19348
rect 25088 19292 25126 19348
rect 25182 19292 25220 19348
rect 25276 19292 25904 19348
rect 25960 19292 25998 19348
rect 26054 19292 26092 19348
rect 26148 19292 26604 19348
rect 26660 19292 26698 19348
rect 26754 19292 26792 19348
rect 26848 19292 29032 19348
rect 29088 19292 29126 19348
rect 29182 19292 29220 19348
rect 29276 19292 29904 19348
rect 29960 19292 29998 19348
rect 30054 19292 30092 19348
rect 30148 19292 30604 19348
rect 30660 19292 30698 19348
rect 30754 19292 30792 19348
rect 30848 19292 33032 19348
rect 33088 19292 33126 19348
rect 33182 19292 33220 19348
rect 33276 19292 33904 19348
rect 33960 19292 33998 19348
rect 34054 19292 34092 19348
rect 34148 19292 34604 19348
rect 34660 19292 34698 19348
rect 34754 19292 34792 19348
rect 34848 19311 36094 19348
rect 36158 19311 36190 19375
rect 36254 19311 36286 19375
rect 36350 19311 36382 19375
rect 36446 19311 36478 19375
rect 34848 19292 36478 19311
rect 1445 19281 36478 19292
rect 37394 19460 37602 19495
rect 41602 19494 42410 19656
rect 42648 19494 42660 19656
rect 41602 19484 42660 19494
rect 37394 19404 37427 19460
rect 37483 19404 37516 19460
rect 37572 19404 37602 19460
rect 37394 19369 37602 19404
rect 37394 19313 37427 19369
rect 37483 19313 37516 19369
rect 37572 19313 37602 19369
rect 37394 19286 37602 19313
rect 1445 19254 36094 19281
rect 1445 19198 1904 19254
rect 1960 19198 1998 19254
rect 2054 19198 2092 19254
rect 2148 19198 2604 19254
rect 2660 19198 2698 19254
rect 2754 19198 2792 19254
rect 2848 19198 5032 19254
rect 5088 19198 5126 19254
rect 5182 19198 5220 19254
rect 5276 19198 5904 19254
rect 5960 19198 5998 19254
rect 6054 19198 6092 19254
rect 6148 19198 6604 19254
rect 6660 19198 6698 19254
rect 6754 19198 6792 19254
rect 6848 19198 9032 19254
rect 9088 19198 9126 19254
rect 9182 19198 9220 19254
rect 9276 19198 9904 19254
rect 9960 19198 9998 19254
rect 10054 19198 10092 19254
rect 10148 19198 10604 19254
rect 10660 19198 10698 19254
rect 10754 19198 10792 19254
rect 10848 19198 13032 19254
rect 13088 19198 13126 19254
rect 13182 19198 13220 19254
rect 13276 19198 13904 19254
rect 13960 19198 13998 19254
rect 14054 19198 14092 19254
rect 14148 19198 14604 19254
rect 14660 19198 14698 19254
rect 14754 19198 14792 19254
rect 14848 19198 17032 19254
rect 17088 19198 17126 19254
rect 17182 19198 17220 19254
rect 17276 19198 17904 19254
rect 17960 19198 17998 19254
rect 18054 19198 18092 19254
rect 18148 19198 18604 19254
rect 18660 19198 18698 19254
rect 18754 19198 18792 19254
rect 18848 19198 21032 19254
rect 21088 19198 21126 19254
rect 21182 19198 21220 19254
rect 21276 19198 21904 19254
rect 21960 19198 21998 19254
rect 22054 19198 22092 19254
rect 22148 19198 22604 19254
rect 22660 19198 22698 19254
rect 22754 19198 22792 19254
rect 22848 19198 25032 19254
rect 25088 19198 25126 19254
rect 25182 19198 25220 19254
rect 25276 19198 25904 19254
rect 25960 19198 25998 19254
rect 26054 19198 26092 19254
rect 26148 19198 26604 19254
rect 26660 19198 26698 19254
rect 26754 19198 26792 19254
rect 26848 19198 29032 19254
rect 29088 19198 29126 19254
rect 29182 19198 29220 19254
rect 29276 19198 29904 19254
rect 29960 19198 29998 19254
rect 30054 19198 30092 19254
rect 30148 19198 30604 19254
rect 30660 19198 30698 19254
rect 30754 19198 30792 19254
rect 30848 19198 33032 19254
rect 33088 19198 33126 19254
rect 33182 19198 33220 19254
rect 33276 19198 33904 19254
rect 33960 19198 33998 19254
rect 34054 19198 34092 19254
rect 34148 19198 34604 19254
rect 34660 19198 34698 19254
rect 34754 19198 34792 19254
rect 34848 19217 36094 19254
rect 36158 19217 36190 19281
rect 36254 19217 36286 19281
rect 36350 19217 36382 19281
rect 36446 19217 36478 19281
rect 42396 19250 42660 19276
rect 34848 19198 36478 19217
rect 1445 19196 36478 19198
rect 0 19182 36478 19196
rect 37444 19212 37602 19227
rect 37444 19160 37451 19212
rect 37503 19160 37542 19212
rect 37594 19160 37602 19212
rect 37444 19110 37602 19160
rect 37444 19058 37451 19110
rect 37503 19058 37542 19110
rect 37594 19058 37602 19110
rect 37444 19007 37602 19058
rect 37444 18955 37452 19007
rect 37504 18955 37543 19007
rect 37595 18955 37602 19007
rect 37444 18914 37602 18955
rect 36540 18870 36954 18890
rect 36540 18836 36561 18870
rect 570 18816 1700 18836
rect 570 18745 591 18816
rect 662 18745 686 18816
rect 757 18745 795 18816
rect 866 18745 890 18816
rect 961 18780 1700 18816
rect 35836 18799 36561 18836
rect 36632 18799 36656 18870
rect 36727 18799 36765 18870
rect 36836 18799 36860 18870
rect 36931 18799 36954 18870
rect 37444 18862 37452 18914
rect 37504 18862 37543 18914
rect 37595 18862 37602 18914
rect 37444 18849 37602 18862
rect 42396 18838 42422 19250
rect 42634 18838 42660 19250
rect 42396 18814 42660 18838
rect 35836 18780 36954 18799
rect 41602 18788 42164 18806
rect 961 18752 984 18780
rect 961 18745 1700 18752
rect 570 18726 1700 18745
rect 620 18724 1700 18726
rect 620 18696 918 18724
rect 41602 18638 41930 18788
rect 42142 18638 42164 18788
rect 41602 18624 42164 18638
rect 570 18502 1700 18522
rect 570 18431 591 18502
rect 662 18431 686 18502
rect 757 18431 795 18502
rect 866 18431 890 18502
rect 961 18494 1700 18502
rect 961 18440 984 18494
rect 961 18431 1700 18440
rect 570 18412 1700 18431
rect 1046 18363 1700 18384
rect 1046 18292 1067 18363
rect 1138 18292 1162 18363
rect 1233 18292 1271 18363
rect 1342 18292 1366 18363
rect 1437 18356 1700 18363
rect 1437 18292 1460 18356
rect 1046 18273 1460 18292
rect 37042 18297 37364 18312
rect 37042 18259 37061 18297
rect 398 18190 404 18242
rect 460 18190 472 18242
rect 528 18230 570 18242
rect 528 18202 1700 18230
rect 35836 18217 37061 18259
rect 37148 18217 37161 18297
rect 37248 18217 37261 18297
rect 37348 18217 37364 18297
rect 35836 18202 37364 18217
rect 41602 18246 42164 18264
rect 528 18190 570 18202
rect 1046 18153 1700 18174
rect 1046 18082 1067 18153
rect 1138 18082 1162 18153
rect 1233 18082 1271 18153
rect 1342 18082 1366 18153
rect 1437 18118 1700 18153
rect 35836 18154 36478 18174
rect 35836 18118 36085 18154
rect 1437 18082 1460 18118
rect 1046 18063 1460 18082
rect 36064 18083 36085 18118
rect 36156 18083 36180 18154
rect 36251 18083 36289 18154
rect 36360 18083 36384 18154
rect 36455 18083 36478 18154
rect 36064 18064 36478 18083
rect 41602 18096 41930 18246
rect 42142 18096 42164 18246
rect 41602 18082 42164 18096
rect 570 17866 984 17886
rect 570 17795 591 17866
rect 662 17795 686 17866
rect 757 17795 795 17866
rect 866 17795 890 17866
rect 961 17832 984 17866
rect 36540 17866 36954 17886
rect 36540 17832 36561 17866
rect 961 17795 1700 17832
rect 570 17776 1700 17795
rect 35836 17795 36561 17832
rect 36632 17795 36656 17866
rect 36727 17795 36765 17866
rect 36836 17795 36860 17866
rect 36931 17795 36954 17866
rect 35836 17776 36954 17795
rect 182 17696 188 17748
rect 244 17720 1700 17748
rect 244 17696 250 17720
rect 41602 17690 42164 17708
rect 41602 17540 41930 17690
rect 42142 17540 42164 17690
rect 41602 17526 42164 17540
rect 0 17490 1700 17518
rect 42396 17492 42660 17518
rect 37444 17452 37602 17467
rect 0 17408 1700 17436
rect 37444 17400 37451 17452
rect 37503 17400 37542 17452
rect 37594 17400 37602 17452
rect 290 17328 296 17380
rect 352 17352 1700 17380
rect 352 17328 358 17352
rect 37444 17350 37602 17400
rect 37042 17293 37364 17308
rect 37042 17255 37061 17293
rect 398 17186 410 17238
rect 524 17226 570 17238
rect 524 17198 1700 17226
rect 35836 17213 37061 17255
rect 37148 17213 37161 17293
rect 37248 17213 37261 17293
rect 37348 17213 37364 17293
rect 35836 17198 37364 17213
rect 37444 17298 37451 17350
rect 37503 17298 37542 17350
rect 37594 17298 37602 17350
rect 37444 17247 37602 17298
rect 524 17186 570 17198
rect 37444 17195 37452 17247
rect 37504 17195 37543 17247
rect 37595 17195 37602 17247
rect 1046 17150 1700 17170
rect 1046 17079 1067 17150
rect 1138 17079 1162 17150
rect 1233 17079 1271 17150
rect 1342 17079 1366 17150
rect 1437 17114 1700 17150
rect 35836 17150 36478 17170
rect 35836 17114 36085 17150
rect 1437 17079 1460 17114
rect 1046 17060 1460 17079
rect 36064 17079 36085 17114
rect 36156 17079 36180 17150
rect 36251 17079 36289 17150
rect 36360 17079 36384 17150
rect 36455 17079 36478 17150
rect 37444 17154 37602 17195
rect 37444 17102 37452 17154
rect 37504 17102 37543 17154
rect 37595 17102 37602 17154
rect 37444 17089 37602 17102
rect 36064 17060 36478 17079
rect 42396 17080 42422 17492
rect 42634 17080 42660 17492
rect 42396 17056 42660 17080
rect 570 16862 984 16882
rect 570 16791 591 16862
rect 662 16791 686 16862
rect 757 16791 795 16862
rect 866 16791 890 16862
rect 961 16828 984 16862
rect 36540 16862 36954 16882
rect 36540 16828 36561 16862
rect 961 16791 1700 16828
rect 570 16772 1700 16791
rect 35836 16791 36561 16828
rect 36632 16791 36656 16862
rect 36727 16791 36765 16862
rect 36836 16791 36860 16862
rect 36931 16791 36954 16862
rect 35836 16772 36954 16791
rect 182 16692 188 16744
rect 244 16716 1700 16744
rect 244 16692 250 16716
rect 37394 16646 37602 16680
rect 37394 16590 37427 16646
rect 37483 16590 37516 16646
rect 37572 16590 37602 16646
rect 37394 16555 37602 16590
rect 0 16486 1700 16514
rect 37394 16499 37427 16555
rect 37483 16499 37516 16555
rect 37572 16499 37602 16555
rect 37394 16464 37602 16499
rect 0 16404 1700 16432
rect 37394 16408 37427 16464
rect 37483 16408 37516 16464
rect 37572 16408 37602 16464
rect 37394 16381 37602 16408
rect 41602 16546 42660 16558
rect 41602 16384 42410 16546
rect 42648 16384 42660 16546
rect 290 16324 296 16376
rect 352 16348 1700 16376
rect 41602 16374 42660 16384
rect 352 16324 358 16348
rect 37042 16289 37364 16304
rect 37042 16251 37061 16289
rect 398 16182 410 16234
rect 524 16222 570 16234
rect 524 16194 1700 16222
rect 35836 16209 37061 16251
rect 37148 16209 37161 16289
rect 37248 16209 37261 16289
rect 37348 16209 37364 16289
rect 35836 16194 37364 16209
rect 524 16182 570 16194
rect 1046 16145 1700 16166
rect 1046 16074 1067 16145
rect 1138 16074 1162 16145
rect 1233 16074 1271 16145
rect 1342 16074 1366 16145
rect 1437 16110 1700 16145
rect 35836 16146 36478 16166
rect 35836 16110 36085 16146
rect 1437 16074 1460 16110
rect 1046 16055 1460 16074
rect 36064 16075 36085 16110
rect 36156 16075 36180 16146
rect 36251 16075 36289 16146
rect 36360 16075 36384 16146
rect 36455 16075 36478 16146
rect 36064 16056 36478 16075
rect 570 15858 984 15878
rect 570 15787 591 15858
rect 662 15787 686 15858
rect 757 15787 795 15858
rect 866 15787 890 15858
rect 961 15824 984 15858
rect 36540 15858 36954 15878
rect 36540 15824 36561 15858
rect 961 15787 1700 15824
rect 570 15768 1700 15787
rect 35836 15787 36561 15824
rect 36632 15787 36656 15858
rect 36727 15787 36765 15858
rect 36836 15787 36860 15858
rect 36931 15787 36954 15858
rect 35836 15768 36954 15787
rect 182 15688 188 15740
rect 244 15712 1700 15740
rect 244 15688 250 15712
rect 41602 15656 42660 15668
rect 0 15482 1700 15510
rect 41602 15494 42410 15656
rect 42648 15494 42660 15656
rect 41602 15484 42660 15494
rect 0 15400 1700 15428
rect 290 15320 296 15372
rect 352 15344 1700 15372
rect 352 15320 358 15344
rect 37042 15285 37364 15300
rect 37042 15247 37061 15285
rect 398 15178 410 15230
rect 524 15218 570 15230
rect 524 15190 1700 15218
rect 35836 15205 37061 15247
rect 37148 15205 37161 15285
rect 37248 15205 37261 15285
rect 37348 15205 37364 15285
rect 42396 15250 42660 15276
rect 35836 15190 37364 15205
rect 37444 15212 37602 15227
rect 524 15178 570 15190
rect 1046 15142 1700 15162
rect 1046 15071 1067 15142
rect 1138 15071 1162 15142
rect 1233 15071 1271 15142
rect 1342 15071 1366 15142
rect 1437 15106 1700 15142
rect 35836 15142 36478 15162
rect 35836 15106 36085 15142
rect 1437 15071 1460 15106
rect 1046 15052 1460 15071
rect 36064 15071 36085 15106
rect 36156 15071 36180 15142
rect 36251 15071 36289 15142
rect 36360 15071 36384 15142
rect 36455 15071 36478 15142
rect 36064 15052 36478 15071
rect 37444 15160 37451 15212
rect 37503 15160 37542 15212
rect 37594 15160 37602 15212
rect 37444 15110 37602 15160
rect 37444 15058 37451 15110
rect 37503 15058 37542 15110
rect 37594 15058 37602 15110
rect 37444 15007 37602 15058
rect 37444 14955 37452 15007
rect 37504 14955 37543 15007
rect 37595 14955 37602 15007
rect 37444 14914 37602 14955
rect 570 14854 984 14874
rect 570 14783 591 14854
rect 662 14783 686 14854
rect 757 14783 795 14854
rect 866 14783 890 14854
rect 961 14820 984 14854
rect 36540 14854 36954 14874
rect 36540 14820 36561 14854
rect 961 14783 1700 14820
rect 570 14764 1700 14783
rect 35836 14783 36561 14820
rect 36632 14783 36656 14854
rect 36727 14783 36765 14854
rect 36836 14783 36860 14854
rect 36931 14783 36954 14854
rect 37444 14862 37452 14914
rect 37504 14862 37543 14914
rect 37595 14862 37602 14914
rect 37444 14849 37602 14862
rect 42396 14838 42422 15250
rect 42634 14838 42660 15250
rect 42396 14814 42660 14838
rect 35836 14764 36954 14783
rect 41602 14788 42164 14806
rect 182 14684 188 14736
rect 244 14708 1700 14736
rect 244 14684 250 14708
rect 41602 14638 41930 14788
rect 42142 14638 42164 14788
rect 41602 14624 42164 14638
rect 0 14478 1700 14506
rect 0 14396 1700 14424
rect 290 14316 296 14368
rect 352 14340 1700 14368
rect 352 14316 358 14340
rect 37042 14281 37364 14296
rect 37042 14243 37061 14281
rect 398 14174 410 14226
rect 524 14214 570 14226
rect 524 14186 1700 14214
rect 35836 14201 37061 14243
rect 37148 14201 37161 14281
rect 37248 14201 37261 14281
rect 37348 14201 37364 14281
rect 35836 14186 37364 14201
rect 41602 14246 42164 14264
rect 524 14174 570 14186
rect 1046 14138 1700 14158
rect 1046 14067 1067 14138
rect 1138 14067 1162 14138
rect 1233 14067 1271 14138
rect 1342 14067 1366 14138
rect 1437 14102 1700 14138
rect 35836 14138 36478 14158
rect 35836 14102 36085 14138
rect 1437 14067 1460 14102
rect 1046 14048 1460 14067
rect 36064 14067 36085 14102
rect 36156 14067 36180 14138
rect 36251 14067 36289 14138
rect 36360 14067 36384 14138
rect 36455 14067 36478 14138
rect 41602 14096 41930 14246
rect 42142 14096 42164 14246
rect 41602 14082 42164 14096
rect 36064 14048 36478 14067
rect 570 13850 984 13870
rect 570 13779 591 13850
rect 662 13779 686 13850
rect 757 13779 795 13850
rect 866 13779 890 13850
rect 961 13816 984 13850
rect 36540 13850 36954 13870
rect 36540 13816 36561 13850
rect 961 13779 1700 13816
rect 570 13760 1700 13779
rect 35836 13779 36561 13816
rect 36632 13779 36656 13850
rect 36727 13779 36765 13850
rect 36836 13779 36860 13850
rect 36931 13779 36954 13850
rect 35836 13760 36954 13779
rect 182 13680 188 13732
rect 244 13704 1700 13732
rect 244 13680 250 13704
rect 41602 13690 42164 13708
rect 41602 13540 41930 13690
rect 42142 13540 42164 13690
rect 41602 13526 42164 13540
rect 0 13474 1700 13502
rect 42396 13492 42660 13518
rect 37444 13452 37602 13467
rect 0 13392 1700 13420
rect 37444 13400 37451 13452
rect 37503 13400 37542 13452
rect 37594 13400 37602 13452
rect 290 13312 296 13364
rect 352 13336 1700 13364
rect 37444 13350 37602 13400
rect 352 13312 358 13336
rect 37444 13298 37451 13350
rect 37503 13298 37542 13350
rect 37594 13298 37602 13350
rect 37042 13277 37364 13292
rect 37042 13239 37061 13277
rect 398 13170 410 13222
rect 524 13210 570 13222
rect 524 13182 1700 13210
rect 35836 13197 37061 13239
rect 37148 13197 37161 13277
rect 37248 13197 37261 13277
rect 37348 13197 37364 13277
rect 35836 13182 37364 13197
rect 37444 13247 37602 13298
rect 37444 13195 37452 13247
rect 37504 13195 37543 13247
rect 37595 13195 37602 13247
rect 524 13170 570 13182
rect 37444 13154 37602 13195
rect 1046 13134 1700 13154
rect 1046 13063 1067 13134
rect 1138 13063 1162 13134
rect 1233 13063 1271 13134
rect 1342 13063 1366 13134
rect 1437 13098 1700 13134
rect 35836 13134 36478 13154
rect 35836 13098 36085 13134
rect 1437 13063 1460 13098
rect 1046 13044 1460 13063
rect 36064 13063 36085 13098
rect 36156 13063 36180 13134
rect 36251 13063 36289 13134
rect 36360 13063 36384 13134
rect 36455 13063 36478 13134
rect 37444 13102 37452 13154
rect 37504 13102 37543 13154
rect 37595 13102 37602 13154
rect 37444 13089 37602 13102
rect 36064 13044 36478 13063
rect 42396 13080 42422 13492
rect 42634 13080 42660 13492
rect 42396 13056 42660 13080
rect 570 12846 984 12866
rect 570 12775 591 12846
rect 662 12775 686 12846
rect 757 12775 795 12846
rect 866 12775 890 12846
rect 961 12812 984 12846
rect 36540 12846 36954 12866
rect 36540 12812 36561 12846
rect 961 12775 1700 12812
rect 570 12756 1700 12775
rect 35836 12775 36561 12812
rect 36632 12775 36656 12846
rect 36727 12775 36765 12846
rect 36836 12775 36860 12846
rect 36931 12775 36954 12846
rect 35836 12756 36954 12775
rect 182 12676 188 12728
rect 244 12700 1700 12728
rect 244 12676 250 12700
rect 37394 12588 37602 12622
rect 37394 12532 37427 12588
rect 37483 12532 37516 12588
rect 37572 12532 37602 12588
rect 0 12470 1700 12498
rect 37394 12497 37602 12532
rect 37394 12441 37427 12497
rect 37483 12441 37516 12497
rect 37572 12441 37602 12497
rect 0 12388 1700 12416
rect 37394 12406 37602 12441
rect 290 12308 296 12360
rect 352 12332 1700 12360
rect 37394 12350 37427 12406
rect 37483 12350 37516 12406
rect 37572 12350 37602 12406
rect 41602 12546 42660 12558
rect 41602 12384 42410 12546
rect 42648 12384 42660 12546
rect 41602 12374 42660 12384
rect 352 12308 358 12332
rect 37394 12323 37602 12350
rect 37042 12273 37364 12288
rect 37042 12235 37061 12273
rect 398 12166 410 12218
rect 524 12206 570 12218
rect 524 12178 1700 12206
rect 35836 12193 37061 12235
rect 37148 12193 37161 12273
rect 37248 12193 37261 12273
rect 37348 12193 37364 12273
rect 35836 12178 37364 12193
rect 524 12166 570 12178
rect 1046 12130 1700 12150
rect 1046 12059 1067 12130
rect 1138 12059 1162 12130
rect 1233 12059 1271 12130
rect 1342 12059 1366 12130
rect 1437 12094 1700 12130
rect 35836 12130 36478 12150
rect 35836 12094 36085 12130
rect 1437 12059 1460 12094
rect 1046 12040 1460 12059
rect 36064 12059 36085 12094
rect 36156 12059 36180 12130
rect 36251 12059 36289 12130
rect 36360 12059 36384 12130
rect 36455 12059 36478 12130
rect 36064 12040 36478 12059
rect 570 11842 984 11862
rect 570 11771 591 11842
rect 662 11771 686 11842
rect 757 11771 795 11842
rect 866 11771 890 11842
rect 961 11808 984 11842
rect 36540 11842 36954 11862
rect 36540 11808 36561 11842
rect 961 11771 1700 11808
rect 570 11752 1700 11771
rect 35836 11771 36561 11808
rect 36632 11771 36656 11842
rect 36727 11771 36765 11842
rect 36836 11771 36860 11842
rect 36931 11771 36954 11842
rect 35836 11752 36954 11771
rect 182 11672 188 11724
rect 244 11696 1700 11724
rect 244 11672 250 11696
rect 41602 11656 42660 11668
rect 41602 11494 42410 11656
rect 42648 11494 42660 11656
rect 0 11466 1700 11494
rect 41602 11484 42660 11494
rect 0 11384 1700 11412
rect 290 11304 296 11356
rect 352 11328 1700 11356
rect 352 11304 358 11328
rect 37042 11269 37364 11284
rect 37042 11231 37061 11269
rect 398 11162 410 11214
rect 524 11202 570 11214
rect 524 11174 1700 11202
rect 35836 11189 37061 11231
rect 37148 11189 37161 11269
rect 37248 11189 37261 11269
rect 37348 11189 37364 11269
rect 42396 11250 42660 11276
rect 35836 11174 37364 11189
rect 37444 11212 37602 11227
rect 524 11162 570 11174
rect 37444 11160 37451 11212
rect 37503 11160 37542 11212
rect 37594 11160 37602 11212
rect 1046 11126 1700 11146
rect 1046 11055 1067 11126
rect 1138 11055 1162 11126
rect 1233 11055 1271 11126
rect 1342 11055 1366 11126
rect 1437 11090 1700 11126
rect 35836 11126 36478 11146
rect 35836 11090 36085 11126
rect 1437 11055 1460 11090
rect 1046 11036 1460 11055
rect 36064 11055 36085 11090
rect 36156 11055 36180 11126
rect 36251 11055 36289 11126
rect 36360 11055 36384 11126
rect 36455 11055 36478 11126
rect 36064 11036 36478 11055
rect 37444 11110 37602 11160
rect 37444 11058 37451 11110
rect 37503 11058 37542 11110
rect 37594 11058 37602 11110
rect 37444 11007 37602 11058
rect 37444 10955 37452 11007
rect 37504 10955 37543 11007
rect 37595 10955 37602 11007
rect 37444 10914 37602 10955
rect 37444 10862 37452 10914
rect 37504 10862 37543 10914
rect 37595 10862 37602 10914
rect 570 10838 984 10858
rect 570 10767 591 10838
rect 662 10767 686 10838
rect 757 10767 795 10838
rect 866 10767 890 10838
rect 961 10804 984 10838
rect 36540 10838 36954 10858
rect 37444 10849 37602 10862
rect 36540 10804 36561 10838
rect 961 10767 1700 10804
rect 570 10748 1700 10767
rect 35836 10767 36561 10804
rect 36632 10767 36656 10838
rect 36727 10767 36765 10838
rect 36836 10767 36860 10838
rect 36931 10767 36954 10838
rect 42396 10838 42422 11250
rect 42634 10838 42660 11250
rect 42396 10814 42660 10838
rect 35836 10748 36954 10767
rect 41602 10788 42164 10806
rect 182 10668 188 10720
rect 244 10692 1700 10720
rect 244 10668 250 10692
rect 41602 10638 41930 10788
rect 42142 10638 42164 10788
rect 41602 10624 42164 10638
rect 0 10462 1700 10490
rect 0 10380 1700 10408
rect 290 10300 296 10352
rect 352 10324 1700 10352
rect 352 10300 358 10324
rect 37042 10265 37364 10280
rect 37042 10227 37061 10265
rect 398 10158 410 10210
rect 524 10198 570 10210
rect 524 10170 1700 10198
rect 35836 10185 37061 10227
rect 37148 10185 37161 10265
rect 37248 10185 37261 10265
rect 37348 10185 37364 10265
rect 35836 10170 37364 10185
rect 41602 10246 42164 10264
rect 524 10158 570 10170
rect 1046 10122 1700 10142
rect 1046 10051 1067 10122
rect 1138 10051 1162 10122
rect 1233 10051 1271 10122
rect 1342 10051 1366 10122
rect 1437 10086 1700 10122
rect 35836 10122 36478 10142
rect 35836 10086 36085 10122
rect 1437 10051 1460 10086
rect 1046 10032 1460 10051
rect 36064 10051 36085 10086
rect 36156 10051 36180 10122
rect 36251 10051 36289 10122
rect 36360 10051 36384 10122
rect 36455 10051 36478 10122
rect 41602 10096 41930 10246
rect 42142 10096 42164 10246
rect 41602 10082 42164 10096
rect 36064 10032 36478 10051
rect 570 9834 984 9854
rect 570 9763 591 9834
rect 662 9763 686 9834
rect 757 9763 795 9834
rect 866 9763 890 9834
rect 961 9800 984 9834
rect 36540 9834 36954 9854
rect 36540 9800 36561 9834
rect 961 9763 1700 9800
rect 570 9744 1700 9763
rect 35836 9763 36561 9800
rect 36632 9763 36656 9834
rect 36727 9763 36765 9834
rect 36836 9763 36860 9834
rect 36931 9763 36954 9834
rect 35836 9744 36954 9763
rect 182 9664 188 9716
rect 244 9688 1700 9716
rect 41602 9690 42164 9708
rect 244 9664 250 9688
rect 41602 9540 41930 9690
rect 42142 9540 42164 9690
rect 41602 9526 42164 9540
rect 42396 9492 42660 9518
rect 0 9458 1700 9486
rect 37444 9452 37602 9467
rect 0 9376 1700 9404
rect 37444 9400 37451 9452
rect 37503 9400 37542 9452
rect 37594 9400 37602 9452
rect 37444 9350 37602 9400
rect 290 9296 296 9348
rect 352 9320 1700 9348
rect 352 9296 358 9320
rect 37444 9298 37451 9350
rect 37503 9298 37542 9350
rect 37594 9298 37602 9350
rect 37042 9261 37364 9276
rect 37042 9223 37061 9261
rect 398 9154 410 9206
rect 524 9194 570 9206
rect 524 9166 1700 9194
rect 35836 9181 37061 9223
rect 37148 9181 37161 9261
rect 37248 9181 37261 9261
rect 37348 9181 37364 9261
rect 35836 9166 37364 9181
rect 37444 9247 37602 9298
rect 37444 9195 37452 9247
rect 37504 9195 37543 9247
rect 37595 9195 37602 9247
rect 524 9154 570 9166
rect 37444 9154 37602 9195
rect 1046 9118 1700 9138
rect 1046 9047 1067 9118
rect 1138 9047 1162 9118
rect 1233 9047 1271 9118
rect 1342 9047 1366 9118
rect 1437 9082 1700 9118
rect 35836 9118 36478 9138
rect 35836 9082 36085 9118
rect 1437 9047 1460 9082
rect 1046 9028 1460 9047
rect 36064 9047 36085 9082
rect 36156 9047 36180 9118
rect 36251 9047 36289 9118
rect 36360 9047 36384 9118
rect 36455 9047 36478 9118
rect 37444 9102 37452 9154
rect 37504 9102 37543 9154
rect 37595 9102 37602 9154
rect 37444 9089 37602 9102
rect 42396 9080 42422 9492
rect 42634 9080 42660 9492
rect 42396 9056 42660 9080
rect 36064 9028 36478 9047
rect 570 8830 984 8850
rect 570 8759 591 8830
rect 662 8759 686 8830
rect 757 8759 795 8830
rect 866 8759 890 8830
rect 961 8796 984 8830
rect 36540 8830 36954 8850
rect 36540 8796 36561 8830
rect 961 8759 1700 8796
rect 570 8740 1700 8759
rect 35836 8759 36561 8796
rect 36632 8759 36656 8830
rect 36727 8759 36765 8830
rect 36836 8759 36860 8830
rect 36931 8759 36954 8830
rect 35836 8740 36954 8759
rect 182 8660 188 8712
rect 244 8684 1700 8712
rect 244 8660 250 8684
rect 41602 8546 42660 8558
rect 37394 8495 37602 8529
rect 0 8454 1700 8482
rect 37394 8439 37427 8495
rect 37483 8439 37516 8495
rect 37572 8439 37602 8495
rect 37394 8404 37602 8439
rect 0 8372 1700 8400
rect 37394 8348 37427 8404
rect 37483 8348 37516 8404
rect 37572 8348 37602 8404
rect 41602 8384 42410 8546
rect 42648 8384 42660 8546
rect 41602 8374 42660 8384
rect 290 8292 296 8344
rect 352 8316 1700 8344
rect 352 8292 358 8316
rect 37394 8313 37602 8348
rect 37042 8257 37364 8272
rect 37042 8219 37061 8257
rect 398 8150 410 8202
rect 524 8190 570 8202
rect 524 8162 1700 8190
rect 35836 8177 37061 8219
rect 37148 8177 37161 8257
rect 37248 8177 37261 8257
rect 37348 8177 37364 8257
rect 37394 8257 37427 8313
rect 37483 8257 37516 8313
rect 37572 8257 37602 8313
rect 37394 8230 37602 8257
rect 35836 8162 37364 8177
rect 524 8150 570 8162
rect 1046 8114 1700 8134
rect 1046 8043 1067 8114
rect 1138 8043 1162 8114
rect 1233 8043 1271 8114
rect 1342 8043 1366 8114
rect 1437 8078 1700 8114
rect 35836 8114 36478 8134
rect 35836 8078 36085 8114
rect 1437 8043 1460 8078
rect 1046 8024 1460 8043
rect 36064 8043 36085 8078
rect 36156 8043 36180 8114
rect 36251 8043 36289 8114
rect 36360 8043 36384 8114
rect 36455 8043 36478 8114
rect 36064 8024 36478 8043
rect 570 7826 984 7846
rect 570 7755 591 7826
rect 662 7755 686 7826
rect 757 7755 795 7826
rect 866 7755 890 7826
rect 961 7792 984 7826
rect 36540 7826 36954 7846
rect 36540 7792 36561 7826
rect 961 7755 1700 7792
rect 570 7736 1700 7755
rect 35836 7755 36561 7792
rect 36632 7755 36656 7826
rect 36727 7755 36765 7826
rect 36836 7755 36860 7826
rect 36931 7755 36954 7826
rect 35836 7736 36954 7755
rect 182 7656 188 7708
rect 244 7680 1700 7708
rect 244 7656 250 7680
rect 41602 7656 42660 7668
rect 41602 7494 42410 7656
rect 42648 7494 42660 7656
rect 41602 7484 42660 7494
rect 0 7450 1700 7478
rect 0 7368 1700 7396
rect 290 7288 296 7340
rect 352 7312 1700 7340
rect 352 7288 358 7312
rect 37042 7253 37364 7268
rect 37042 7215 37061 7253
rect 398 7146 410 7198
rect 524 7186 570 7198
rect 524 7158 1700 7186
rect 35836 7173 37061 7215
rect 37148 7173 37161 7253
rect 37248 7173 37261 7253
rect 37348 7173 37364 7253
rect 42396 7250 42660 7276
rect 35836 7158 37364 7173
rect 37444 7212 37602 7227
rect 37444 7160 37451 7212
rect 37503 7160 37542 7212
rect 37594 7160 37602 7212
rect 524 7146 570 7158
rect 1046 7110 1700 7130
rect 1046 7039 1067 7110
rect 1138 7039 1162 7110
rect 1233 7039 1271 7110
rect 1342 7039 1366 7110
rect 1437 7074 1700 7110
rect 35836 7110 36478 7130
rect 35836 7074 36085 7110
rect 1437 7039 1460 7074
rect 1046 7020 1460 7039
rect 36064 7039 36085 7074
rect 36156 7039 36180 7110
rect 36251 7039 36289 7110
rect 36360 7039 36384 7110
rect 36455 7039 36478 7110
rect 36064 7020 36478 7039
rect 37444 7110 37602 7160
rect 37444 7058 37451 7110
rect 37503 7058 37542 7110
rect 37594 7058 37602 7110
rect 37444 7007 37602 7058
rect 37444 6955 37452 7007
rect 37504 6955 37543 7007
rect 37595 6955 37602 7007
rect 37444 6914 37602 6955
rect 37444 6862 37452 6914
rect 37504 6862 37543 6914
rect 37595 6862 37602 6914
rect 37444 6849 37602 6862
rect 570 6822 984 6842
rect 570 6751 591 6822
rect 662 6751 686 6822
rect 757 6751 795 6822
rect 866 6751 890 6822
rect 961 6788 984 6822
rect 36540 6822 36954 6842
rect 36540 6788 36561 6822
rect 961 6751 1700 6788
rect 570 6732 1700 6751
rect 35836 6751 36561 6788
rect 36632 6751 36656 6822
rect 36727 6751 36765 6822
rect 36836 6751 36860 6822
rect 36931 6751 36954 6822
rect 42396 6838 42422 7250
rect 42634 6838 42660 7250
rect 42396 6814 42660 6838
rect 35836 6732 36954 6751
rect 41602 6788 42164 6806
rect 182 6652 188 6704
rect 244 6676 1700 6704
rect 244 6652 250 6676
rect 41602 6638 41930 6788
rect 42142 6638 42164 6788
rect 41602 6624 42164 6638
rect 0 6446 1700 6474
rect 0 6364 1700 6392
rect 290 6284 296 6336
rect 352 6308 1700 6336
rect 352 6284 358 6308
rect 37042 6249 37364 6264
rect 37042 6211 37061 6249
rect 398 6142 410 6194
rect 524 6182 570 6194
rect 524 6154 1700 6182
rect 35836 6169 37061 6211
rect 37148 6169 37161 6249
rect 37248 6169 37261 6249
rect 37348 6169 37364 6249
rect 35836 6154 37364 6169
rect 41602 6246 42164 6264
rect 524 6142 570 6154
rect 1046 6106 1700 6126
rect 1046 6035 1067 6106
rect 1138 6035 1162 6106
rect 1233 6035 1271 6106
rect 1342 6035 1366 6106
rect 1437 6070 1700 6106
rect 35836 6106 36478 6126
rect 35836 6070 36085 6106
rect 1437 6035 1460 6070
rect 1046 6016 1460 6035
rect 36064 6035 36085 6070
rect 36156 6035 36180 6106
rect 36251 6035 36289 6106
rect 36360 6035 36384 6106
rect 36455 6035 36478 6106
rect 41602 6096 41930 6246
rect 42142 6096 42164 6246
rect 41602 6082 42164 6096
rect 36064 6016 36478 6035
rect 570 5818 984 5838
rect 570 5747 591 5818
rect 662 5747 686 5818
rect 757 5747 795 5818
rect 866 5747 890 5818
rect 961 5784 984 5818
rect 36540 5818 36954 5838
rect 36540 5784 36561 5818
rect 961 5747 1700 5784
rect 570 5728 1700 5747
rect 35836 5747 36561 5784
rect 36632 5747 36656 5818
rect 36727 5747 36765 5818
rect 36836 5747 36860 5818
rect 36931 5747 36954 5818
rect 35836 5728 36954 5747
rect 182 5648 188 5700
rect 244 5672 1700 5700
rect 41602 5690 42164 5708
rect 244 5648 250 5672
rect 41602 5540 41930 5690
rect 42142 5540 42164 5690
rect 41602 5526 42164 5540
rect 42396 5492 42660 5518
rect 0 5442 1700 5470
rect 37444 5452 37602 5467
rect 37444 5400 37451 5452
rect 37503 5400 37542 5452
rect 37594 5400 37602 5452
rect 0 5360 1700 5388
rect 37444 5350 37602 5400
rect 290 5280 296 5332
rect 352 5304 1700 5332
rect 352 5280 358 5304
rect 37444 5298 37451 5350
rect 37503 5298 37542 5350
rect 37594 5298 37602 5350
rect 37042 5245 37364 5260
rect 37042 5207 37061 5245
rect 398 5138 410 5190
rect 524 5178 570 5190
rect 524 5150 1700 5178
rect 35836 5165 37061 5207
rect 37148 5165 37161 5245
rect 37248 5165 37261 5245
rect 37348 5165 37364 5245
rect 35836 5150 37364 5165
rect 37444 5247 37602 5298
rect 37444 5195 37452 5247
rect 37504 5195 37543 5247
rect 37595 5195 37602 5247
rect 37444 5154 37602 5195
rect 524 5138 570 5150
rect 1046 5102 1700 5122
rect 1046 5031 1067 5102
rect 1138 5031 1162 5102
rect 1233 5031 1271 5102
rect 1342 5031 1366 5102
rect 1437 5066 1700 5102
rect 35836 5102 36478 5122
rect 35836 5066 36085 5102
rect 1437 5031 1460 5066
rect 1046 5012 1460 5031
rect 36064 5031 36085 5066
rect 36156 5031 36180 5102
rect 36251 5031 36289 5102
rect 36360 5031 36384 5102
rect 36455 5031 36478 5102
rect 37444 5102 37452 5154
rect 37504 5102 37543 5154
rect 37595 5102 37602 5154
rect 37444 5089 37602 5102
rect 42396 5080 42422 5492
rect 42634 5080 42660 5492
rect 42396 5056 42660 5080
rect 36064 5012 36478 5031
rect 570 4814 984 4834
rect 570 4743 591 4814
rect 662 4743 686 4814
rect 757 4743 795 4814
rect 866 4743 890 4814
rect 961 4780 984 4814
rect 36540 4814 36954 4834
rect 36540 4780 36561 4814
rect 961 4743 1700 4780
rect 570 4724 1700 4743
rect 35836 4743 36561 4780
rect 36632 4743 36656 4814
rect 36727 4743 36765 4814
rect 36836 4743 36860 4814
rect 36931 4743 36954 4814
rect 35836 4724 36954 4743
rect 182 4644 188 4696
rect 244 4668 1700 4696
rect 244 4644 250 4668
rect 41602 4546 42660 4558
rect 0 4438 1700 4466
rect 41602 4384 42410 4546
rect 42648 4384 42660 4546
rect 0 4356 1700 4384
rect 41602 4374 42660 4384
rect 290 4276 296 4328
rect 352 4300 1700 4328
rect 352 4276 358 4300
rect 37042 4241 37364 4256
rect 37042 4203 37061 4241
rect 398 4134 410 4186
rect 524 4174 570 4186
rect 524 4146 1700 4174
rect 35836 4161 37061 4203
rect 37148 4161 37161 4241
rect 37248 4161 37261 4241
rect 37348 4161 37364 4241
rect 35836 4146 37364 4161
rect 524 4134 570 4146
rect 1046 4098 1700 4118
rect 1046 4027 1067 4098
rect 1138 4027 1162 4098
rect 1233 4027 1271 4098
rect 1342 4027 1366 4098
rect 1437 4062 1700 4098
rect 35836 4098 36478 4118
rect 35836 4062 36085 4098
rect 1437 4027 1460 4062
rect 1046 4008 1460 4027
rect 36064 4027 36085 4062
rect 36156 4027 36180 4098
rect 36251 4027 36289 4098
rect 36360 4027 36384 4098
rect 36455 4027 36478 4098
rect 36064 4008 36478 4027
rect 570 3810 984 3830
rect 570 3739 591 3810
rect 662 3739 686 3810
rect 757 3739 795 3810
rect 866 3739 890 3810
rect 961 3776 984 3810
rect 36540 3810 36954 3830
rect 36540 3776 36561 3810
rect 961 3739 1700 3776
rect 570 3720 1700 3739
rect 35836 3739 36561 3776
rect 36632 3739 36656 3810
rect 36727 3739 36765 3810
rect 36836 3739 36860 3810
rect 36931 3739 36954 3810
rect 35836 3720 36954 3739
rect 182 3640 188 3692
rect 244 3664 1700 3692
rect 244 3640 250 3664
rect 41602 3656 42660 3668
rect 37394 3583 37602 3617
rect 37394 3527 37427 3583
rect 37483 3527 37516 3583
rect 37572 3527 37602 3583
rect 37394 3492 37602 3527
rect 0 3434 1700 3462
rect 37394 3436 37427 3492
rect 37483 3436 37516 3492
rect 37572 3436 37602 3492
rect 41602 3494 42410 3656
rect 42648 3494 42660 3656
rect 41602 3484 42660 3494
rect 37394 3401 37602 3436
rect 0 3352 1700 3380
rect 37394 3345 37427 3401
rect 37483 3345 37516 3401
rect 37572 3345 37602 3401
rect 290 3272 296 3324
rect 352 3296 1700 3324
rect 37394 3318 37602 3345
rect 352 3272 358 3296
rect 37042 3237 37364 3252
rect 42396 3250 42660 3276
rect 37042 3199 37061 3237
rect 398 3130 410 3182
rect 524 3170 570 3182
rect 524 3142 1700 3170
rect 35836 3157 37061 3199
rect 37148 3157 37161 3237
rect 37248 3157 37261 3237
rect 37348 3157 37364 3237
rect 35836 3142 37364 3157
rect 37444 3222 37602 3237
rect 37444 3170 37451 3222
rect 37503 3170 37542 3222
rect 37594 3170 37602 3222
rect 524 3130 570 3142
rect 37444 3120 37602 3170
rect 1046 3092 1700 3114
rect 1046 3021 1067 3092
rect 1138 3021 1162 3092
rect 1233 3021 1271 3092
rect 1342 3021 1366 3092
rect 1437 3058 1700 3092
rect 35836 3094 36478 3114
rect 35836 3058 36085 3094
rect 1437 3021 1460 3058
rect 1046 3002 1460 3021
rect 36064 3023 36085 3058
rect 36156 3023 36180 3094
rect 36251 3023 36289 3094
rect 36360 3023 36384 3094
rect 36455 3023 36478 3094
rect 36064 3004 36478 3023
rect 37444 3068 37451 3120
rect 37503 3068 37542 3120
rect 37594 3068 37602 3120
rect 37444 3017 37602 3068
rect 37444 2965 37452 3017
rect 37504 2965 37543 3017
rect 37595 2965 37602 3017
rect 37444 2924 37602 2965
rect 37444 2872 37452 2924
rect 37504 2872 37543 2924
rect 37595 2872 37602 2924
rect 37444 2859 37602 2872
rect 42396 2838 42422 3250
rect 42634 2838 42660 3250
rect 570 2806 984 2826
rect 570 2735 591 2806
rect 662 2735 686 2806
rect 757 2735 795 2806
rect 866 2735 890 2806
rect 961 2772 984 2806
rect 36540 2806 36954 2826
rect 42396 2814 42660 2838
rect 36540 2772 36561 2806
rect 961 2735 1700 2772
rect 570 2716 1700 2735
rect 35836 2735 36561 2772
rect 36632 2735 36656 2806
rect 36727 2735 36765 2806
rect 36836 2735 36860 2806
rect 36931 2735 36954 2806
rect 35836 2716 36954 2735
rect 41602 2788 42164 2806
rect 182 2636 188 2688
rect 244 2660 1700 2688
rect 244 2636 250 2660
rect 41602 2638 41930 2788
rect 42142 2638 42164 2788
rect 41602 2624 42164 2638
rect 0 2430 1700 2458
rect 0 2348 1700 2376
rect 290 2268 296 2320
rect 352 2292 1700 2320
rect 352 2268 358 2292
rect 37042 2233 37364 2248
rect 37042 2195 37061 2233
rect 398 2126 410 2178
rect 524 2166 570 2178
rect 524 2138 1700 2166
rect 35836 2153 37061 2195
rect 37148 2153 37161 2233
rect 37248 2153 37261 2233
rect 37348 2153 37364 2233
rect 35836 2138 37364 2153
rect 41602 2246 42164 2264
rect 524 2126 570 2138
rect 1046 2089 1700 2110
rect 1046 2018 1067 2089
rect 1138 2018 1162 2089
rect 1233 2018 1271 2089
rect 1342 2018 1366 2089
rect 1437 2054 1700 2089
rect 35836 2090 36478 2110
rect 35836 2054 36085 2090
rect 1437 2018 1460 2054
rect 1046 1999 1460 2018
rect 36064 2019 36085 2054
rect 36156 2019 36180 2090
rect 36251 2019 36289 2090
rect 36360 2019 36384 2090
rect 36455 2019 36478 2090
rect 41602 2096 41930 2246
rect 42142 2096 42164 2246
rect 41602 2082 42164 2096
rect 36064 2000 36478 2019
rect 36540 1802 36954 1822
rect 36540 1768 36561 1802
rect 570 1748 1700 1768
rect 570 1677 591 1748
rect 662 1677 686 1748
rect 757 1677 795 1748
rect 866 1677 890 1748
rect 961 1712 1700 1748
rect 35836 1731 36561 1768
rect 36632 1731 36656 1802
rect 36727 1731 36765 1802
rect 36836 1731 36860 1802
rect 36931 1731 36954 1802
rect 35836 1712 36954 1731
rect 961 1684 984 1712
rect 41602 1690 42164 1708
rect 961 1677 1700 1684
rect 570 1658 1700 1677
rect 620 1656 1700 1658
rect 620 1628 918 1656
rect 41602 1540 41930 1690
rect 42142 1540 42164 1690
rect 41602 1526 42164 1540
rect 42396 1492 42660 1518
rect 1046 1434 1700 1454
rect 1046 1363 1067 1434
rect 1138 1363 1162 1434
rect 1233 1363 1271 1434
rect 1342 1363 1366 1434
rect 1437 1426 1700 1434
rect 37444 1452 37602 1467
rect 1437 1372 1460 1426
rect 37444 1400 37451 1452
rect 37503 1400 37542 1452
rect 37594 1400 37602 1452
rect 1437 1363 1700 1372
rect 1046 1344 1700 1363
rect 37444 1350 37602 1400
rect 1046 1324 1460 1344
rect 1046 1253 1067 1324
rect 1138 1253 1162 1324
rect 1233 1253 1271 1324
rect 1342 1253 1366 1324
rect 1437 1316 1460 1324
rect 1437 1288 1700 1316
rect 37444 1298 37451 1350
rect 37503 1298 37542 1350
rect 37594 1298 37602 1350
rect 1437 1253 1460 1288
rect 1046 1234 1460 1253
rect 37444 1247 37602 1298
rect 37042 1229 37364 1244
rect 37042 1191 37061 1229
rect 398 1122 410 1174
rect 524 1162 570 1174
rect 524 1134 1700 1162
rect 35836 1149 37061 1191
rect 37148 1149 37161 1229
rect 37248 1149 37261 1229
rect 37348 1149 37364 1229
rect 35836 1134 37364 1149
rect 37444 1195 37452 1247
rect 37504 1195 37543 1247
rect 37595 1195 37602 1247
rect 37444 1154 37602 1195
rect 524 1122 570 1134
rect 1046 1085 1700 1106
rect 1046 1014 1067 1085
rect 1138 1014 1162 1085
rect 1233 1014 1271 1085
rect 1342 1014 1366 1085
rect 1437 1050 1700 1085
rect 35836 1086 36478 1106
rect 37444 1102 37452 1154
rect 37504 1102 37543 1154
rect 37595 1102 37602 1154
rect 37444 1089 37602 1102
rect 35836 1050 36085 1086
rect 1437 1014 1460 1050
rect 1046 995 1460 1014
rect 36064 1015 36085 1050
rect 36156 1015 36180 1086
rect 36251 1015 36289 1086
rect 36360 1015 36384 1086
rect 36455 1015 36478 1086
rect 42396 1080 42422 1492
rect 42634 1080 42660 1492
rect 42396 1056 42660 1080
rect 36064 996 36478 1015
rect 2554 893 2670 914
rect 2554 859 2565 893
rect 2662 859 2670 893
rect 2554 832 2670 859
rect 3558 909 3674 914
rect 3558 857 3569 909
rect 3666 857 3674 909
rect 3558 845 3674 857
rect 4194 911 4310 914
rect 4194 859 4205 911
rect 4302 859 4310 911
rect 4194 847 4310 859
rect 4562 910 4678 914
rect 4562 858 4573 910
rect 4670 858 4678 910
rect 4562 846 4678 858
rect 5566 910 5682 914
rect 5566 858 5577 910
rect 5674 858 5682 910
rect 5566 846 5682 858
rect 6570 910 6686 914
rect 6570 858 6581 910
rect 6678 858 6686 910
rect 6570 846 6686 858
rect 7574 910 7690 914
rect 7574 858 7585 910
rect 7682 858 7690 910
rect 7574 846 7690 858
rect 8578 910 8694 914
rect 8578 858 8589 910
rect 8686 858 8694 910
rect 8578 846 8694 858
rect 9582 910 9698 914
rect 9582 858 9593 910
rect 9690 858 9698 910
rect 9582 846 9698 858
rect 10586 910 10702 914
rect 10586 858 10597 910
rect 10694 858 10702 910
rect 10586 846 10702 858
rect 11590 910 11706 914
rect 11590 858 11601 910
rect 11698 858 11706 910
rect 11590 846 11706 858
rect 12594 910 12710 914
rect 12594 858 12605 910
rect 12702 858 12710 910
rect 12594 846 12710 858
rect 13598 910 13714 914
rect 13598 858 13609 910
rect 13706 858 13714 910
rect 13598 846 13714 858
rect 14602 910 14718 914
rect 14602 858 14613 910
rect 14710 858 14718 910
rect 14602 846 14718 858
rect 15606 910 15722 914
rect 15606 858 15617 910
rect 15714 858 15722 910
rect 15606 846 15722 858
rect 16610 910 16726 914
rect 16610 858 16621 910
rect 16718 858 16726 910
rect 16610 846 16726 858
rect 17614 910 17730 914
rect 17614 858 17625 910
rect 17722 858 17730 910
rect 17614 846 17730 858
rect 18244 911 18360 914
rect 18244 859 18255 911
rect 18352 859 18360 911
rect 18244 847 18360 859
rect 18618 910 18734 914
rect 18618 858 18629 910
rect 18726 858 18734 910
rect 18618 846 18734 858
rect 19250 911 19366 914
rect 19250 859 19261 911
rect 19358 859 19366 911
rect 19250 847 19366 859
rect 19622 910 19738 914
rect 19622 858 19633 910
rect 19730 858 19738 910
rect 19622 846 19738 858
rect 20246 911 20362 914
rect 20246 859 20257 911
rect 20354 859 20362 911
rect 20246 847 20362 859
rect 20626 910 20742 914
rect 20626 858 20637 910
rect 20734 858 20742 910
rect 20626 846 20742 858
rect 21630 910 21746 914
rect 21630 858 21641 910
rect 21738 858 21746 910
rect 21630 846 21746 858
rect 22634 910 22750 914
rect 22634 858 22645 910
rect 22742 858 22750 910
rect 22634 846 22750 858
rect 23638 910 23754 914
rect 23638 858 23649 910
rect 23746 858 23754 910
rect 23638 846 23754 858
rect 24642 910 24758 914
rect 24642 858 24653 910
rect 24750 858 24758 910
rect 24642 846 24758 858
rect 25646 910 25762 914
rect 25646 858 25657 910
rect 25754 858 25762 910
rect 25646 846 25762 858
rect 26650 910 26766 914
rect 26650 858 26661 910
rect 26758 858 26766 910
rect 26650 846 26766 858
rect 27654 910 27770 914
rect 27654 858 27665 910
rect 27762 858 27770 910
rect 27654 846 27770 858
rect 28658 892 28774 914
rect 28658 858 28669 892
rect 28766 858 28774 892
rect 28658 846 28774 858
rect 29662 910 29778 914
rect 29662 858 29673 910
rect 29770 858 29778 910
rect 29662 846 29778 858
rect 30666 910 30782 914
rect 30666 858 30677 910
rect 30774 858 30782 910
rect 30666 846 30782 858
rect 31670 910 31786 914
rect 31670 858 31681 910
rect 31778 858 31786 910
rect 31670 846 31786 858
rect 32674 910 32790 914
rect 32674 858 32685 910
rect 32782 858 32790 910
rect 32674 846 32790 858
rect 33600 910 33716 914
rect 33600 858 33611 910
rect 33708 858 33716 910
rect 34105 908 34145 914
rect 34682 910 34798 914
rect 33600 846 33716 858
rect 34083 907 34147 908
rect 34083 855 34089 907
rect 34141 855 34147 907
rect 34083 854 34147 855
rect 34682 858 34693 910
rect 34790 858 34798 910
rect 34682 846 34798 858
rect 37394 875 37602 909
rect 570 812 2670 832
rect 570 741 591 812
rect 662 741 686 812
rect 757 741 795 812
rect 866 741 890 812
rect 961 790 2670 812
rect 27848 801 28774 846
rect 37394 819 37427 875
rect 37483 819 37516 875
rect 37572 819 37602 875
rect 27848 795 27912 801
rect 961 772 984 790
rect 961 741 983 772
rect 27848 743 27854 795
rect 27906 743 27912 795
rect 27848 742 27912 743
rect 37394 784 37602 819
rect 570 722 983 741
rect 29672 739 29736 740
rect 29672 734 29678 739
rect 28052 719 29678 734
rect 28052 667 28058 719
rect 28110 687 29678 719
rect 29730 687 29736 739
rect 28110 686 29736 687
rect 37394 728 37427 784
rect 37483 728 37516 784
rect 37572 728 37602 784
rect 37394 693 37602 728
rect 28110 667 28116 686
rect 28052 666 28116 667
rect 30690 651 30754 652
rect 28251 649 28315 650
rect 28251 597 28257 649
rect 28309 648 28315 649
rect 30690 648 30696 651
rect 28309 600 30696 648
rect 28309 597 28315 600
rect 30690 599 30696 600
rect 30748 599 30754 651
rect 37394 637 37427 693
rect 37483 637 37516 693
rect 37572 637 37602 693
rect 37394 610 37602 637
rect 30690 598 30754 599
rect 28251 596 28315 597
rect 31696 575 31760 576
rect 28455 570 28519 571
rect 31696 570 31702 575
rect 28455 518 28461 570
rect 28513 523 31702 570
rect 31754 523 31760 575
rect 41847 557 42660 558
rect 41602 546 42660 557
rect 28513 522 31760 523
rect 36540 526 36954 546
rect 28513 518 28519 522
rect 28455 517 28519 518
rect 32700 499 32764 500
rect 32700 494 32706 499
rect 28659 493 32706 494
rect 28659 441 28665 493
rect 28717 447 32706 493
rect 32758 447 32764 499
rect 36540 493 36561 526
rect 28717 446 32764 447
rect 35678 487 36561 493
rect 35678 453 35690 487
rect 35724 455 36561 487
rect 36632 455 36656 526
rect 36727 455 36765 526
rect 36836 455 36860 526
rect 36931 455 36954 526
rect 35724 453 36954 455
rect 28717 441 28723 446
rect 35678 445 36954 453
rect 28659 440 28723 441
rect 36540 436 36954 445
rect 33628 423 33692 424
rect 33628 418 33634 423
rect 28863 417 33634 418
rect 28863 365 28869 417
rect 28921 371 33634 417
rect 33686 371 33692 423
rect 41602 384 42410 546
rect 42648 384 42660 546
rect 41602 374 42660 384
rect 41602 373 41847 374
rect 28921 370 33692 371
rect 28921 365 28927 370
rect 28863 364 28927 365
rect 34680 347 34744 348
rect 34680 342 34686 347
rect 29067 341 34686 342
rect 29067 289 29073 341
rect 29125 295 34686 341
rect 34738 295 34744 347
rect 29125 294 34744 295
rect 29125 289 29131 294
rect 29067 288 29131 289
rect 34082 120 42810 124
rect 34082 68 34088 120
rect 34141 68 42810 120
rect 34082 56 42810 68
rect 34082 4 34088 56
rect 34141 8 42810 56
rect 34141 4 34147 8
rect 34082 3 34147 4
<< via1 >>
rect 42410 23494 42648 23656
rect 42422 22838 42634 23250
rect 41930 22638 42142 22788
rect 41930 22096 42142 22246
rect 41930 21540 42142 21690
rect 42422 21080 42634 21492
rect 42410 20384 42648 20546
rect 1898 19946 2160 20104
rect 5026 19946 5288 20104
rect 5898 19946 6160 20104
rect 9026 19946 9288 20104
rect 9898 19946 10160 20104
rect 13026 19946 13288 20104
rect 13898 19946 14160 20104
rect 17026 19946 17288 20104
rect 17898 19946 18160 20104
rect 21026 19946 21288 20104
rect 21898 19946 22160 20104
rect 25026 19946 25288 20104
rect 25898 19946 26160 20104
rect 29026 19946 29288 20104
rect 29898 19946 30160 20104
rect 33026 19946 33288 20104
rect 33898 19946 34160 20104
rect 37026 19980 37288 20104
rect 587 19634 969 19889
rect 3444 19638 3770 19882
rect 7444 19638 7770 19882
rect 11444 19638 11770 19882
rect 15444 19638 15770 19882
rect 19444 19638 19770 19882
rect 23444 19638 23770 19882
rect 27444 19638 27770 19882
rect 31444 19638 31770 19882
rect 35426 19783 35490 19847
rect 35522 19783 35586 19847
rect 35618 19783 35682 19847
rect 35714 19783 35778 19847
rect 36570 19821 36634 19885
rect 36666 19821 36730 19885
rect 36762 19821 36826 19885
rect 36858 19821 36922 19885
rect 35426 19689 35490 19753
rect 35522 19689 35586 19753
rect 35618 19689 35682 19753
rect 35714 19689 35778 19753
rect 36570 19727 36634 19791
rect 36666 19727 36730 19791
rect 36762 19727 36826 19791
rect 36858 19727 36922 19791
rect 37427 19495 37483 19551
rect 37516 19495 37572 19551
rect 1063 19196 1445 19451
rect 1904 19386 1960 19442
rect 1998 19386 2054 19442
rect 2092 19386 2148 19442
rect 5032 19386 5088 19442
rect 5126 19386 5182 19442
rect 5220 19386 5276 19442
rect 5904 19386 5960 19442
rect 5998 19386 6054 19442
rect 6092 19386 6148 19442
rect 9032 19386 9088 19442
rect 9126 19386 9182 19442
rect 9220 19386 9276 19442
rect 9904 19386 9960 19442
rect 9998 19386 10054 19442
rect 10092 19386 10148 19442
rect 13032 19386 13088 19442
rect 13126 19386 13182 19442
rect 13220 19386 13276 19442
rect 13904 19386 13960 19442
rect 13998 19386 14054 19442
rect 14092 19386 14148 19442
rect 17032 19386 17088 19442
rect 17126 19386 17182 19442
rect 17220 19386 17276 19442
rect 17904 19386 17960 19442
rect 17998 19386 18054 19442
rect 18092 19386 18148 19442
rect 21032 19386 21088 19442
rect 21126 19386 21182 19442
rect 21220 19386 21276 19442
rect 21904 19386 21960 19442
rect 21998 19386 22054 19442
rect 22092 19386 22148 19442
rect 25032 19386 25088 19442
rect 25126 19386 25182 19442
rect 25220 19386 25276 19442
rect 25904 19386 25960 19442
rect 25998 19386 26054 19442
rect 26092 19386 26148 19442
rect 29032 19386 29088 19442
rect 29126 19386 29182 19442
rect 29220 19386 29276 19442
rect 29904 19386 29960 19442
rect 29998 19386 30054 19442
rect 30092 19386 30148 19442
rect 33032 19386 33088 19442
rect 33126 19386 33182 19442
rect 33220 19386 33276 19442
rect 33904 19386 33960 19442
rect 33998 19386 34054 19442
rect 34092 19386 34148 19442
rect 1904 19292 1960 19348
rect 1998 19292 2054 19348
rect 2092 19292 2148 19348
rect 5032 19292 5088 19348
rect 5126 19292 5182 19348
rect 5220 19292 5276 19348
rect 5904 19292 5960 19348
rect 5998 19292 6054 19348
rect 6092 19292 6148 19348
rect 9032 19292 9088 19348
rect 9126 19292 9182 19348
rect 9220 19292 9276 19348
rect 9904 19292 9960 19348
rect 9998 19292 10054 19348
rect 10092 19292 10148 19348
rect 13032 19292 13088 19348
rect 13126 19292 13182 19348
rect 13220 19292 13276 19348
rect 13904 19292 13960 19348
rect 13998 19292 14054 19348
rect 14092 19292 14148 19348
rect 17032 19292 17088 19348
rect 17126 19292 17182 19348
rect 17220 19292 17276 19348
rect 17904 19292 17960 19348
rect 17998 19292 18054 19348
rect 18092 19292 18148 19348
rect 21032 19292 21088 19348
rect 21126 19292 21182 19348
rect 21220 19292 21276 19348
rect 21904 19292 21960 19348
rect 21998 19292 22054 19348
rect 22092 19292 22148 19348
rect 25032 19292 25088 19348
rect 25126 19292 25182 19348
rect 25220 19292 25276 19348
rect 25904 19292 25960 19348
rect 25998 19292 26054 19348
rect 26092 19292 26148 19348
rect 29032 19292 29088 19348
rect 29126 19292 29182 19348
rect 29220 19292 29276 19348
rect 29904 19292 29960 19348
rect 29998 19292 30054 19348
rect 30092 19292 30148 19348
rect 33032 19292 33088 19348
rect 33126 19292 33182 19348
rect 33220 19292 33276 19348
rect 33904 19292 33960 19348
rect 33998 19292 34054 19348
rect 34092 19292 34148 19348
rect 36094 19311 36158 19375
rect 36190 19311 36254 19375
rect 36286 19311 36350 19375
rect 36382 19311 36446 19375
rect 42410 19494 42648 19656
rect 37427 19404 37483 19460
rect 37516 19404 37572 19460
rect 37427 19313 37483 19369
rect 37516 19313 37572 19369
rect 1904 19198 1960 19254
rect 1998 19198 2054 19254
rect 2092 19198 2148 19254
rect 5032 19198 5088 19254
rect 5126 19198 5182 19254
rect 5220 19198 5276 19254
rect 5904 19198 5960 19254
rect 5998 19198 6054 19254
rect 6092 19198 6148 19254
rect 9032 19198 9088 19254
rect 9126 19198 9182 19254
rect 9220 19198 9276 19254
rect 9904 19198 9960 19254
rect 9998 19198 10054 19254
rect 10092 19198 10148 19254
rect 13032 19198 13088 19254
rect 13126 19198 13182 19254
rect 13220 19198 13276 19254
rect 13904 19198 13960 19254
rect 13998 19198 14054 19254
rect 14092 19198 14148 19254
rect 17032 19198 17088 19254
rect 17126 19198 17182 19254
rect 17220 19198 17276 19254
rect 17904 19198 17960 19254
rect 17998 19198 18054 19254
rect 18092 19198 18148 19254
rect 21032 19198 21088 19254
rect 21126 19198 21182 19254
rect 21220 19198 21276 19254
rect 21904 19198 21960 19254
rect 21998 19198 22054 19254
rect 22092 19198 22148 19254
rect 25032 19198 25088 19254
rect 25126 19198 25182 19254
rect 25220 19198 25276 19254
rect 25904 19198 25960 19254
rect 25998 19198 26054 19254
rect 26092 19198 26148 19254
rect 29032 19198 29088 19254
rect 29126 19198 29182 19254
rect 29220 19198 29276 19254
rect 29904 19198 29960 19254
rect 29998 19198 30054 19254
rect 30092 19198 30148 19254
rect 33032 19198 33088 19254
rect 33126 19198 33182 19254
rect 33220 19198 33276 19254
rect 33904 19198 33960 19254
rect 33998 19198 34054 19254
rect 34092 19198 34148 19254
rect 36094 19217 36158 19281
rect 36190 19217 36254 19281
rect 36286 19217 36350 19281
rect 36382 19217 36446 19281
rect 37451 19160 37503 19212
rect 37542 19160 37594 19212
rect 37451 19058 37503 19110
rect 37542 19058 37594 19110
rect 37452 18955 37504 19007
rect 37543 18955 37595 19007
rect 591 18745 662 18816
rect 686 18745 757 18816
rect 795 18745 866 18816
rect 890 18745 961 18816
rect 36561 18799 36632 18870
rect 36656 18799 36727 18870
rect 36765 18799 36836 18870
rect 36860 18799 36931 18870
rect 37452 18862 37504 18914
rect 37543 18862 37595 18914
rect 42422 18838 42634 19250
rect 41930 18638 42142 18788
rect 591 18431 662 18502
rect 686 18431 757 18502
rect 795 18431 866 18502
rect 890 18431 961 18502
rect 1067 18292 1138 18363
rect 1162 18292 1233 18363
rect 1271 18292 1342 18363
rect 1366 18292 1437 18363
rect 404 18190 460 18242
rect 472 18190 528 18242
rect 37061 18217 37148 18297
rect 37161 18217 37248 18297
rect 37261 18217 37348 18297
rect 1067 18082 1138 18153
rect 1162 18082 1233 18153
rect 1271 18082 1342 18153
rect 1366 18082 1437 18153
rect 36085 18083 36156 18154
rect 36180 18083 36251 18154
rect 36289 18083 36360 18154
rect 36384 18083 36455 18154
rect 41930 18096 42142 18246
rect 591 17795 662 17866
rect 686 17795 757 17866
rect 795 17795 866 17866
rect 890 17795 961 17866
rect 36561 17795 36632 17866
rect 36656 17795 36727 17866
rect 36765 17795 36836 17866
rect 36860 17795 36931 17866
rect 188 17696 244 17748
rect 41930 17540 42142 17690
rect 37451 17400 37503 17452
rect 37542 17400 37594 17452
rect 296 17328 352 17380
rect 410 17186 524 17238
rect 37061 17213 37148 17293
rect 37161 17213 37248 17293
rect 37261 17213 37348 17293
rect 37451 17298 37503 17350
rect 37542 17298 37594 17350
rect 37452 17195 37504 17247
rect 37543 17195 37595 17247
rect 1067 17079 1138 17150
rect 1162 17079 1233 17150
rect 1271 17079 1342 17150
rect 1366 17079 1437 17150
rect 36085 17079 36156 17150
rect 36180 17079 36251 17150
rect 36289 17079 36360 17150
rect 36384 17079 36455 17150
rect 37452 17102 37504 17154
rect 37543 17102 37595 17154
rect 42422 17080 42634 17492
rect 591 16791 662 16862
rect 686 16791 757 16862
rect 795 16791 866 16862
rect 890 16791 961 16862
rect 36561 16791 36632 16862
rect 36656 16791 36727 16862
rect 36765 16791 36836 16862
rect 36860 16791 36931 16862
rect 188 16692 244 16744
rect 37427 16590 37483 16646
rect 37516 16590 37572 16646
rect 37427 16499 37483 16555
rect 37516 16499 37572 16555
rect 37427 16408 37483 16464
rect 37516 16408 37572 16464
rect 42410 16384 42648 16546
rect 296 16324 352 16376
rect 410 16182 524 16234
rect 37061 16209 37148 16289
rect 37161 16209 37248 16289
rect 37261 16209 37348 16289
rect 1067 16074 1138 16145
rect 1162 16074 1233 16145
rect 1271 16074 1342 16145
rect 1366 16074 1437 16145
rect 36085 16075 36156 16146
rect 36180 16075 36251 16146
rect 36289 16075 36360 16146
rect 36384 16075 36455 16146
rect 591 15787 662 15858
rect 686 15787 757 15858
rect 795 15787 866 15858
rect 890 15787 961 15858
rect 36561 15787 36632 15858
rect 36656 15787 36727 15858
rect 36765 15787 36836 15858
rect 36860 15787 36931 15858
rect 188 15688 244 15740
rect 42410 15494 42648 15656
rect 296 15320 352 15372
rect 410 15178 524 15230
rect 37061 15205 37148 15285
rect 37161 15205 37248 15285
rect 37261 15205 37348 15285
rect 1067 15071 1138 15142
rect 1162 15071 1233 15142
rect 1271 15071 1342 15142
rect 1366 15071 1437 15142
rect 36085 15071 36156 15142
rect 36180 15071 36251 15142
rect 36289 15071 36360 15142
rect 36384 15071 36455 15142
rect 37451 15160 37503 15212
rect 37542 15160 37594 15212
rect 37451 15058 37503 15110
rect 37542 15058 37594 15110
rect 37452 14955 37504 15007
rect 37543 14955 37595 15007
rect 591 14783 662 14854
rect 686 14783 757 14854
rect 795 14783 866 14854
rect 890 14783 961 14854
rect 36561 14783 36632 14854
rect 36656 14783 36727 14854
rect 36765 14783 36836 14854
rect 36860 14783 36931 14854
rect 37452 14862 37504 14914
rect 37543 14862 37595 14914
rect 42422 14838 42634 15250
rect 188 14684 244 14736
rect 41930 14638 42142 14788
rect 296 14316 352 14368
rect 410 14174 524 14226
rect 37061 14201 37148 14281
rect 37161 14201 37248 14281
rect 37261 14201 37348 14281
rect 1067 14067 1138 14138
rect 1162 14067 1233 14138
rect 1271 14067 1342 14138
rect 1366 14067 1437 14138
rect 36085 14067 36156 14138
rect 36180 14067 36251 14138
rect 36289 14067 36360 14138
rect 36384 14067 36455 14138
rect 41930 14096 42142 14246
rect 591 13779 662 13850
rect 686 13779 757 13850
rect 795 13779 866 13850
rect 890 13779 961 13850
rect 36561 13779 36632 13850
rect 36656 13779 36727 13850
rect 36765 13779 36836 13850
rect 36860 13779 36931 13850
rect 188 13680 244 13732
rect 41930 13540 42142 13690
rect 37451 13400 37503 13452
rect 37542 13400 37594 13452
rect 296 13312 352 13364
rect 37451 13298 37503 13350
rect 37542 13298 37594 13350
rect 410 13170 524 13222
rect 37061 13197 37148 13277
rect 37161 13197 37248 13277
rect 37261 13197 37348 13277
rect 37452 13195 37504 13247
rect 37543 13195 37595 13247
rect 1067 13063 1138 13134
rect 1162 13063 1233 13134
rect 1271 13063 1342 13134
rect 1366 13063 1437 13134
rect 36085 13063 36156 13134
rect 36180 13063 36251 13134
rect 36289 13063 36360 13134
rect 36384 13063 36455 13134
rect 37452 13102 37504 13154
rect 37543 13102 37595 13154
rect 42422 13080 42634 13492
rect 591 12775 662 12846
rect 686 12775 757 12846
rect 795 12775 866 12846
rect 890 12775 961 12846
rect 36561 12775 36632 12846
rect 36656 12775 36727 12846
rect 36765 12775 36836 12846
rect 36860 12775 36931 12846
rect 188 12676 244 12728
rect 37427 12532 37483 12588
rect 37516 12532 37572 12588
rect 37427 12441 37483 12497
rect 37516 12441 37572 12497
rect 296 12308 352 12360
rect 37427 12350 37483 12406
rect 37516 12350 37572 12406
rect 42410 12384 42648 12546
rect 410 12166 524 12218
rect 37061 12193 37148 12273
rect 37161 12193 37248 12273
rect 37261 12193 37348 12273
rect 1067 12059 1138 12130
rect 1162 12059 1233 12130
rect 1271 12059 1342 12130
rect 1366 12059 1437 12130
rect 36085 12059 36156 12130
rect 36180 12059 36251 12130
rect 36289 12059 36360 12130
rect 36384 12059 36455 12130
rect 591 11771 662 11842
rect 686 11771 757 11842
rect 795 11771 866 11842
rect 890 11771 961 11842
rect 36561 11771 36632 11842
rect 36656 11771 36727 11842
rect 36765 11771 36836 11842
rect 36860 11771 36931 11842
rect 188 11672 244 11724
rect 42410 11494 42648 11656
rect 296 11304 352 11356
rect 410 11162 524 11214
rect 37061 11189 37148 11269
rect 37161 11189 37248 11269
rect 37261 11189 37348 11269
rect 37451 11160 37503 11212
rect 37542 11160 37594 11212
rect 1067 11055 1138 11126
rect 1162 11055 1233 11126
rect 1271 11055 1342 11126
rect 1366 11055 1437 11126
rect 36085 11055 36156 11126
rect 36180 11055 36251 11126
rect 36289 11055 36360 11126
rect 36384 11055 36455 11126
rect 37451 11058 37503 11110
rect 37542 11058 37594 11110
rect 37452 10955 37504 11007
rect 37543 10955 37595 11007
rect 37452 10862 37504 10914
rect 37543 10862 37595 10914
rect 591 10767 662 10838
rect 686 10767 757 10838
rect 795 10767 866 10838
rect 890 10767 961 10838
rect 36561 10767 36632 10838
rect 36656 10767 36727 10838
rect 36765 10767 36836 10838
rect 36860 10767 36931 10838
rect 42422 10838 42634 11250
rect 188 10668 244 10720
rect 41930 10638 42142 10788
rect 296 10300 352 10352
rect 410 10158 524 10210
rect 37061 10185 37148 10265
rect 37161 10185 37248 10265
rect 37261 10185 37348 10265
rect 1067 10051 1138 10122
rect 1162 10051 1233 10122
rect 1271 10051 1342 10122
rect 1366 10051 1437 10122
rect 36085 10051 36156 10122
rect 36180 10051 36251 10122
rect 36289 10051 36360 10122
rect 36384 10051 36455 10122
rect 41930 10096 42142 10246
rect 591 9763 662 9834
rect 686 9763 757 9834
rect 795 9763 866 9834
rect 890 9763 961 9834
rect 36561 9763 36632 9834
rect 36656 9763 36727 9834
rect 36765 9763 36836 9834
rect 36860 9763 36931 9834
rect 188 9664 244 9716
rect 41930 9540 42142 9690
rect 37451 9400 37503 9452
rect 37542 9400 37594 9452
rect 296 9296 352 9348
rect 37451 9298 37503 9350
rect 37542 9298 37594 9350
rect 410 9154 524 9206
rect 37061 9181 37148 9261
rect 37161 9181 37248 9261
rect 37261 9181 37348 9261
rect 37452 9195 37504 9247
rect 37543 9195 37595 9247
rect 1067 9047 1138 9118
rect 1162 9047 1233 9118
rect 1271 9047 1342 9118
rect 1366 9047 1437 9118
rect 36085 9047 36156 9118
rect 36180 9047 36251 9118
rect 36289 9047 36360 9118
rect 36384 9047 36455 9118
rect 37452 9102 37504 9154
rect 37543 9102 37595 9154
rect 42422 9080 42634 9492
rect 591 8759 662 8830
rect 686 8759 757 8830
rect 795 8759 866 8830
rect 890 8759 961 8830
rect 36561 8759 36632 8830
rect 36656 8759 36727 8830
rect 36765 8759 36836 8830
rect 36860 8759 36931 8830
rect 188 8660 244 8712
rect 37427 8439 37483 8495
rect 37516 8439 37572 8495
rect 37427 8348 37483 8404
rect 37516 8348 37572 8404
rect 42410 8384 42648 8546
rect 296 8292 352 8344
rect 410 8150 524 8202
rect 37061 8177 37148 8257
rect 37161 8177 37248 8257
rect 37261 8177 37348 8257
rect 37427 8257 37483 8313
rect 37516 8257 37572 8313
rect 1067 8043 1138 8114
rect 1162 8043 1233 8114
rect 1271 8043 1342 8114
rect 1366 8043 1437 8114
rect 36085 8043 36156 8114
rect 36180 8043 36251 8114
rect 36289 8043 36360 8114
rect 36384 8043 36455 8114
rect 591 7755 662 7826
rect 686 7755 757 7826
rect 795 7755 866 7826
rect 890 7755 961 7826
rect 36561 7755 36632 7826
rect 36656 7755 36727 7826
rect 36765 7755 36836 7826
rect 36860 7755 36931 7826
rect 188 7656 244 7708
rect 42410 7494 42648 7656
rect 296 7288 352 7340
rect 410 7146 524 7198
rect 37061 7173 37148 7253
rect 37161 7173 37248 7253
rect 37261 7173 37348 7253
rect 37451 7160 37503 7212
rect 37542 7160 37594 7212
rect 1067 7039 1138 7110
rect 1162 7039 1233 7110
rect 1271 7039 1342 7110
rect 1366 7039 1437 7110
rect 36085 7039 36156 7110
rect 36180 7039 36251 7110
rect 36289 7039 36360 7110
rect 36384 7039 36455 7110
rect 37451 7058 37503 7110
rect 37542 7058 37594 7110
rect 37452 6955 37504 7007
rect 37543 6955 37595 7007
rect 37452 6862 37504 6914
rect 37543 6862 37595 6914
rect 591 6751 662 6822
rect 686 6751 757 6822
rect 795 6751 866 6822
rect 890 6751 961 6822
rect 36561 6751 36632 6822
rect 36656 6751 36727 6822
rect 36765 6751 36836 6822
rect 36860 6751 36931 6822
rect 42422 6838 42634 7250
rect 188 6652 244 6704
rect 41930 6638 42142 6788
rect 296 6284 352 6336
rect 410 6142 524 6194
rect 37061 6169 37148 6249
rect 37161 6169 37248 6249
rect 37261 6169 37348 6249
rect 1067 6035 1138 6106
rect 1162 6035 1233 6106
rect 1271 6035 1342 6106
rect 1366 6035 1437 6106
rect 36085 6035 36156 6106
rect 36180 6035 36251 6106
rect 36289 6035 36360 6106
rect 36384 6035 36455 6106
rect 41930 6096 42142 6246
rect 591 5747 662 5818
rect 686 5747 757 5818
rect 795 5747 866 5818
rect 890 5747 961 5818
rect 36561 5747 36632 5818
rect 36656 5747 36727 5818
rect 36765 5747 36836 5818
rect 36860 5747 36931 5818
rect 188 5648 244 5700
rect 41930 5540 42142 5690
rect 37451 5400 37503 5452
rect 37542 5400 37594 5452
rect 296 5280 352 5332
rect 37451 5298 37503 5350
rect 37542 5298 37594 5350
rect 410 5138 524 5190
rect 37061 5165 37148 5245
rect 37161 5165 37248 5245
rect 37261 5165 37348 5245
rect 37452 5195 37504 5247
rect 37543 5195 37595 5247
rect 1067 5031 1138 5102
rect 1162 5031 1233 5102
rect 1271 5031 1342 5102
rect 1366 5031 1437 5102
rect 36085 5031 36156 5102
rect 36180 5031 36251 5102
rect 36289 5031 36360 5102
rect 36384 5031 36455 5102
rect 37452 5102 37504 5154
rect 37543 5102 37595 5154
rect 42422 5080 42634 5492
rect 591 4743 662 4814
rect 686 4743 757 4814
rect 795 4743 866 4814
rect 890 4743 961 4814
rect 36561 4743 36632 4814
rect 36656 4743 36727 4814
rect 36765 4743 36836 4814
rect 36860 4743 36931 4814
rect 188 4644 244 4696
rect 42410 4384 42648 4546
rect 296 4276 352 4328
rect 410 4134 524 4186
rect 37061 4161 37148 4241
rect 37161 4161 37248 4241
rect 37261 4161 37348 4241
rect 1067 4027 1138 4098
rect 1162 4027 1233 4098
rect 1271 4027 1342 4098
rect 1366 4027 1437 4098
rect 36085 4027 36156 4098
rect 36180 4027 36251 4098
rect 36289 4027 36360 4098
rect 36384 4027 36455 4098
rect 591 3739 662 3810
rect 686 3739 757 3810
rect 795 3739 866 3810
rect 890 3739 961 3810
rect 36561 3739 36632 3810
rect 36656 3739 36727 3810
rect 36765 3739 36836 3810
rect 36860 3739 36931 3810
rect 188 3640 244 3692
rect 37427 3527 37483 3583
rect 37516 3527 37572 3583
rect 37427 3436 37483 3492
rect 37516 3436 37572 3492
rect 42410 3494 42648 3656
rect 37427 3345 37483 3401
rect 37516 3345 37572 3401
rect 296 3272 352 3324
rect 410 3130 524 3182
rect 37061 3157 37148 3237
rect 37161 3157 37248 3237
rect 37261 3157 37348 3237
rect 37451 3170 37503 3222
rect 37542 3170 37594 3222
rect 1067 3021 1138 3092
rect 1162 3021 1233 3092
rect 1271 3021 1342 3092
rect 1366 3021 1437 3092
rect 36085 3023 36156 3094
rect 36180 3023 36251 3094
rect 36289 3023 36360 3094
rect 36384 3023 36455 3094
rect 37451 3068 37503 3120
rect 37542 3068 37594 3120
rect 37452 2965 37504 3017
rect 37543 2965 37595 3017
rect 37452 2872 37504 2924
rect 37543 2872 37595 2924
rect 42422 2838 42634 3250
rect 591 2735 662 2806
rect 686 2735 757 2806
rect 795 2735 866 2806
rect 890 2735 961 2806
rect 36561 2735 36632 2806
rect 36656 2735 36727 2806
rect 36765 2735 36836 2806
rect 36860 2735 36931 2806
rect 188 2636 244 2688
rect 41930 2638 42142 2788
rect 296 2268 352 2320
rect 410 2126 524 2178
rect 37061 2153 37148 2233
rect 37161 2153 37248 2233
rect 37261 2153 37348 2233
rect 1067 2018 1138 2089
rect 1162 2018 1233 2089
rect 1271 2018 1342 2089
rect 1366 2018 1437 2089
rect 36085 2019 36156 2090
rect 36180 2019 36251 2090
rect 36289 2019 36360 2090
rect 36384 2019 36455 2090
rect 41930 2096 42142 2246
rect 591 1677 662 1748
rect 686 1677 757 1748
rect 795 1677 866 1748
rect 890 1677 961 1748
rect 36561 1731 36632 1802
rect 36656 1731 36727 1802
rect 36765 1731 36836 1802
rect 36860 1731 36931 1802
rect 41930 1540 42142 1690
rect 1067 1363 1138 1434
rect 1162 1363 1233 1434
rect 1271 1363 1342 1434
rect 1366 1363 1437 1434
rect 37451 1400 37503 1452
rect 37542 1400 37594 1452
rect 1067 1253 1138 1324
rect 1162 1253 1233 1324
rect 1271 1253 1342 1324
rect 1366 1253 1437 1324
rect 37451 1298 37503 1350
rect 37542 1298 37594 1350
rect 410 1122 524 1174
rect 37061 1149 37148 1229
rect 37161 1149 37248 1229
rect 37261 1149 37348 1229
rect 37452 1195 37504 1247
rect 37543 1195 37595 1247
rect 1067 1014 1138 1085
rect 1162 1014 1233 1085
rect 1271 1014 1342 1085
rect 1366 1014 1437 1085
rect 37452 1102 37504 1154
rect 37543 1102 37595 1154
rect 36085 1015 36156 1086
rect 36180 1015 36251 1086
rect 36289 1015 36360 1086
rect 36384 1015 36455 1086
rect 42422 1080 42634 1492
rect 3569 891 3666 909
rect 3569 857 3666 891
rect 4205 893 4302 911
rect 4205 859 4302 893
rect 4573 892 4670 910
rect 4573 858 4670 892
rect 5577 892 5674 910
rect 5577 858 5674 892
rect 6581 892 6678 910
rect 6581 858 6678 892
rect 7585 892 7682 910
rect 7585 858 7682 892
rect 8589 892 8686 910
rect 8589 858 8686 892
rect 9593 892 9690 910
rect 9593 858 9690 892
rect 10597 892 10694 910
rect 10597 858 10694 892
rect 11601 892 11698 910
rect 11601 858 11698 892
rect 12605 892 12702 910
rect 12605 858 12702 892
rect 13609 892 13706 910
rect 13609 858 13706 892
rect 14613 892 14710 910
rect 14613 858 14710 892
rect 15617 892 15714 910
rect 15617 858 15714 892
rect 16621 892 16718 910
rect 16621 858 16718 892
rect 17625 892 17722 910
rect 17625 858 17722 892
rect 18255 893 18352 911
rect 18255 859 18352 893
rect 18629 892 18726 910
rect 18629 858 18726 892
rect 19261 893 19358 911
rect 19261 859 19358 893
rect 19633 892 19730 910
rect 19633 858 19730 892
rect 20257 893 20354 911
rect 20257 859 20354 893
rect 20637 892 20734 910
rect 20637 858 20734 892
rect 21641 892 21738 910
rect 21641 858 21738 892
rect 22645 892 22742 910
rect 22645 858 22742 892
rect 23649 892 23746 910
rect 23649 858 23746 892
rect 24653 892 24750 910
rect 24653 858 24750 892
rect 25657 892 25754 910
rect 25657 858 25754 892
rect 26661 892 26758 910
rect 26661 858 26758 892
rect 27665 892 27762 910
rect 27665 858 27762 892
rect 29673 892 29770 910
rect 29673 858 29770 892
rect 30677 893 30774 910
rect 30677 858 30774 893
rect 31681 893 31778 910
rect 31681 858 31778 893
rect 32685 893 32782 910
rect 32685 858 32782 893
rect 33611 893 33708 910
rect 33611 858 33708 893
rect 34089 855 34141 907
rect 34693 893 34790 910
rect 34693 858 34790 893
rect 591 741 662 812
rect 686 741 757 812
rect 795 741 866 812
rect 890 741 961 812
rect 37427 819 37483 875
rect 37516 819 37572 875
rect 27854 743 27906 795
rect 28058 667 28110 719
rect 29678 687 29730 739
rect 37427 728 37483 784
rect 37516 728 37572 784
rect 28257 597 28309 649
rect 30696 599 30748 651
rect 37427 637 37483 693
rect 37516 637 37572 693
rect 28461 518 28513 570
rect 31702 523 31754 575
rect 28665 441 28717 493
rect 32706 447 32758 499
rect 36561 455 36632 526
rect 36656 455 36727 526
rect 36765 455 36836 526
rect 36860 455 36931 526
rect 28869 365 28921 417
rect 33634 371 33686 423
rect 42410 384 42648 546
rect 29073 289 29125 341
rect 34686 295 34738 347
rect 34088 68 34141 120
rect 34088 4 34141 56
<< metal2 >>
rect 41602 23656 42660 23668
rect 41602 23494 42410 23656
rect 42648 23494 42660 23656
rect 41602 23484 42660 23494
rect 42396 23250 42660 23276
rect 42396 22838 42422 23250
rect 42634 22838 42660 23250
rect 42396 22814 42660 22838
rect 41602 22788 42164 22806
rect 41602 22638 41930 22788
rect 42142 22638 42164 22788
rect 41602 22624 42164 22638
rect 41602 22246 42164 22264
rect 41602 22096 41930 22246
rect 42142 22096 42164 22246
rect 41602 22082 42164 22096
rect 41602 21690 42164 21708
rect 41602 21540 41930 21690
rect 42142 21540 42164 21690
rect 41602 21526 42164 21540
rect 42396 21492 42660 21518
rect 42396 21080 42422 21492
rect 42634 21080 42660 21492
rect 42396 21056 42660 21080
rect 41602 20546 42660 20558
rect 41602 20384 42410 20546
rect 42648 20384 42660 20546
rect 41602 20374 42660 20384
rect 1884 20104 2176 20120
rect 1884 19946 1898 20104
rect 2160 19946 2176 20104
rect 1884 19934 2176 19946
rect 5012 20104 5304 20120
rect 5012 19946 5026 20104
rect 5288 19946 5304 20104
rect 5012 19934 5304 19946
rect 5884 20104 6176 20120
rect 5884 19946 5898 20104
rect 6160 19946 6176 20104
rect 5884 19934 6176 19946
rect 9012 20104 9304 20120
rect 9012 19946 9026 20104
rect 9288 19946 9304 20104
rect 9012 19934 9304 19946
rect 9884 20104 10176 20120
rect 9884 19946 9898 20104
rect 10160 19946 10176 20104
rect 9884 19934 10176 19946
rect 13012 20104 13304 20120
rect 13012 19946 13026 20104
rect 13288 19946 13304 20104
rect 13012 19934 13304 19946
rect 13884 20104 14176 20120
rect 13884 19946 13898 20104
rect 14160 19946 14176 20104
rect 13884 19934 14176 19946
rect 17012 20104 17304 20120
rect 17012 19946 17026 20104
rect 17288 19946 17304 20104
rect 17012 19934 17304 19946
rect 17884 20104 18176 20120
rect 17884 19946 17898 20104
rect 18160 19946 18176 20104
rect 17884 19934 18176 19946
rect 21012 20104 21304 20120
rect 21012 19946 21026 20104
rect 21288 19946 21304 20104
rect 21012 19934 21304 19946
rect 21884 20104 22176 20120
rect 21884 19946 21898 20104
rect 22160 19946 22176 20104
rect 21884 19934 22176 19946
rect 25012 20104 25304 20120
rect 25012 19946 25026 20104
rect 25288 19946 25304 20104
rect 25012 19934 25304 19946
rect 25884 20104 26176 20120
rect 25884 19946 25898 20104
rect 26160 19946 26176 20104
rect 25884 19934 26176 19946
rect 29012 20104 29304 20120
rect 29012 19946 29026 20104
rect 29288 19946 29304 20104
rect 29012 19934 29304 19946
rect 29884 20104 30176 20120
rect 29884 19946 29898 20104
rect 30160 19946 30176 20104
rect 29884 19934 30176 19946
rect 33012 20104 33304 20120
rect 33012 19946 33026 20104
rect 33288 19946 33304 20104
rect 33012 19934 33304 19946
rect 33884 20104 34176 20120
rect 33884 19946 33898 20104
rect 34160 19946 34176 20104
rect 37012 20104 37304 20120
rect 37012 19980 37026 20104
rect 37288 19980 37304 20104
rect 37012 19968 37304 19980
rect 33884 19934 34176 19946
rect 570 19889 984 19900
rect 570 19634 587 19889
rect 969 19634 984 19889
rect 570 19620 984 19634
rect 1046 19620 1460 19900
rect 3420 19882 3790 19900
rect 3420 19638 3444 19882
rect 3770 19638 3790 19882
rect 3420 19620 3790 19638
rect 7420 19882 7790 19900
rect 7420 19638 7444 19882
rect 7770 19638 7790 19882
rect 7420 19620 7790 19638
rect 11420 19882 11790 19900
rect 11420 19638 11444 19882
rect 11770 19638 11790 19882
rect 11420 19620 11790 19638
rect 15420 19882 15790 19900
rect 15420 19638 15444 19882
rect 15770 19638 15790 19882
rect 15420 19620 15790 19638
rect 19420 19882 19790 19900
rect 19420 19638 19444 19882
rect 19770 19638 19790 19882
rect 19420 19620 19790 19638
rect 23420 19882 23790 19900
rect 23420 19638 23444 19882
rect 23770 19638 23790 19882
rect 23420 19620 23790 19638
rect 27420 19882 27790 19900
rect 27420 19638 27444 19882
rect 27770 19638 27790 19882
rect 27420 19620 27790 19638
rect 31420 19882 31790 19900
rect 31420 19638 31444 19882
rect 31770 19638 31790 19882
rect 36540 19885 36954 19900
rect 35396 19847 35810 19862
rect 35396 19783 35426 19847
rect 35490 19783 35522 19847
rect 35586 19783 35618 19847
rect 35682 19783 35714 19847
rect 35778 19783 35810 19847
rect 35396 19753 35810 19783
rect 35396 19689 35426 19753
rect 35490 19689 35522 19753
rect 35586 19689 35618 19753
rect 35682 19689 35714 19753
rect 35778 19689 35810 19753
rect 36540 19821 36570 19885
rect 36634 19821 36666 19885
rect 36730 19821 36762 19885
rect 36826 19821 36858 19885
rect 36922 19821 36954 19885
rect 36540 19791 36954 19821
rect 36540 19727 36570 19791
rect 36634 19727 36666 19791
rect 36730 19727 36762 19791
rect 36826 19727 36858 19791
rect 36922 19727 36954 19791
rect 36540 19692 36954 19727
rect 35396 19655 35810 19689
rect 31420 19620 31790 19638
rect 36064 19557 36478 19585
rect 36064 19493 36094 19557
rect 36158 19493 36190 19557
rect 36254 19493 36286 19557
rect 36350 19493 36382 19557
rect 36446 19493 36478 19557
rect 36064 19466 36478 19493
rect 1046 19451 1460 19462
rect 1046 19196 1063 19451
rect 1445 19196 1460 19451
rect 1046 19182 1460 19196
rect 1884 19442 2176 19462
rect 1884 19386 1904 19442
rect 1960 19386 1998 19442
rect 2054 19386 2092 19442
rect 2148 19386 2176 19442
rect 1884 19348 2176 19386
rect 1884 19292 1904 19348
rect 1960 19292 1998 19348
rect 2054 19292 2092 19348
rect 2148 19292 2176 19348
rect 1884 19254 2176 19292
rect 1884 19198 1904 19254
rect 1960 19198 1998 19254
rect 2054 19198 2092 19254
rect 2148 19198 2176 19254
rect 1884 19182 2176 19198
rect 5012 19442 5304 19462
rect 5012 19386 5032 19442
rect 5088 19386 5126 19442
rect 5182 19386 5220 19442
rect 5276 19386 5304 19442
rect 5012 19348 5304 19386
rect 5012 19292 5032 19348
rect 5088 19292 5126 19348
rect 5182 19292 5220 19348
rect 5276 19292 5304 19348
rect 5012 19254 5304 19292
rect 5012 19198 5032 19254
rect 5088 19198 5126 19254
rect 5182 19198 5220 19254
rect 5276 19198 5304 19254
rect 5012 19182 5304 19198
rect 5884 19442 6176 19462
rect 5884 19386 5904 19442
rect 5960 19386 5998 19442
rect 6054 19386 6092 19442
rect 6148 19386 6176 19442
rect 5884 19348 6176 19386
rect 5884 19292 5904 19348
rect 5960 19292 5998 19348
rect 6054 19292 6092 19348
rect 6148 19292 6176 19348
rect 5884 19254 6176 19292
rect 5884 19198 5904 19254
rect 5960 19198 5998 19254
rect 6054 19198 6092 19254
rect 6148 19198 6176 19254
rect 5884 19182 6176 19198
rect 9012 19442 9304 19462
rect 9012 19386 9032 19442
rect 9088 19386 9126 19442
rect 9182 19386 9220 19442
rect 9276 19386 9304 19442
rect 9012 19348 9304 19386
rect 9012 19292 9032 19348
rect 9088 19292 9126 19348
rect 9182 19292 9220 19348
rect 9276 19292 9304 19348
rect 9012 19254 9304 19292
rect 9012 19198 9032 19254
rect 9088 19198 9126 19254
rect 9182 19198 9220 19254
rect 9276 19198 9304 19254
rect 9012 19182 9304 19198
rect 9884 19442 10176 19462
rect 9884 19386 9904 19442
rect 9960 19386 9998 19442
rect 10054 19386 10092 19442
rect 10148 19386 10176 19442
rect 9884 19348 10176 19386
rect 9884 19292 9904 19348
rect 9960 19292 9998 19348
rect 10054 19292 10092 19348
rect 10148 19292 10176 19348
rect 9884 19254 10176 19292
rect 9884 19198 9904 19254
rect 9960 19198 9998 19254
rect 10054 19198 10092 19254
rect 10148 19198 10176 19254
rect 9884 19182 10176 19198
rect 13012 19442 13304 19462
rect 13012 19386 13032 19442
rect 13088 19386 13126 19442
rect 13182 19386 13220 19442
rect 13276 19386 13304 19442
rect 13012 19348 13304 19386
rect 13012 19292 13032 19348
rect 13088 19292 13126 19348
rect 13182 19292 13220 19348
rect 13276 19292 13304 19348
rect 13012 19254 13304 19292
rect 13012 19198 13032 19254
rect 13088 19198 13126 19254
rect 13182 19198 13220 19254
rect 13276 19198 13304 19254
rect 13012 19182 13304 19198
rect 13884 19442 14176 19462
rect 13884 19386 13904 19442
rect 13960 19386 13998 19442
rect 14054 19386 14092 19442
rect 14148 19386 14176 19442
rect 13884 19348 14176 19386
rect 13884 19292 13904 19348
rect 13960 19292 13998 19348
rect 14054 19292 14092 19348
rect 14148 19292 14176 19348
rect 13884 19254 14176 19292
rect 13884 19198 13904 19254
rect 13960 19198 13998 19254
rect 14054 19198 14092 19254
rect 14148 19198 14176 19254
rect 13884 19182 14176 19198
rect 17012 19442 17304 19462
rect 17012 19386 17032 19442
rect 17088 19386 17126 19442
rect 17182 19386 17220 19442
rect 17276 19386 17304 19442
rect 17012 19348 17304 19386
rect 17012 19292 17032 19348
rect 17088 19292 17126 19348
rect 17182 19292 17220 19348
rect 17276 19292 17304 19348
rect 17012 19254 17304 19292
rect 17012 19198 17032 19254
rect 17088 19198 17126 19254
rect 17182 19198 17220 19254
rect 17276 19198 17304 19254
rect 17012 19182 17304 19198
rect 17884 19442 18176 19462
rect 17884 19386 17904 19442
rect 17960 19386 17998 19442
rect 18054 19386 18092 19442
rect 18148 19386 18176 19442
rect 17884 19348 18176 19386
rect 17884 19292 17904 19348
rect 17960 19292 17998 19348
rect 18054 19292 18092 19348
rect 18148 19292 18176 19348
rect 17884 19254 18176 19292
rect 17884 19198 17904 19254
rect 17960 19198 17998 19254
rect 18054 19198 18092 19254
rect 18148 19198 18176 19254
rect 17884 19182 18176 19198
rect 21012 19442 21304 19462
rect 21012 19386 21032 19442
rect 21088 19386 21126 19442
rect 21182 19386 21220 19442
rect 21276 19386 21304 19442
rect 21012 19348 21304 19386
rect 21012 19292 21032 19348
rect 21088 19292 21126 19348
rect 21182 19292 21220 19348
rect 21276 19292 21304 19348
rect 21012 19254 21304 19292
rect 21012 19198 21032 19254
rect 21088 19198 21126 19254
rect 21182 19198 21220 19254
rect 21276 19198 21304 19254
rect 21012 19182 21304 19198
rect 21884 19442 22176 19462
rect 21884 19386 21904 19442
rect 21960 19386 21998 19442
rect 22054 19386 22092 19442
rect 22148 19386 22176 19442
rect 21884 19348 22176 19386
rect 21884 19292 21904 19348
rect 21960 19292 21998 19348
rect 22054 19292 22092 19348
rect 22148 19292 22176 19348
rect 21884 19254 22176 19292
rect 21884 19198 21904 19254
rect 21960 19198 21998 19254
rect 22054 19198 22092 19254
rect 22148 19198 22176 19254
rect 21884 19182 22176 19198
rect 25012 19442 25304 19462
rect 25012 19386 25032 19442
rect 25088 19386 25126 19442
rect 25182 19386 25220 19442
rect 25276 19386 25304 19442
rect 25012 19348 25304 19386
rect 25012 19292 25032 19348
rect 25088 19292 25126 19348
rect 25182 19292 25220 19348
rect 25276 19292 25304 19348
rect 25012 19254 25304 19292
rect 25012 19198 25032 19254
rect 25088 19198 25126 19254
rect 25182 19198 25220 19254
rect 25276 19198 25304 19254
rect 25012 19182 25304 19198
rect 25884 19442 26176 19462
rect 25884 19386 25904 19442
rect 25960 19386 25998 19442
rect 26054 19386 26092 19442
rect 26148 19386 26176 19442
rect 25884 19348 26176 19386
rect 25884 19292 25904 19348
rect 25960 19292 25998 19348
rect 26054 19292 26092 19348
rect 26148 19292 26176 19348
rect 25884 19254 26176 19292
rect 25884 19198 25904 19254
rect 25960 19198 25998 19254
rect 26054 19198 26092 19254
rect 26148 19198 26176 19254
rect 25884 19182 26176 19198
rect 29012 19442 29304 19462
rect 29012 19386 29032 19442
rect 29088 19386 29126 19442
rect 29182 19386 29220 19442
rect 29276 19386 29304 19442
rect 29012 19348 29304 19386
rect 29012 19292 29032 19348
rect 29088 19292 29126 19348
rect 29182 19292 29220 19348
rect 29276 19292 29304 19348
rect 29012 19254 29304 19292
rect 29012 19198 29032 19254
rect 29088 19198 29126 19254
rect 29182 19198 29220 19254
rect 29276 19198 29304 19254
rect 29012 19182 29304 19198
rect 29884 19442 30176 19462
rect 29884 19386 29904 19442
rect 29960 19386 29998 19442
rect 30054 19386 30092 19442
rect 30148 19386 30176 19442
rect 29884 19348 30176 19386
rect 29884 19292 29904 19348
rect 29960 19292 29998 19348
rect 30054 19292 30092 19348
rect 30148 19292 30176 19348
rect 29884 19254 30176 19292
rect 29884 19198 29904 19254
rect 29960 19198 29998 19254
rect 30054 19198 30092 19254
rect 30148 19198 30176 19254
rect 29884 19182 30176 19198
rect 33012 19442 33304 19462
rect 33012 19386 33032 19442
rect 33088 19386 33126 19442
rect 33182 19386 33220 19442
rect 33276 19386 33304 19442
rect 33012 19348 33304 19386
rect 33012 19292 33032 19348
rect 33088 19292 33126 19348
rect 33182 19292 33220 19348
rect 33276 19292 33304 19348
rect 33012 19254 33304 19292
rect 33012 19198 33032 19254
rect 33088 19198 33126 19254
rect 33182 19198 33220 19254
rect 33276 19198 33304 19254
rect 33012 19182 33304 19198
rect 33884 19442 34176 19462
rect 33884 19386 33904 19442
rect 33960 19386 33998 19442
rect 34054 19386 34092 19442
rect 34148 19386 34176 19442
rect 33884 19348 34176 19386
rect 33884 19292 33904 19348
rect 33960 19292 33998 19348
rect 34054 19292 34092 19348
rect 34148 19292 34176 19348
rect 33884 19254 34176 19292
rect 33884 19198 33904 19254
rect 33960 19198 33998 19254
rect 34054 19198 34092 19254
rect 34148 19198 34176 19254
rect 33884 19182 34176 19198
rect 36064 19402 36094 19466
rect 36158 19402 36190 19466
rect 36254 19402 36286 19466
rect 36350 19402 36382 19466
rect 36446 19402 36478 19466
rect 36064 19375 36478 19402
rect 36064 19311 36094 19375
rect 36158 19311 36190 19375
rect 36254 19311 36286 19375
rect 36350 19311 36382 19375
rect 36446 19311 36478 19375
rect 36064 19281 36478 19311
rect 36064 19217 36094 19281
rect 36158 19217 36190 19281
rect 36254 19217 36286 19281
rect 36350 19217 36382 19281
rect 36446 19217 36478 19281
rect 36064 19182 36478 19217
rect 182 17748 250 18986
rect 182 17696 188 17748
rect 244 17696 250 17748
rect 182 16744 250 17696
rect 182 16692 188 16744
rect 244 16692 250 16744
rect 182 15740 250 16692
rect 182 15688 188 15740
rect 244 15688 250 15740
rect 182 14736 250 15688
rect 182 14684 188 14736
rect 244 14684 250 14736
rect 182 13732 250 14684
rect 182 13680 188 13732
rect 244 13680 250 13732
rect 182 12728 250 13680
rect 182 12676 188 12728
rect 244 12676 250 12728
rect 182 11724 250 12676
rect 182 11672 188 11724
rect 244 11672 250 11724
rect 182 10720 250 11672
rect 182 10668 188 10720
rect 244 10668 250 10720
rect 182 9716 250 10668
rect 182 9664 188 9716
rect 244 9664 250 9716
rect 182 8712 250 9664
rect 182 8660 188 8712
rect 244 8660 250 8712
rect 182 7708 250 8660
rect 182 7656 188 7708
rect 244 7656 250 7708
rect 182 6704 250 7656
rect 182 6652 188 6704
rect 244 6652 250 6704
rect 182 5700 250 6652
rect 182 5648 188 5700
rect 244 5648 250 5700
rect 182 4696 250 5648
rect 182 4644 188 4696
rect 244 4644 250 4696
rect 182 3692 250 4644
rect 182 3640 188 3692
rect 244 3640 250 3692
rect 182 2688 250 3640
rect 182 2636 188 2688
rect 244 2636 250 2688
rect 182 0 250 2636
rect 290 17380 358 18986
rect 290 17328 296 17380
rect 352 17328 358 17380
rect 290 16376 358 17328
rect 290 16324 296 16376
rect 352 16324 358 16376
rect 290 15372 358 16324
rect 290 15320 296 15372
rect 352 15320 358 15372
rect 290 14368 358 15320
rect 290 14316 296 14368
rect 352 14316 358 14368
rect 290 13364 358 14316
rect 290 13312 296 13364
rect 352 13312 358 13364
rect 290 12360 358 13312
rect 290 12308 296 12360
rect 352 12308 358 12360
rect 290 11356 358 12308
rect 290 11304 296 11356
rect 352 11304 358 11356
rect 290 10352 358 11304
rect 290 10300 296 10352
rect 352 10300 358 10352
rect 290 9348 358 10300
rect 290 9296 296 9348
rect 352 9296 358 9348
rect 290 8344 358 9296
rect 290 8292 296 8344
rect 352 8292 358 8344
rect 290 7340 358 8292
rect 290 7288 296 7340
rect 352 7288 358 7340
rect 290 6336 358 7288
rect 290 6284 296 6336
rect 352 6284 358 6336
rect 290 5332 358 6284
rect 290 5280 296 5332
rect 352 5280 358 5332
rect 290 4328 358 5280
rect 290 4276 296 4328
rect 352 4276 358 4328
rect 290 3324 358 4276
rect 290 3272 296 3324
rect 352 3272 358 3324
rect 290 2320 358 3272
rect 290 2268 296 2320
rect 352 2268 358 2320
rect 290 0 358 2268
rect 398 18242 534 18986
rect 36540 18870 36954 18890
rect 570 18816 984 18836
rect 570 18745 591 18816
rect 662 18745 686 18816
rect 757 18745 795 18816
rect 866 18745 890 18816
rect 961 18745 984 18816
rect 36540 18799 36561 18870
rect 36632 18799 36656 18870
rect 36727 18799 36765 18870
rect 36836 18799 36860 18870
rect 36931 18799 36954 18870
rect 36540 18780 36954 18799
rect 570 18726 984 18745
rect 570 18502 984 18522
rect 570 18431 591 18502
rect 662 18431 686 18502
rect 757 18431 795 18502
rect 866 18431 890 18502
rect 961 18431 984 18502
rect 570 18412 984 18431
rect 1046 18363 1460 18383
rect 1046 18292 1067 18363
rect 1138 18292 1162 18363
rect 1233 18292 1271 18363
rect 1342 18292 1366 18363
rect 1437 18292 1460 18363
rect 1046 18273 1460 18292
rect 37042 18297 37364 19901
rect 41602 19656 42660 19668
rect 37394 19551 37602 19585
rect 37394 19495 37427 19551
rect 37483 19495 37516 19551
rect 37572 19495 37602 19551
rect 37394 19460 37602 19495
rect 41602 19494 42410 19656
rect 42648 19494 42660 19656
rect 41602 19484 42660 19494
rect 37394 19404 37427 19460
rect 37483 19404 37516 19460
rect 37572 19404 37602 19460
rect 37394 19369 37602 19404
rect 37394 19313 37427 19369
rect 37483 19313 37516 19369
rect 37572 19313 37602 19369
rect 37394 19286 37602 19313
rect 37444 19212 37602 19286
rect 37444 19160 37451 19212
rect 37503 19160 37542 19212
rect 37594 19160 37602 19212
rect 37444 19110 37602 19160
rect 37444 19058 37451 19110
rect 37503 19058 37542 19110
rect 37594 19058 37602 19110
rect 37444 19007 37602 19058
rect 37444 18955 37452 19007
rect 37504 18955 37543 19007
rect 37595 18955 37602 19007
rect 37444 18914 37602 18955
rect 37444 18862 37452 18914
rect 37504 18862 37543 18914
rect 37595 18862 37602 18914
rect 37444 18849 37602 18862
rect 42396 19250 42660 19276
rect 42396 18838 42422 19250
rect 42634 18838 42660 19250
rect 42396 18814 42660 18838
rect 41602 18788 42164 18806
rect 41602 18638 41930 18788
rect 42142 18638 42164 18788
rect 41602 18624 42164 18638
rect 398 18190 404 18242
rect 460 18190 472 18242
rect 528 18190 534 18242
rect 398 17238 534 18190
rect 37042 18217 37061 18297
rect 37148 18217 37161 18297
rect 37248 18217 37261 18297
rect 37348 18217 37364 18297
rect 1046 18153 1460 18173
rect 1046 18082 1067 18153
rect 1138 18082 1162 18153
rect 1233 18082 1271 18153
rect 1342 18082 1366 18153
rect 1437 18082 1460 18153
rect 1046 18063 1460 18082
rect 36064 18154 36478 18174
rect 36064 18083 36085 18154
rect 36156 18083 36180 18154
rect 36251 18083 36289 18154
rect 36360 18083 36384 18154
rect 36455 18083 36478 18154
rect 36064 18064 36478 18083
rect 570 17866 984 17886
rect 570 17795 591 17866
rect 662 17795 686 17866
rect 757 17795 795 17866
rect 866 17795 890 17866
rect 961 17795 984 17866
rect 570 17776 984 17795
rect 36540 17866 36954 17886
rect 36540 17795 36561 17866
rect 36632 17795 36656 17866
rect 36727 17795 36765 17866
rect 36836 17795 36860 17866
rect 36931 17795 36954 17866
rect 36540 17776 36954 17795
rect 398 17186 410 17238
rect 524 17186 534 17238
rect 398 16234 534 17186
rect 37042 17293 37364 18217
rect 37392 18307 37602 18332
rect 37392 18243 37431 18307
rect 37495 18243 37602 18307
rect 37392 18195 37602 18243
rect 37392 18131 37430 18195
rect 37494 18131 37602 18195
rect 37392 18077 37602 18131
rect 41602 18246 42164 18264
rect 41602 18096 41930 18246
rect 42142 18096 42164 18246
rect 41602 18082 42164 18096
rect 37392 18013 37430 18077
rect 37494 18013 37602 18077
rect 37392 17988 37602 18013
rect 41602 17690 42164 17708
rect 41602 17540 41930 17690
rect 42142 17540 42164 17690
rect 41602 17526 42164 17540
rect 37042 17213 37061 17293
rect 37148 17213 37161 17293
rect 37248 17213 37261 17293
rect 37348 17213 37364 17293
rect 1046 17150 1460 17170
rect 1046 17079 1067 17150
rect 1138 17079 1162 17150
rect 1233 17079 1271 17150
rect 1342 17079 1366 17150
rect 1437 17079 1460 17150
rect 1046 17060 1460 17079
rect 36064 17150 36478 17170
rect 36064 17079 36085 17150
rect 36156 17079 36180 17150
rect 36251 17079 36289 17150
rect 36360 17079 36384 17150
rect 36455 17079 36478 17150
rect 36064 17060 36478 17079
rect 570 16862 984 16882
rect 570 16791 591 16862
rect 662 16791 686 16862
rect 757 16791 795 16862
rect 866 16791 890 16862
rect 961 16791 984 16862
rect 570 16772 984 16791
rect 36540 16862 36954 16882
rect 36540 16791 36561 16862
rect 36632 16791 36656 16862
rect 36727 16791 36765 16862
rect 36836 16791 36860 16862
rect 36931 16791 36954 16862
rect 36540 16772 36954 16791
rect 36064 16652 36478 16680
rect 36064 16588 36094 16652
rect 36158 16588 36190 16652
rect 36254 16588 36286 16652
rect 36350 16588 36382 16652
rect 36446 16588 36478 16652
rect 36064 16561 36478 16588
rect 36064 16497 36094 16561
rect 36158 16497 36190 16561
rect 36254 16497 36286 16561
rect 36350 16497 36382 16561
rect 36446 16497 36478 16561
rect 36064 16470 36478 16497
rect 36064 16406 36094 16470
rect 36158 16406 36190 16470
rect 36254 16406 36286 16470
rect 36350 16406 36382 16470
rect 36446 16406 36478 16470
rect 36064 16381 36478 16406
rect 398 16182 410 16234
rect 524 16182 534 16234
rect 398 15230 534 16182
rect 37042 16289 37364 17213
rect 37444 17452 37602 17498
rect 37444 17400 37451 17452
rect 37503 17400 37542 17452
rect 37594 17400 37602 17452
rect 37444 17350 37602 17400
rect 37444 17298 37451 17350
rect 37503 17298 37542 17350
rect 37594 17298 37602 17350
rect 37444 17247 37602 17298
rect 37444 17195 37452 17247
rect 37504 17195 37543 17247
rect 37595 17195 37602 17247
rect 37444 17154 37602 17195
rect 37444 17102 37452 17154
rect 37504 17102 37543 17154
rect 37595 17102 37602 17154
rect 37444 17089 37602 17102
rect 42396 17492 42660 17518
rect 42396 17080 42422 17492
rect 42634 17080 42660 17492
rect 42396 17056 42660 17080
rect 37444 16680 37602 17056
rect 37394 16646 37602 16680
rect 37394 16590 37427 16646
rect 37483 16590 37516 16646
rect 37572 16590 37602 16646
rect 37394 16555 37602 16590
rect 37394 16499 37427 16555
rect 37483 16499 37516 16555
rect 37572 16499 37602 16555
rect 37394 16464 37602 16499
rect 37394 16408 37427 16464
rect 37483 16408 37516 16464
rect 37572 16408 37602 16464
rect 37394 16381 37602 16408
rect 37042 16209 37061 16289
rect 37148 16209 37161 16289
rect 37248 16209 37261 16289
rect 37348 16209 37364 16289
rect 1046 16145 1460 16165
rect 1046 16074 1067 16145
rect 1138 16074 1162 16145
rect 1233 16074 1271 16145
rect 1342 16074 1366 16145
rect 1437 16074 1460 16145
rect 1046 16055 1460 16074
rect 36064 16146 36478 16166
rect 36064 16075 36085 16146
rect 36156 16075 36180 16146
rect 36251 16075 36289 16146
rect 36360 16075 36384 16146
rect 36455 16075 36478 16146
rect 36064 16056 36478 16075
rect 570 15858 984 15878
rect 570 15787 591 15858
rect 662 15787 686 15858
rect 757 15787 795 15858
rect 866 15787 890 15858
rect 961 15787 984 15858
rect 570 15768 984 15787
rect 36540 15858 36954 15878
rect 36540 15787 36561 15858
rect 36632 15787 36656 15858
rect 36727 15787 36765 15858
rect 36836 15787 36860 15858
rect 36931 15787 36954 15858
rect 36540 15768 36954 15787
rect 398 15178 410 15230
rect 524 15178 534 15230
rect 398 14226 534 15178
rect 37042 15285 37364 16209
rect 37042 15205 37061 15285
rect 37148 15205 37161 15285
rect 37248 15205 37261 15285
rect 37348 15205 37364 15285
rect 1046 15142 1460 15162
rect 1046 15071 1067 15142
rect 1138 15071 1162 15142
rect 1233 15071 1271 15142
rect 1342 15071 1366 15142
rect 1437 15071 1460 15142
rect 1046 15052 1460 15071
rect 36064 15142 36478 15162
rect 36064 15071 36085 15142
rect 36156 15071 36180 15142
rect 36251 15071 36289 15142
rect 36360 15071 36384 15142
rect 36455 15071 36478 15142
rect 36064 15052 36478 15071
rect 570 14854 984 14874
rect 570 14783 591 14854
rect 662 14783 686 14854
rect 757 14783 795 14854
rect 866 14783 890 14854
rect 961 14783 984 14854
rect 570 14764 984 14783
rect 36540 14854 36954 14874
rect 36540 14783 36561 14854
rect 36632 14783 36656 14854
rect 36727 14783 36765 14854
rect 36836 14783 36860 14854
rect 36931 14783 36954 14854
rect 36540 14764 36954 14783
rect 398 14174 410 14226
rect 524 14174 534 14226
rect 398 13222 534 14174
rect 37042 14281 37364 15205
rect 37444 15212 37602 16381
rect 41602 16546 42660 16558
rect 41602 16384 42410 16546
rect 42648 16384 42660 16546
rect 41602 16374 42660 16384
rect 41602 15656 42660 15668
rect 41602 15494 42410 15656
rect 42648 15494 42660 15656
rect 41602 15484 42660 15494
rect 37444 15160 37451 15212
rect 37503 15160 37542 15212
rect 37594 15160 37602 15212
rect 37444 15110 37602 15160
rect 37444 15058 37451 15110
rect 37503 15058 37542 15110
rect 37594 15058 37602 15110
rect 37444 15007 37602 15058
rect 37444 14955 37452 15007
rect 37504 14955 37543 15007
rect 37595 14955 37602 15007
rect 37444 14914 37602 14955
rect 37444 14862 37452 14914
rect 37504 14862 37543 14914
rect 37595 14862 37602 14914
rect 37444 14850 37602 14862
rect 42396 15250 42660 15276
rect 42396 14838 42422 15250
rect 42634 14838 42660 15250
rect 42396 14814 42660 14838
rect 41602 14788 42164 14806
rect 41602 14638 41930 14788
rect 42142 14638 42164 14788
rect 41602 14624 42164 14638
rect 37042 14201 37061 14281
rect 37148 14201 37161 14281
rect 37248 14201 37261 14281
rect 37348 14201 37364 14281
rect 1046 14138 1460 14158
rect 1046 14067 1067 14138
rect 1138 14067 1162 14138
rect 1233 14067 1271 14138
rect 1342 14067 1366 14138
rect 1437 14067 1460 14138
rect 1046 14048 1460 14067
rect 36064 14138 36478 14158
rect 36064 14067 36085 14138
rect 36156 14067 36180 14138
rect 36251 14067 36289 14138
rect 36360 14067 36384 14138
rect 36455 14067 36478 14138
rect 36064 14048 36478 14067
rect 570 13850 984 13870
rect 570 13779 591 13850
rect 662 13779 686 13850
rect 757 13779 795 13850
rect 866 13779 890 13850
rect 961 13779 984 13850
rect 570 13760 984 13779
rect 36540 13850 36954 13870
rect 36540 13779 36561 13850
rect 36632 13779 36656 13850
rect 36727 13779 36765 13850
rect 36836 13779 36860 13850
rect 36931 13779 36954 13850
rect 36540 13760 36954 13779
rect 398 13170 410 13222
rect 524 13170 534 13222
rect 398 12218 534 13170
rect 37042 13277 37364 14201
rect 37392 14307 37602 14332
rect 37392 14243 37431 14307
rect 37495 14243 37602 14307
rect 37392 14195 37602 14243
rect 37392 14131 37430 14195
rect 37494 14131 37602 14195
rect 37392 14077 37602 14131
rect 41602 14246 42164 14264
rect 41602 14096 41930 14246
rect 42142 14096 42164 14246
rect 41602 14082 42164 14096
rect 37392 14013 37430 14077
rect 37494 14013 37602 14077
rect 37392 13988 37602 14013
rect 41602 13690 42164 13708
rect 41602 13540 41930 13690
rect 42142 13540 42164 13690
rect 41602 13526 42164 13540
rect 37042 13197 37061 13277
rect 37148 13197 37161 13277
rect 37248 13197 37261 13277
rect 37348 13197 37364 13277
rect 1046 13134 1460 13154
rect 1046 13063 1067 13134
rect 1138 13063 1162 13134
rect 1233 13063 1271 13134
rect 1342 13063 1366 13134
rect 1437 13063 1460 13134
rect 1046 13044 1460 13063
rect 36064 13134 36478 13154
rect 36064 13063 36085 13134
rect 36156 13063 36180 13134
rect 36251 13063 36289 13134
rect 36360 13063 36384 13134
rect 36455 13063 36478 13134
rect 36064 13044 36478 13063
rect 570 12846 984 12866
rect 570 12775 591 12846
rect 662 12775 686 12846
rect 757 12775 795 12846
rect 866 12775 890 12846
rect 961 12775 984 12846
rect 570 12756 984 12775
rect 36540 12846 36954 12866
rect 36540 12775 36561 12846
rect 36632 12775 36656 12846
rect 36727 12775 36765 12846
rect 36836 12775 36860 12846
rect 36931 12775 36954 12846
rect 36540 12756 36954 12775
rect 36064 12594 36478 12622
rect 36064 12530 36094 12594
rect 36158 12530 36190 12594
rect 36254 12530 36286 12594
rect 36350 12530 36382 12594
rect 36446 12530 36478 12594
rect 36064 12503 36478 12530
rect 36064 12439 36094 12503
rect 36158 12439 36190 12503
rect 36254 12439 36286 12503
rect 36350 12439 36382 12503
rect 36446 12439 36478 12503
rect 36064 12412 36478 12439
rect 36064 12348 36094 12412
rect 36158 12348 36190 12412
rect 36254 12348 36286 12412
rect 36350 12348 36382 12412
rect 36446 12348 36478 12412
rect 36064 12323 36478 12348
rect 398 12166 410 12218
rect 524 12166 534 12218
rect 398 11214 534 12166
rect 37042 12273 37364 13197
rect 37444 13452 37602 13498
rect 37444 13400 37451 13452
rect 37503 13400 37542 13452
rect 37594 13400 37602 13452
rect 37444 13350 37602 13400
rect 37444 13298 37451 13350
rect 37503 13298 37542 13350
rect 37594 13298 37602 13350
rect 37444 13247 37602 13298
rect 37444 13195 37452 13247
rect 37504 13195 37543 13247
rect 37595 13195 37602 13247
rect 37444 13154 37602 13195
rect 37444 13102 37452 13154
rect 37504 13102 37543 13154
rect 37595 13102 37602 13154
rect 37444 12622 37602 13102
rect 42396 13492 42660 13518
rect 42396 13080 42422 13492
rect 42634 13080 42660 13492
rect 42396 13056 42660 13080
rect 37394 12588 37602 12622
rect 37394 12532 37427 12588
rect 37483 12532 37516 12588
rect 37572 12532 37602 12588
rect 37394 12497 37602 12532
rect 37394 12441 37427 12497
rect 37483 12441 37516 12497
rect 37572 12441 37602 12497
rect 37394 12406 37602 12441
rect 37394 12350 37427 12406
rect 37483 12350 37516 12406
rect 37572 12350 37602 12406
rect 41602 12546 42660 12558
rect 41602 12384 42410 12546
rect 42648 12384 42660 12546
rect 41602 12374 42660 12384
rect 37394 12323 37602 12350
rect 37042 12193 37061 12273
rect 37148 12193 37161 12273
rect 37248 12193 37261 12273
rect 37348 12193 37364 12273
rect 1046 12130 1460 12150
rect 1046 12059 1067 12130
rect 1138 12059 1162 12130
rect 1233 12059 1271 12130
rect 1342 12059 1366 12130
rect 1437 12059 1460 12130
rect 1046 12040 1460 12059
rect 36064 12130 36478 12150
rect 36064 12059 36085 12130
rect 36156 12059 36180 12130
rect 36251 12059 36289 12130
rect 36360 12059 36384 12130
rect 36455 12059 36478 12130
rect 36064 12040 36478 12059
rect 570 11842 984 11862
rect 570 11771 591 11842
rect 662 11771 686 11842
rect 757 11771 795 11842
rect 866 11771 890 11842
rect 961 11771 984 11842
rect 570 11752 984 11771
rect 36540 11842 36954 11862
rect 36540 11771 36561 11842
rect 36632 11771 36656 11842
rect 36727 11771 36765 11842
rect 36836 11771 36860 11842
rect 36931 11771 36954 11842
rect 36540 11752 36954 11771
rect 398 11162 410 11214
rect 524 11162 534 11214
rect 398 10210 534 11162
rect 37042 11269 37364 12193
rect 37042 11189 37061 11269
rect 37148 11189 37161 11269
rect 37248 11189 37261 11269
rect 37348 11189 37364 11269
rect 1046 11126 1460 11146
rect 1046 11055 1067 11126
rect 1138 11055 1162 11126
rect 1233 11055 1271 11126
rect 1342 11055 1366 11126
rect 1437 11055 1460 11126
rect 1046 11036 1460 11055
rect 36064 11126 36478 11146
rect 36064 11055 36085 11126
rect 36156 11055 36180 11126
rect 36251 11055 36289 11126
rect 36360 11055 36384 11126
rect 36455 11055 36478 11126
rect 36064 11036 36478 11055
rect 570 10838 984 10858
rect 570 10767 591 10838
rect 662 10767 686 10838
rect 757 10767 795 10838
rect 866 10767 890 10838
rect 961 10767 984 10838
rect 570 10748 984 10767
rect 36540 10838 36954 10858
rect 36540 10767 36561 10838
rect 36632 10767 36656 10838
rect 36727 10767 36765 10838
rect 36836 10767 36860 10838
rect 36931 10767 36954 10838
rect 36540 10748 36954 10767
rect 398 10158 410 10210
rect 524 10158 534 10210
rect 398 9206 534 10158
rect 37042 10265 37364 11189
rect 37444 11212 37602 12323
rect 41602 11656 42660 11668
rect 41602 11494 42410 11656
rect 42648 11494 42660 11656
rect 41602 11484 42660 11494
rect 37444 11160 37451 11212
rect 37503 11160 37542 11212
rect 37594 11160 37602 11212
rect 37444 11110 37602 11160
rect 37444 11058 37451 11110
rect 37503 11058 37542 11110
rect 37594 11058 37602 11110
rect 37444 11007 37602 11058
rect 37444 10955 37452 11007
rect 37504 10955 37543 11007
rect 37595 10955 37602 11007
rect 37444 10914 37602 10955
rect 37444 10862 37452 10914
rect 37504 10862 37543 10914
rect 37595 10862 37602 10914
rect 37444 10849 37602 10862
rect 42396 11250 42660 11276
rect 42396 10838 42422 11250
rect 42634 10838 42660 11250
rect 42396 10814 42660 10838
rect 41602 10788 42164 10806
rect 41602 10638 41930 10788
rect 42142 10638 42164 10788
rect 41602 10624 42164 10638
rect 37042 10185 37061 10265
rect 37148 10185 37161 10265
rect 37248 10185 37261 10265
rect 37348 10185 37364 10265
rect 1046 10122 1460 10142
rect 1046 10051 1067 10122
rect 1138 10051 1162 10122
rect 1233 10051 1271 10122
rect 1342 10051 1366 10122
rect 1437 10051 1460 10122
rect 1046 10032 1460 10051
rect 36064 10122 36478 10142
rect 36064 10051 36085 10122
rect 36156 10051 36180 10122
rect 36251 10051 36289 10122
rect 36360 10051 36384 10122
rect 36455 10051 36478 10122
rect 36064 10032 36478 10051
rect 570 9834 984 9854
rect 570 9763 591 9834
rect 662 9763 686 9834
rect 757 9763 795 9834
rect 866 9763 890 9834
rect 961 9763 984 9834
rect 570 9744 984 9763
rect 36540 9834 36954 9854
rect 36540 9763 36561 9834
rect 36632 9763 36656 9834
rect 36727 9763 36765 9834
rect 36836 9763 36860 9834
rect 36931 9763 36954 9834
rect 36540 9744 36954 9763
rect 398 9154 410 9206
rect 524 9154 534 9206
rect 398 8202 534 9154
rect 37042 9261 37364 10185
rect 37392 10307 37602 10332
rect 37392 10243 37431 10307
rect 37495 10243 37602 10307
rect 37392 10195 37602 10243
rect 37392 10131 37430 10195
rect 37494 10131 37602 10195
rect 37392 10077 37602 10131
rect 41602 10246 42164 10264
rect 41602 10096 41930 10246
rect 42142 10096 42164 10246
rect 41602 10082 42164 10096
rect 37392 10013 37430 10077
rect 37494 10013 37602 10077
rect 37392 9988 37602 10013
rect 41602 9690 42164 9708
rect 41602 9540 41930 9690
rect 42142 9540 42164 9690
rect 41602 9526 42164 9540
rect 37042 9181 37061 9261
rect 37148 9181 37161 9261
rect 37248 9181 37261 9261
rect 37348 9181 37364 9261
rect 1046 9118 1460 9138
rect 1046 9047 1067 9118
rect 1138 9047 1162 9118
rect 1233 9047 1271 9118
rect 1342 9047 1366 9118
rect 1437 9047 1460 9118
rect 1046 9028 1460 9047
rect 36064 9118 36478 9138
rect 36064 9047 36085 9118
rect 36156 9047 36180 9118
rect 36251 9047 36289 9118
rect 36360 9047 36384 9118
rect 36455 9047 36478 9118
rect 36064 9028 36478 9047
rect 570 8830 984 8850
rect 570 8759 591 8830
rect 662 8759 686 8830
rect 757 8759 795 8830
rect 866 8759 890 8830
rect 961 8759 984 8830
rect 570 8740 984 8759
rect 36540 8830 36954 8850
rect 36540 8759 36561 8830
rect 36632 8759 36656 8830
rect 36727 8759 36765 8830
rect 36836 8759 36860 8830
rect 36931 8759 36954 8830
rect 36540 8740 36954 8759
rect 36064 8501 36478 8529
rect 36064 8437 36094 8501
rect 36158 8437 36190 8501
rect 36254 8437 36286 8501
rect 36350 8437 36382 8501
rect 36446 8437 36478 8501
rect 36064 8410 36478 8437
rect 36064 8346 36094 8410
rect 36158 8346 36190 8410
rect 36254 8346 36286 8410
rect 36350 8346 36382 8410
rect 36446 8346 36478 8410
rect 36064 8319 36478 8346
rect 36064 8255 36094 8319
rect 36158 8255 36190 8319
rect 36254 8255 36286 8319
rect 36350 8255 36382 8319
rect 36446 8255 36478 8319
rect 36064 8230 36478 8255
rect 37042 8257 37364 9181
rect 37444 9452 37602 9498
rect 37444 9400 37451 9452
rect 37503 9400 37542 9452
rect 37594 9400 37602 9452
rect 37444 9350 37602 9400
rect 37444 9298 37451 9350
rect 37503 9298 37542 9350
rect 37594 9298 37602 9350
rect 37444 9247 37602 9298
rect 37444 9195 37452 9247
rect 37504 9195 37543 9247
rect 37595 9195 37602 9247
rect 37444 9154 37602 9195
rect 37444 9102 37452 9154
rect 37504 9102 37543 9154
rect 37595 9102 37602 9154
rect 37444 8529 37602 9102
rect 42396 9492 42660 9518
rect 42396 9080 42422 9492
rect 42634 9080 42660 9492
rect 42396 9056 42660 9080
rect 398 8150 410 8202
rect 524 8150 534 8202
rect 398 7198 534 8150
rect 37042 8177 37061 8257
rect 37148 8177 37161 8257
rect 37248 8177 37261 8257
rect 37348 8177 37364 8257
rect 37394 8495 37602 8529
rect 37394 8439 37427 8495
rect 37483 8439 37516 8495
rect 37572 8439 37602 8495
rect 37394 8404 37602 8439
rect 37394 8348 37427 8404
rect 37483 8348 37516 8404
rect 37572 8348 37602 8404
rect 41602 8546 42660 8558
rect 41602 8384 42410 8546
rect 42648 8384 42660 8546
rect 41602 8374 42660 8384
rect 37394 8313 37602 8348
rect 37394 8257 37427 8313
rect 37483 8257 37516 8313
rect 37572 8257 37602 8313
rect 37394 8230 37602 8257
rect 1046 8114 1460 8134
rect 1046 8043 1067 8114
rect 1138 8043 1162 8114
rect 1233 8043 1271 8114
rect 1342 8043 1366 8114
rect 1437 8043 1460 8114
rect 1046 8024 1460 8043
rect 36064 8114 36478 8134
rect 36064 8043 36085 8114
rect 36156 8043 36180 8114
rect 36251 8043 36289 8114
rect 36360 8043 36384 8114
rect 36455 8043 36478 8114
rect 36064 8024 36478 8043
rect 570 7826 984 7846
rect 570 7755 591 7826
rect 662 7755 686 7826
rect 757 7755 795 7826
rect 866 7755 890 7826
rect 961 7755 984 7826
rect 570 7736 984 7755
rect 36540 7826 36954 7846
rect 36540 7755 36561 7826
rect 36632 7755 36656 7826
rect 36727 7755 36765 7826
rect 36836 7755 36860 7826
rect 36931 7755 36954 7826
rect 36540 7736 36954 7755
rect 398 7146 410 7198
rect 524 7146 534 7198
rect 398 6194 534 7146
rect 37042 7253 37364 8177
rect 37042 7173 37061 7253
rect 37148 7173 37161 7253
rect 37248 7173 37261 7253
rect 37348 7173 37364 7253
rect 1046 7110 1460 7130
rect 1046 7039 1067 7110
rect 1138 7039 1162 7110
rect 1233 7039 1271 7110
rect 1342 7039 1366 7110
rect 1437 7039 1460 7110
rect 1046 7020 1460 7039
rect 36064 7110 36478 7130
rect 36064 7039 36085 7110
rect 36156 7039 36180 7110
rect 36251 7039 36289 7110
rect 36360 7039 36384 7110
rect 36455 7039 36478 7110
rect 36064 7020 36478 7039
rect 570 6822 984 6842
rect 570 6751 591 6822
rect 662 6751 686 6822
rect 757 6751 795 6822
rect 866 6751 890 6822
rect 961 6751 984 6822
rect 570 6732 984 6751
rect 36540 6822 36954 6842
rect 36540 6751 36561 6822
rect 36632 6751 36656 6822
rect 36727 6751 36765 6822
rect 36836 6751 36860 6822
rect 36931 6751 36954 6822
rect 36540 6732 36954 6751
rect 398 6142 410 6194
rect 524 6142 534 6194
rect 398 5190 534 6142
rect 37042 6249 37364 7173
rect 37444 7212 37602 8230
rect 41602 7656 42660 7668
rect 41602 7494 42410 7656
rect 42648 7494 42660 7656
rect 41602 7484 42660 7494
rect 37444 7160 37451 7212
rect 37503 7160 37542 7212
rect 37594 7160 37602 7212
rect 37444 7110 37602 7160
rect 37444 7058 37451 7110
rect 37503 7058 37542 7110
rect 37594 7058 37602 7110
rect 37444 7007 37602 7058
rect 37444 6955 37452 7007
rect 37504 6955 37543 7007
rect 37595 6955 37602 7007
rect 37444 6914 37602 6955
rect 37444 6862 37452 6914
rect 37504 6862 37543 6914
rect 37595 6862 37602 6914
rect 37444 6849 37602 6862
rect 42396 7250 42660 7276
rect 42396 6838 42422 7250
rect 42634 6838 42660 7250
rect 42396 6814 42660 6838
rect 41602 6788 42164 6806
rect 41602 6638 41930 6788
rect 42142 6638 42164 6788
rect 41602 6624 42164 6638
rect 37042 6169 37061 6249
rect 37148 6169 37161 6249
rect 37248 6169 37261 6249
rect 37348 6169 37364 6249
rect 1046 6106 1460 6126
rect 1046 6035 1067 6106
rect 1138 6035 1162 6106
rect 1233 6035 1271 6106
rect 1342 6035 1366 6106
rect 1437 6035 1460 6106
rect 1046 6016 1460 6035
rect 36064 6106 36478 6126
rect 36064 6035 36085 6106
rect 36156 6035 36180 6106
rect 36251 6035 36289 6106
rect 36360 6035 36384 6106
rect 36455 6035 36478 6106
rect 36064 6016 36478 6035
rect 570 5818 984 5838
rect 570 5747 591 5818
rect 662 5747 686 5818
rect 757 5747 795 5818
rect 866 5747 890 5818
rect 961 5747 984 5818
rect 570 5728 984 5747
rect 36540 5818 36954 5838
rect 36540 5747 36561 5818
rect 36632 5747 36656 5818
rect 36727 5747 36765 5818
rect 36836 5747 36860 5818
rect 36931 5747 36954 5818
rect 36540 5728 36954 5747
rect 398 5138 410 5190
rect 524 5138 534 5190
rect 398 4186 534 5138
rect 37042 5245 37364 6169
rect 37392 6305 37602 6330
rect 37392 6241 37431 6305
rect 37495 6241 37602 6305
rect 37392 6193 37602 6241
rect 37392 6129 37430 6193
rect 37494 6129 37602 6193
rect 37392 6075 37602 6129
rect 41602 6246 42164 6264
rect 41602 6096 41930 6246
rect 42142 6096 42164 6246
rect 41602 6082 42164 6096
rect 37392 6011 37430 6075
rect 37494 6011 37602 6075
rect 37392 5986 37602 6011
rect 41602 5690 42164 5708
rect 41602 5540 41930 5690
rect 42142 5540 42164 5690
rect 41602 5526 42164 5540
rect 37042 5165 37061 5245
rect 37148 5165 37161 5245
rect 37248 5165 37261 5245
rect 37348 5165 37364 5245
rect 1046 5102 1460 5122
rect 1046 5031 1067 5102
rect 1138 5031 1162 5102
rect 1233 5031 1271 5102
rect 1342 5031 1366 5102
rect 1437 5031 1460 5102
rect 1046 5012 1460 5031
rect 36064 5102 36478 5122
rect 36064 5031 36085 5102
rect 36156 5031 36180 5102
rect 36251 5031 36289 5102
rect 36360 5031 36384 5102
rect 36455 5031 36478 5102
rect 36064 5012 36478 5031
rect 570 4814 984 4834
rect 570 4743 591 4814
rect 662 4743 686 4814
rect 757 4743 795 4814
rect 866 4743 890 4814
rect 961 4743 984 4814
rect 570 4724 984 4743
rect 36540 4814 36954 4834
rect 36540 4743 36561 4814
rect 36632 4743 36656 4814
rect 36727 4743 36765 4814
rect 36836 4743 36860 4814
rect 36931 4743 36954 4814
rect 36540 4724 36954 4743
rect 398 4134 410 4186
rect 524 4134 534 4186
rect 398 3182 534 4134
rect 37042 4241 37364 5165
rect 37042 4161 37061 4241
rect 37148 4161 37161 4241
rect 37248 4161 37261 4241
rect 37348 4161 37364 4241
rect 1046 4098 1460 4118
rect 1046 4027 1067 4098
rect 1138 4027 1162 4098
rect 1233 4027 1271 4098
rect 1342 4027 1366 4098
rect 1437 4027 1460 4098
rect 1046 4008 1460 4027
rect 36064 4098 36478 4118
rect 36064 4027 36085 4098
rect 36156 4027 36180 4098
rect 36251 4027 36289 4098
rect 36360 4027 36384 4098
rect 36455 4027 36478 4098
rect 36064 4008 36478 4027
rect 570 3810 984 3830
rect 570 3739 591 3810
rect 662 3739 686 3810
rect 757 3739 795 3810
rect 866 3739 890 3810
rect 961 3739 984 3810
rect 570 3720 984 3739
rect 36540 3810 36954 3830
rect 36540 3739 36561 3810
rect 36632 3739 36656 3810
rect 36727 3739 36765 3810
rect 36836 3739 36860 3810
rect 36931 3739 36954 3810
rect 36540 3720 36954 3739
rect 36064 3589 36478 3617
rect 36064 3525 36094 3589
rect 36158 3525 36190 3589
rect 36254 3525 36286 3589
rect 36350 3525 36382 3589
rect 36446 3525 36478 3589
rect 36064 3498 36478 3525
rect 36064 3434 36094 3498
rect 36158 3434 36190 3498
rect 36254 3434 36286 3498
rect 36350 3434 36382 3498
rect 36446 3434 36478 3498
rect 36064 3407 36478 3434
rect 36064 3343 36094 3407
rect 36158 3343 36190 3407
rect 36254 3343 36286 3407
rect 36350 3343 36382 3407
rect 36446 3343 36478 3407
rect 36064 3318 36478 3343
rect 398 3130 410 3182
rect 524 3130 534 3182
rect 398 2178 534 3130
rect 37042 3237 37364 4161
rect 37444 5452 37602 5498
rect 37444 5400 37451 5452
rect 37503 5400 37542 5452
rect 37594 5400 37602 5452
rect 37444 5350 37602 5400
rect 37444 5298 37451 5350
rect 37503 5298 37542 5350
rect 37594 5298 37602 5350
rect 37444 5247 37602 5298
rect 37444 5195 37452 5247
rect 37504 5195 37543 5247
rect 37595 5195 37602 5247
rect 37444 5154 37602 5195
rect 37444 5102 37452 5154
rect 37504 5102 37543 5154
rect 37595 5102 37602 5154
rect 37444 3617 37602 5102
rect 42396 5492 42660 5518
rect 42396 5080 42422 5492
rect 42634 5080 42660 5492
rect 42396 5056 42660 5080
rect 41602 4546 42660 4558
rect 41602 4384 42410 4546
rect 42648 4384 42660 4546
rect 41602 4374 42660 4384
rect 37394 3583 37602 3617
rect 37394 3527 37427 3583
rect 37483 3527 37516 3583
rect 37572 3527 37602 3583
rect 37394 3492 37602 3527
rect 37394 3436 37427 3492
rect 37483 3436 37516 3492
rect 37572 3436 37602 3492
rect 41602 3656 42660 3668
rect 41602 3494 42410 3656
rect 42648 3494 42660 3656
rect 41602 3484 42660 3494
rect 37394 3401 37602 3436
rect 37394 3345 37427 3401
rect 37483 3345 37516 3401
rect 37572 3345 37602 3401
rect 37394 3318 37602 3345
rect 37042 3157 37061 3237
rect 37148 3157 37161 3237
rect 37248 3157 37261 3237
rect 37348 3157 37364 3237
rect 1046 3092 1460 3112
rect 1046 3021 1067 3092
rect 1138 3021 1162 3092
rect 1233 3021 1271 3092
rect 1342 3021 1366 3092
rect 1437 3021 1460 3092
rect 1046 3002 1460 3021
rect 36064 3094 36478 3114
rect 36064 3023 36085 3094
rect 36156 3023 36180 3094
rect 36251 3023 36289 3094
rect 36360 3023 36384 3094
rect 36455 3023 36478 3094
rect 36064 3004 36478 3023
rect 570 2806 984 2826
rect 570 2735 591 2806
rect 662 2735 686 2806
rect 757 2735 795 2806
rect 866 2735 890 2806
rect 961 2735 984 2806
rect 570 2716 984 2735
rect 36540 2806 36954 2826
rect 36540 2735 36561 2806
rect 36632 2735 36656 2806
rect 36727 2735 36765 2806
rect 36836 2735 36860 2806
rect 36931 2735 36954 2806
rect 36540 2716 36954 2735
rect 398 2126 410 2178
rect 524 2126 534 2178
rect 398 1174 534 2126
rect 37042 2233 37364 3157
rect 37444 3222 37602 3318
rect 37444 3170 37451 3222
rect 37503 3170 37542 3222
rect 37594 3170 37602 3222
rect 37444 3120 37602 3170
rect 37444 3068 37451 3120
rect 37503 3068 37542 3120
rect 37594 3068 37602 3120
rect 37444 3017 37602 3068
rect 37444 2965 37452 3017
rect 37504 2965 37543 3017
rect 37595 2965 37602 3017
rect 37444 2924 37602 2965
rect 37444 2872 37452 2924
rect 37504 2872 37543 2924
rect 37595 2872 37602 2924
rect 37444 2834 37602 2872
rect 42396 3250 42660 3276
rect 42396 2838 42422 3250
rect 42634 2838 42660 3250
rect 42396 2814 42660 2838
rect 41602 2788 42164 2806
rect 41602 2638 41930 2788
rect 42142 2638 42164 2788
rect 41602 2624 42164 2638
rect 37042 2153 37061 2233
rect 37148 2153 37161 2233
rect 37248 2153 37261 2233
rect 37348 2153 37364 2233
rect 1046 2089 1460 2109
rect 1046 2018 1067 2089
rect 1138 2018 1162 2089
rect 1233 2018 1271 2089
rect 1342 2018 1366 2089
rect 1437 2018 1460 2089
rect 1046 1999 1460 2018
rect 36064 2090 36478 2110
rect 36064 2019 36085 2090
rect 36156 2019 36180 2090
rect 36251 2019 36289 2090
rect 36360 2019 36384 2090
rect 36455 2019 36478 2090
rect 36064 2000 36478 2019
rect 36540 1802 36954 1822
rect 570 1748 984 1768
rect 570 1677 591 1748
rect 662 1677 686 1748
rect 757 1677 795 1748
rect 866 1677 890 1748
rect 961 1677 984 1748
rect 36540 1731 36561 1802
rect 36632 1731 36656 1802
rect 36727 1731 36765 1802
rect 36836 1731 36860 1802
rect 36931 1731 36954 1802
rect 36540 1712 36954 1731
rect 570 1658 984 1677
rect 1046 1434 1460 1454
rect 1046 1363 1067 1434
rect 1138 1363 1162 1434
rect 1233 1363 1271 1434
rect 1342 1363 1366 1434
rect 1437 1363 1460 1434
rect 1046 1324 1460 1363
rect 1046 1253 1067 1324
rect 1138 1253 1162 1324
rect 1233 1253 1271 1324
rect 1342 1253 1366 1324
rect 1437 1253 1460 1324
rect 1046 1234 1460 1253
rect 398 1122 410 1174
rect 524 1122 534 1174
rect 398 0 534 1122
rect 37042 1229 37364 2153
rect 37392 2311 37602 2336
rect 37392 2247 37431 2311
rect 37495 2247 37602 2311
rect 37392 2199 37602 2247
rect 37392 2135 37430 2199
rect 37494 2135 37602 2199
rect 37392 2081 37602 2135
rect 41602 2246 42164 2264
rect 41602 2096 41930 2246
rect 42142 2096 42164 2246
rect 41602 2082 42164 2096
rect 37392 2017 37430 2081
rect 37494 2017 37602 2081
rect 37392 1992 37602 2017
rect 41602 1690 42164 1708
rect 41602 1540 41930 1690
rect 42142 1540 42164 1690
rect 41602 1526 42164 1540
rect 37042 1149 37061 1229
rect 37148 1149 37161 1229
rect 37248 1149 37261 1229
rect 37348 1149 37364 1229
rect 1046 1085 1460 1105
rect 1046 1014 1067 1085
rect 1138 1014 1162 1085
rect 1233 1014 1271 1085
rect 1342 1014 1366 1085
rect 1437 1014 1460 1085
rect 1046 995 1460 1014
rect 36064 1086 36478 1106
rect 36064 1015 36085 1086
rect 36156 1015 36180 1086
rect 36251 1015 36289 1086
rect 36360 1015 36384 1086
rect 36455 1015 36478 1086
rect 36064 996 36478 1015
rect 3558 909 3674 914
rect 3558 857 3569 909
rect 3666 857 3674 909
rect 3558 845 3674 857
rect 4194 911 4310 914
rect 4194 859 4205 911
rect 4302 859 4310 911
rect 4194 847 4310 859
rect 4562 910 4678 914
rect 4562 858 4573 910
rect 4670 858 4678 910
rect 570 812 984 832
rect 570 741 591 812
rect 662 741 686 812
rect 757 741 795 812
rect 866 741 890 812
rect 961 772 984 812
rect 961 741 983 772
rect 570 722 983 741
rect 3558 0 3592 845
rect 4230 0 4264 847
rect 4562 846 4678 858
rect 5566 910 5682 914
rect 5566 858 5577 910
rect 5674 858 5682 910
rect 5566 846 5682 858
rect 6570 910 6686 914
rect 6570 858 6581 910
rect 6678 858 6686 910
rect 6570 846 6686 858
rect 7574 910 7690 914
rect 7574 858 7585 910
rect 7682 858 7690 910
rect 7574 846 7690 858
rect 8578 910 8694 914
rect 8578 858 8589 910
rect 8686 858 8694 910
rect 8578 846 8694 858
rect 9582 910 9698 914
rect 9582 858 9593 910
rect 9690 858 9698 910
rect 9582 846 9698 858
rect 10586 910 10702 914
rect 10586 858 10597 910
rect 10694 858 10702 910
rect 10586 846 10702 858
rect 11590 910 11706 914
rect 11590 858 11601 910
rect 11698 858 11706 910
rect 11590 846 11706 858
rect 12594 910 12710 914
rect 12594 858 12605 910
rect 12702 858 12710 910
rect 12594 846 12710 858
rect 13598 910 13714 914
rect 13598 858 13609 910
rect 13706 858 13714 910
rect 13598 846 13714 858
rect 14602 910 14718 914
rect 14602 858 14613 910
rect 14710 858 14718 910
rect 14602 846 14718 858
rect 15606 910 15722 914
rect 15606 858 15617 910
rect 15714 858 15722 910
rect 15606 846 15722 858
rect 16610 910 16726 914
rect 16610 858 16621 910
rect 16718 858 16726 910
rect 16610 846 16726 858
rect 17614 910 17730 914
rect 17614 858 17625 910
rect 17722 858 17730 910
rect 17614 846 17730 858
rect 18244 911 18360 914
rect 18244 859 18255 911
rect 18352 859 18360 911
rect 18244 847 18360 859
rect 18618 910 18734 914
rect 18618 858 18629 910
rect 18726 858 18734 910
rect 4562 0 4596 846
rect 5566 0 5600 846
rect 6570 0 6604 846
rect 7574 0 7608 846
rect 8578 0 8612 846
rect 9582 0 9616 846
rect 10586 0 10620 846
rect 11590 0 11624 846
rect 12594 0 12628 846
rect 13598 0 13632 846
rect 14602 0 14636 846
rect 15606 0 15640 846
rect 16610 0 16644 846
rect 17614 0 17648 846
rect 18286 0 18320 847
rect 18618 846 18734 858
rect 19250 911 19366 914
rect 19250 859 19261 911
rect 19358 859 19366 911
rect 19250 847 19366 859
rect 19622 910 19738 914
rect 19622 858 19633 910
rect 19730 858 19738 910
rect 18618 0 18652 846
rect 19290 0 19324 847
rect 19622 846 19738 858
rect 20246 911 20362 914
rect 20246 859 20257 911
rect 20354 859 20362 911
rect 20246 847 20362 859
rect 20626 910 20742 914
rect 20626 858 20637 910
rect 20734 858 20742 910
rect 19622 0 19656 846
rect 20294 0 20328 847
rect 20626 846 20742 858
rect 21630 910 21746 914
rect 21630 858 21641 910
rect 21738 858 21746 910
rect 21630 846 21746 858
rect 22634 910 22750 914
rect 22634 858 22645 910
rect 22742 858 22750 910
rect 22634 846 22750 858
rect 23638 910 23754 914
rect 23638 858 23649 910
rect 23746 858 23754 910
rect 23638 846 23754 858
rect 24642 910 24758 914
rect 24642 858 24653 910
rect 24750 858 24758 910
rect 24642 846 24758 858
rect 25646 910 25762 914
rect 25646 858 25657 910
rect 25754 858 25762 910
rect 25646 846 25762 858
rect 26650 910 26766 914
rect 26650 858 26661 910
rect 26758 858 26766 910
rect 26650 846 26766 858
rect 27654 910 27770 914
rect 27654 858 27665 910
rect 27762 858 27770 910
rect 27654 846 27770 858
rect 29662 910 29778 914
rect 29662 858 29673 910
rect 29770 858 29778 910
rect 29662 846 29778 858
rect 30666 910 30782 914
rect 30666 858 30677 910
rect 30774 858 30782 910
rect 30666 846 30782 858
rect 31670 910 31786 914
rect 31670 858 31681 910
rect 31778 858 31786 910
rect 31670 846 31786 858
rect 32674 910 32790 914
rect 32674 858 32685 910
rect 32782 858 32790 910
rect 32674 846 32790 858
rect 33600 910 33716 914
rect 33600 858 33611 910
rect 33708 858 33716 910
rect 33600 846 33716 858
rect 34082 907 34147 908
rect 34082 855 34089 907
rect 34141 855 34147 907
rect 20626 0 20660 846
rect 21630 0 21664 846
rect 22634 0 22668 846
rect 23638 0 23672 846
rect 24642 0 24676 846
rect 25646 0 25680 846
rect 26650 0 26684 846
rect 27654 0 27688 846
rect 27848 795 27912 796
rect 27848 743 27854 795
rect 27906 743 27912 795
rect 27848 742 27912 743
rect 27858 0 27892 742
rect 29672 739 29738 846
rect 28052 719 28116 720
rect 28052 667 28058 719
rect 28110 667 28116 719
rect 29672 687 29678 739
rect 29730 687 29738 739
rect 29672 684 29738 687
rect 28052 666 28116 667
rect 28062 0 28096 666
rect 30686 651 30754 846
rect 28251 649 28315 650
rect 28251 597 28257 649
rect 28309 597 28315 649
rect 28251 596 28315 597
rect 30686 599 30696 651
rect 30748 599 30754 651
rect 30686 596 30754 599
rect 28266 0 28300 596
rect 31694 575 31762 846
rect 28455 570 28519 571
rect 28455 518 28461 570
rect 28513 518 28519 570
rect 31694 523 31702 575
rect 31754 523 31762 575
rect 31694 522 31762 523
rect 28455 517 28519 518
rect 28470 0 28504 517
rect 32698 499 32764 846
rect 28659 493 28723 494
rect 28659 441 28665 493
rect 28717 441 28723 493
rect 32698 447 32706 499
rect 32758 447 32764 499
rect 32698 444 32764 447
rect 28659 440 28723 441
rect 28674 0 28708 440
rect 33628 423 33692 846
rect 28863 417 28927 418
rect 28863 365 28869 417
rect 28921 365 28927 417
rect 33628 371 33634 423
rect 33686 371 33692 423
rect 33628 370 33692 371
rect 28863 364 28927 365
rect 28878 0 28912 364
rect 29067 341 29131 342
rect 29067 289 29073 341
rect 29125 289 29131 341
rect 29067 288 29131 289
rect 29082 0 29116 288
rect 34082 120 34147 855
rect 34082 68 34088 120
rect 34141 68 34147 120
rect 34082 56 34147 68
rect 34082 4 34088 56
rect 34141 4 34147 56
rect 34082 3 34147 4
rect 34180 0 34219 914
rect 34554 0 34593 914
rect 34680 910 34798 914
rect 34680 858 34693 910
rect 34790 858 34798 910
rect 34680 846 34798 858
rect 36064 881 36478 909
rect 34680 347 34744 846
rect 36064 817 36094 881
rect 36158 817 36190 881
rect 36254 817 36286 881
rect 36350 817 36382 881
rect 36446 817 36478 881
rect 36064 790 36478 817
rect 36064 726 36094 790
rect 36158 726 36190 790
rect 36254 726 36286 790
rect 36350 726 36382 790
rect 36446 726 36478 790
rect 36064 699 36478 726
rect 36064 635 36094 699
rect 36158 635 36190 699
rect 36254 635 36286 699
rect 36350 635 36382 699
rect 36446 635 36478 699
rect 36064 610 36478 635
rect 36540 526 36954 546
rect 36540 455 36561 526
rect 36632 455 36656 526
rect 36727 455 36765 526
rect 36836 455 36860 526
rect 36931 455 36954 526
rect 36540 436 36954 455
rect 34680 295 34686 347
rect 34738 295 34744 347
rect 34680 294 34744 295
rect 37042 174 37364 1149
rect 37444 1452 37602 1498
rect 37444 1400 37451 1452
rect 37503 1400 37542 1452
rect 37594 1400 37602 1452
rect 37444 1350 37602 1400
rect 37444 1298 37451 1350
rect 37503 1298 37542 1350
rect 37594 1298 37602 1350
rect 37444 1247 37602 1298
rect 37444 1195 37452 1247
rect 37504 1195 37543 1247
rect 37595 1195 37602 1247
rect 37444 1154 37602 1195
rect 37444 1102 37452 1154
rect 37504 1102 37543 1154
rect 37595 1102 37602 1154
rect 37444 909 37602 1102
rect 42396 1492 42660 1518
rect 42396 1080 42422 1492
rect 42634 1080 42660 1492
rect 42396 1056 42660 1080
rect 37394 875 37602 909
rect 37394 819 37427 875
rect 37483 819 37516 875
rect 37572 819 37602 875
rect 37394 784 37602 819
rect 37394 728 37427 784
rect 37483 728 37516 784
rect 37572 728 37602 784
rect 37394 693 37602 728
rect 37394 637 37427 693
rect 37483 637 37516 693
rect 37572 637 37602 693
rect 37394 610 37602 637
rect 41847 557 42660 558
rect 41602 546 42660 557
rect 41602 384 42410 546
rect 42648 384 42660 546
rect 41602 374 42660 384
rect 41602 373 41847 374
<< via2 >>
rect 42410 23494 42648 23656
rect 42422 22838 42634 23250
rect 41930 22638 42142 22788
rect 41930 22096 42142 22246
rect 41930 21540 42142 21690
rect 42422 21080 42634 21492
rect 42410 20384 42648 20546
rect 1898 19946 2160 20104
rect 5026 19946 5288 20104
rect 5898 19946 6160 20104
rect 9026 19946 9288 20104
rect 9898 19946 10160 20104
rect 13026 19946 13288 20104
rect 13898 19946 14160 20104
rect 17026 19946 17288 20104
rect 17898 19946 18160 20104
rect 21026 19946 21288 20104
rect 21898 19946 22160 20104
rect 25026 19946 25288 20104
rect 25898 19946 26160 20104
rect 29026 19946 29288 20104
rect 29898 19946 30160 20104
rect 33026 19946 33288 20104
rect 33898 19946 34160 20104
rect 37026 19980 37288 20104
rect 587 19634 969 19889
rect 3444 19638 3770 19882
rect 7444 19638 7770 19882
rect 11444 19638 11770 19882
rect 15444 19638 15770 19882
rect 19444 19638 19770 19882
rect 23444 19638 23770 19882
rect 27444 19638 27770 19882
rect 31444 19638 31770 19882
rect 35426 19783 35490 19847
rect 35522 19783 35586 19847
rect 35618 19783 35682 19847
rect 35714 19783 35778 19847
rect 35426 19689 35490 19753
rect 35522 19689 35586 19753
rect 35618 19689 35682 19753
rect 35714 19689 35778 19753
rect 36570 19821 36634 19885
rect 36666 19821 36730 19885
rect 36762 19821 36826 19885
rect 36858 19821 36922 19885
rect 36570 19727 36634 19791
rect 36666 19727 36730 19791
rect 36762 19727 36826 19791
rect 36858 19727 36922 19791
rect 36094 19493 36158 19557
rect 36190 19493 36254 19557
rect 36286 19493 36350 19557
rect 36382 19493 36446 19557
rect 1063 19196 1445 19451
rect 1904 19386 1960 19442
rect 1998 19386 2054 19442
rect 2092 19386 2148 19442
rect 1904 19292 1960 19348
rect 1998 19292 2054 19348
rect 2092 19292 2148 19348
rect 1904 19198 1960 19254
rect 1998 19198 2054 19254
rect 2092 19198 2148 19254
rect 5032 19386 5088 19442
rect 5126 19386 5182 19442
rect 5220 19386 5276 19442
rect 5032 19292 5088 19348
rect 5126 19292 5182 19348
rect 5220 19292 5276 19348
rect 5032 19198 5088 19254
rect 5126 19198 5182 19254
rect 5220 19198 5276 19254
rect 5904 19386 5960 19442
rect 5998 19386 6054 19442
rect 6092 19386 6148 19442
rect 5904 19292 5960 19348
rect 5998 19292 6054 19348
rect 6092 19292 6148 19348
rect 5904 19198 5960 19254
rect 5998 19198 6054 19254
rect 6092 19198 6148 19254
rect 9032 19386 9088 19442
rect 9126 19386 9182 19442
rect 9220 19386 9276 19442
rect 9032 19292 9088 19348
rect 9126 19292 9182 19348
rect 9220 19292 9276 19348
rect 9032 19198 9088 19254
rect 9126 19198 9182 19254
rect 9220 19198 9276 19254
rect 9904 19386 9960 19442
rect 9998 19386 10054 19442
rect 10092 19386 10148 19442
rect 9904 19292 9960 19348
rect 9998 19292 10054 19348
rect 10092 19292 10148 19348
rect 9904 19198 9960 19254
rect 9998 19198 10054 19254
rect 10092 19198 10148 19254
rect 13032 19386 13088 19442
rect 13126 19386 13182 19442
rect 13220 19386 13276 19442
rect 13032 19292 13088 19348
rect 13126 19292 13182 19348
rect 13220 19292 13276 19348
rect 13032 19198 13088 19254
rect 13126 19198 13182 19254
rect 13220 19198 13276 19254
rect 13904 19386 13960 19442
rect 13998 19386 14054 19442
rect 14092 19386 14148 19442
rect 13904 19292 13960 19348
rect 13998 19292 14054 19348
rect 14092 19292 14148 19348
rect 13904 19198 13960 19254
rect 13998 19198 14054 19254
rect 14092 19198 14148 19254
rect 17032 19386 17088 19442
rect 17126 19386 17182 19442
rect 17220 19386 17276 19442
rect 17032 19292 17088 19348
rect 17126 19292 17182 19348
rect 17220 19292 17276 19348
rect 17032 19198 17088 19254
rect 17126 19198 17182 19254
rect 17220 19198 17276 19254
rect 17904 19386 17960 19442
rect 17998 19386 18054 19442
rect 18092 19386 18148 19442
rect 17904 19292 17960 19348
rect 17998 19292 18054 19348
rect 18092 19292 18148 19348
rect 17904 19198 17960 19254
rect 17998 19198 18054 19254
rect 18092 19198 18148 19254
rect 21032 19386 21088 19442
rect 21126 19386 21182 19442
rect 21220 19386 21276 19442
rect 21032 19292 21088 19348
rect 21126 19292 21182 19348
rect 21220 19292 21276 19348
rect 21032 19198 21088 19254
rect 21126 19198 21182 19254
rect 21220 19198 21276 19254
rect 21904 19386 21960 19442
rect 21998 19386 22054 19442
rect 22092 19386 22148 19442
rect 21904 19292 21960 19348
rect 21998 19292 22054 19348
rect 22092 19292 22148 19348
rect 21904 19198 21960 19254
rect 21998 19198 22054 19254
rect 22092 19198 22148 19254
rect 25032 19386 25088 19442
rect 25126 19386 25182 19442
rect 25220 19386 25276 19442
rect 25032 19292 25088 19348
rect 25126 19292 25182 19348
rect 25220 19292 25276 19348
rect 25032 19198 25088 19254
rect 25126 19198 25182 19254
rect 25220 19198 25276 19254
rect 25904 19386 25960 19442
rect 25998 19386 26054 19442
rect 26092 19386 26148 19442
rect 25904 19292 25960 19348
rect 25998 19292 26054 19348
rect 26092 19292 26148 19348
rect 25904 19198 25960 19254
rect 25998 19198 26054 19254
rect 26092 19198 26148 19254
rect 29032 19386 29088 19442
rect 29126 19386 29182 19442
rect 29220 19386 29276 19442
rect 29032 19292 29088 19348
rect 29126 19292 29182 19348
rect 29220 19292 29276 19348
rect 29032 19198 29088 19254
rect 29126 19198 29182 19254
rect 29220 19198 29276 19254
rect 29904 19386 29960 19442
rect 29998 19386 30054 19442
rect 30092 19386 30148 19442
rect 29904 19292 29960 19348
rect 29998 19292 30054 19348
rect 30092 19292 30148 19348
rect 29904 19198 29960 19254
rect 29998 19198 30054 19254
rect 30092 19198 30148 19254
rect 33032 19386 33088 19442
rect 33126 19386 33182 19442
rect 33220 19386 33276 19442
rect 33032 19292 33088 19348
rect 33126 19292 33182 19348
rect 33220 19292 33276 19348
rect 33032 19198 33088 19254
rect 33126 19198 33182 19254
rect 33220 19198 33276 19254
rect 33904 19386 33960 19442
rect 33998 19386 34054 19442
rect 34092 19386 34148 19442
rect 33904 19292 33960 19348
rect 33998 19292 34054 19348
rect 34092 19292 34148 19348
rect 33904 19198 33960 19254
rect 33998 19198 34054 19254
rect 34092 19198 34148 19254
rect 36094 19402 36158 19466
rect 36190 19402 36254 19466
rect 36286 19402 36350 19466
rect 36382 19402 36446 19466
rect 36094 19311 36158 19375
rect 36190 19311 36254 19375
rect 36286 19311 36350 19375
rect 36382 19311 36446 19375
rect 36094 19217 36158 19281
rect 36190 19217 36254 19281
rect 36286 19217 36350 19281
rect 36382 19217 36446 19281
rect 591 18745 662 18816
rect 686 18745 757 18816
rect 795 18745 866 18816
rect 890 18745 961 18816
rect 36561 18799 36632 18870
rect 36656 18799 36727 18870
rect 36765 18799 36836 18870
rect 36860 18799 36931 18870
rect 591 18431 662 18502
rect 686 18431 757 18502
rect 795 18431 866 18502
rect 890 18431 961 18502
rect 1067 18292 1138 18363
rect 1162 18292 1233 18363
rect 1271 18292 1342 18363
rect 1366 18292 1437 18363
rect 37427 19495 37483 19551
rect 42410 19494 42648 19656
rect 37427 19404 37483 19460
rect 37427 19313 37483 19369
rect 42422 18838 42634 19250
rect 41930 18638 42142 18788
rect 1067 18082 1138 18153
rect 1162 18082 1233 18153
rect 1271 18082 1342 18153
rect 1366 18082 1437 18153
rect 36085 18083 36156 18154
rect 36180 18083 36251 18154
rect 36289 18083 36360 18154
rect 36384 18083 36455 18154
rect 591 17795 662 17866
rect 686 17795 757 17866
rect 795 17795 866 17866
rect 890 17795 961 17866
rect 36561 17795 36632 17866
rect 36656 17795 36727 17866
rect 36765 17795 36836 17866
rect 36860 17795 36931 17866
rect 37431 18243 37495 18307
rect 37430 18131 37494 18195
rect 41930 18096 42142 18246
rect 37430 18013 37494 18077
rect 41930 17540 42142 17690
rect 1067 17079 1138 17150
rect 1162 17079 1233 17150
rect 1271 17079 1342 17150
rect 1366 17079 1437 17150
rect 36085 17079 36156 17150
rect 36180 17079 36251 17150
rect 36289 17079 36360 17150
rect 36384 17079 36455 17150
rect 591 16791 662 16862
rect 686 16791 757 16862
rect 795 16791 866 16862
rect 890 16791 961 16862
rect 36561 16791 36632 16862
rect 36656 16791 36727 16862
rect 36765 16791 36836 16862
rect 36860 16791 36931 16862
rect 36094 16588 36158 16652
rect 36190 16588 36254 16652
rect 36286 16588 36350 16652
rect 36382 16588 36446 16652
rect 36094 16497 36158 16561
rect 36190 16497 36254 16561
rect 36286 16497 36350 16561
rect 36382 16497 36446 16561
rect 36094 16406 36158 16470
rect 36190 16406 36254 16470
rect 36286 16406 36350 16470
rect 36382 16406 36446 16470
rect 42422 17080 42634 17492
rect 37427 16590 37483 16646
rect 37427 16499 37483 16555
rect 37427 16408 37483 16464
rect 1067 16074 1138 16145
rect 1162 16074 1233 16145
rect 1271 16074 1342 16145
rect 1366 16074 1437 16145
rect 36085 16075 36156 16146
rect 36180 16075 36251 16146
rect 36289 16075 36360 16146
rect 36384 16075 36455 16146
rect 591 15787 662 15858
rect 686 15787 757 15858
rect 795 15787 866 15858
rect 890 15787 961 15858
rect 36561 15787 36632 15858
rect 36656 15787 36727 15858
rect 36765 15787 36836 15858
rect 36860 15787 36931 15858
rect 1067 15071 1138 15142
rect 1162 15071 1233 15142
rect 1271 15071 1342 15142
rect 1366 15071 1437 15142
rect 36085 15071 36156 15142
rect 36180 15071 36251 15142
rect 36289 15071 36360 15142
rect 36384 15071 36455 15142
rect 591 14783 662 14854
rect 686 14783 757 14854
rect 795 14783 866 14854
rect 890 14783 961 14854
rect 36561 14783 36632 14854
rect 36656 14783 36727 14854
rect 36765 14783 36836 14854
rect 36860 14783 36931 14854
rect 42410 16384 42648 16546
rect 42410 15494 42648 15656
rect 42422 14838 42634 15250
rect 41930 14638 42142 14788
rect 1067 14067 1138 14138
rect 1162 14067 1233 14138
rect 1271 14067 1342 14138
rect 1366 14067 1437 14138
rect 36085 14067 36156 14138
rect 36180 14067 36251 14138
rect 36289 14067 36360 14138
rect 36384 14067 36455 14138
rect 591 13779 662 13850
rect 686 13779 757 13850
rect 795 13779 866 13850
rect 890 13779 961 13850
rect 36561 13779 36632 13850
rect 36656 13779 36727 13850
rect 36765 13779 36836 13850
rect 36860 13779 36931 13850
rect 37431 14243 37495 14307
rect 37430 14131 37494 14195
rect 41930 14096 42142 14246
rect 37430 14013 37494 14077
rect 41930 13540 42142 13690
rect 1067 13063 1138 13134
rect 1162 13063 1233 13134
rect 1271 13063 1342 13134
rect 1366 13063 1437 13134
rect 36085 13063 36156 13134
rect 36180 13063 36251 13134
rect 36289 13063 36360 13134
rect 36384 13063 36455 13134
rect 591 12775 662 12846
rect 686 12775 757 12846
rect 795 12775 866 12846
rect 890 12775 961 12846
rect 36561 12775 36632 12846
rect 36656 12775 36727 12846
rect 36765 12775 36836 12846
rect 36860 12775 36931 12846
rect 36094 12530 36158 12594
rect 36190 12530 36254 12594
rect 36286 12530 36350 12594
rect 36382 12530 36446 12594
rect 36094 12439 36158 12503
rect 36190 12439 36254 12503
rect 36286 12439 36350 12503
rect 36382 12439 36446 12503
rect 36094 12348 36158 12412
rect 36190 12348 36254 12412
rect 36286 12348 36350 12412
rect 36382 12348 36446 12412
rect 42422 13080 42634 13492
rect 37427 12532 37483 12588
rect 37427 12441 37483 12497
rect 37427 12350 37483 12406
rect 42410 12384 42648 12546
rect 1067 12059 1138 12130
rect 1162 12059 1233 12130
rect 1271 12059 1342 12130
rect 1366 12059 1437 12130
rect 36085 12059 36156 12130
rect 36180 12059 36251 12130
rect 36289 12059 36360 12130
rect 36384 12059 36455 12130
rect 591 11771 662 11842
rect 686 11771 757 11842
rect 795 11771 866 11842
rect 890 11771 961 11842
rect 36561 11771 36632 11842
rect 36656 11771 36727 11842
rect 36765 11771 36836 11842
rect 36860 11771 36931 11842
rect 1067 11055 1138 11126
rect 1162 11055 1233 11126
rect 1271 11055 1342 11126
rect 1366 11055 1437 11126
rect 36085 11055 36156 11126
rect 36180 11055 36251 11126
rect 36289 11055 36360 11126
rect 36384 11055 36455 11126
rect 591 10767 662 10838
rect 686 10767 757 10838
rect 795 10767 866 10838
rect 890 10767 961 10838
rect 36561 10767 36632 10838
rect 36656 10767 36727 10838
rect 36765 10767 36836 10838
rect 36860 10767 36931 10838
rect 42410 11494 42648 11656
rect 42422 10838 42634 11250
rect 41930 10638 42142 10788
rect 1067 10051 1138 10122
rect 1162 10051 1233 10122
rect 1271 10051 1342 10122
rect 1366 10051 1437 10122
rect 36085 10051 36156 10122
rect 36180 10051 36251 10122
rect 36289 10051 36360 10122
rect 36384 10051 36455 10122
rect 591 9763 662 9834
rect 686 9763 757 9834
rect 795 9763 866 9834
rect 890 9763 961 9834
rect 36561 9763 36632 9834
rect 36656 9763 36727 9834
rect 36765 9763 36836 9834
rect 36860 9763 36931 9834
rect 37431 10243 37495 10307
rect 37430 10131 37494 10195
rect 41930 10096 42142 10246
rect 37430 10013 37494 10077
rect 41930 9540 42142 9690
rect 1067 9047 1138 9118
rect 1162 9047 1233 9118
rect 1271 9047 1342 9118
rect 1366 9047 1437 9118
rect 36085 9047 36156 9118
rect 36180 9047 36251 9118
rect 36289 9047 36360 9118
rect 36384 9047 36455 9118
rect 591 8759 662 8830
rect 686 8759 757 8830
rect 795 8759 866 8830
rect 890 8759 961 8830
rect 36561 8759 36632 8830
rect 36656 8759 36727 8830
rect 36765 8759 36836 8830
rect 36860 8759 36931 8830
rect 36094 8437 36158 8501
rect 36190 8437 36254 8501
rect 36286 8437 36350 8501
rect 36382 8437 36446 8501
rect 36094 8346 36158 8410
rect 36190 8346 36254 8410
rect 36286 8346 36350 8410
rect 36382 8346 36446 8410
rect 36094 8255 36158 8319
rect 36190 8255 36254 8319
rect 36286 8255 36350 8319
rect 36382 8255 36446 8319
rect 42422 9080 42634 9492
rect 37427 8439 37483 8495
rect 37427 8348 37483 8404
rect 42410 8384 42648 8546
rect 37427 8257 37483 8313
rect 1067 8043 1138 8114
rect 1162 8043 1233 8114
rect 1271 8043 1342 8114
rect 1366 8043 1437 8114
rect 36085 8043 36156 8114
rect 36180 8043 36251 8114
rect 36289 8043 36360 8114
rect 36384 8043 36455 8114
rect 591 7755 662 7826
rect 686 7755 757 7826
rect 795 7755 866 7826
rect 890 7755 961 7826
rect 36561 7755 36632 7826
rect 36656 7755 36727 7826
rect 36765 7755 36836 7826
rect 36860 7755 36931 7826
rect 1067 7039 1138 7110
rect 1162 7039 1233 7110
rect 1271 7039 1342 7110
rect 1366 7039 1437 7110
rect 36085 7039 36156 7110
rect 36180 7039 36251 7110
rect 36289 7039 36360 7110
rect 36384 7039 36455 7110
rect 591 6751 662 6822
rect 686 6751 757 6822
rect 795 6751 866 6822
rect 890 6751 961 6822
rect 36561 6751 36632 6822
rect 36656 6751 36727 6822
rect 36765 6751 36836 6822
rect 36860 6751 36931 6822
rect 42410 7494 42648 7656
rect 42422 6838 42634 7250
rect 41930 6638 42142 6788
rect 1067 6035 1138 6106
rect 1162 6035 1233 6106
rect 1271 6035 1342 6106
rect 1366 6035 1437 6106
rect 36085 6035 36156 6106
rect 36180 6035 36251 6106
rect 36289 6035 36360 6106
rect 36384 6035 36455 6106
rect 591 5747 662 5818
rect 686 5747 757 5818
rect 795 5747 866 5818
rect 890 5747 961 5818
rect 36561 5747 36632 5818
rect 36656 5747 36727 5818
rect 36765 5747 36836 5818
rect 36860 5747 36931 5818
rect 37431 6241 37495 6305
rect 37430 6129 37494 6193
rect 41930 6096 42142 6246
rect 37430 6011 37494 6075
rect 41930 5540 42142 5690
rect 1067 5031 1138 5102
rect 1162 5031 1233 5102
rect 1271 5031 1342 5102
rect 1366 5031 1437 5102
rect 36085 5031 36156 5102
rect 36180 5031 36251 5102
rect 36289 5031 36360 5102
rect 36384 5031 36455 5102
rect 591 4743 662 4814
rect 686 4743 757 4814
rect 795 4743 866 4814
rect 890 4743 961 4814
rect 36561 4743 36632 4814
rect 36656 4743 36727 4814
rect 36765 4743 36836 4814
rect 36860 4743 36931 4814
rect 1067 4027 1138 4098
rect 1162 4027 1233 4098
rect 1271 4027 1342 4098
rect 1366 4027 1437 4098
rect 36085 4027 36156 4098
rect 36180 4027 36251 4098
rect 36289 4027 36360 4098
rect 36384 4027 36455 4098
rect 591 3739 662 3810
rect 686 3739 757 3810
rect 795 3739 866 3810
rect 890 3739 961 3810
rect 36561 3739 36632 3810
rect 36656 3739 36727 3810
rect 36765 3739 36836 3810
rect 36860 3739 36931 3810
rect 36094 3525 36158 3589
rect 36190 3525 36254 3589
rect 36286 3525 36350 3589
rect 36382 3525 36446 3589
rect 36094 3434 36158 3498
rect 36190 3434 36254 3498
rect 36286 3434 36350 3498
rect 36382 3434 36446 3498
rect 36094 3343 36158 3407
rect 36190 3343 36254 3407
rect 36286 3343 36350 3407
rect 36382 3343 36446 3407
rect 42422 5080 42634 5492
rect 42410 4384 42648 4546
rect 37427 3527 37483 3583
rect 37427 3436 37483 3492
rect 42410 3494 42648 3656
rect 37427 3345 37483 3401
rect 1067 3021 1138 3092
rect 1162 3021 1233 3092
rect 1271 3021 1342 3092
rect 1366 3021 1437 3092
rect 36085 3023 36156 3094
rect 36180 3023 36251 3094
rect 36289 3023 36360 3094
rect 36384 3023 36455 3094
rect 591 2735 662 2806
rect 686 2735 757 2806
rect 795 2735 866 2806
rect 890 2735 961 2806
rect 36561 2735 36632 2806
rect 36656 2735 36727 2806
rect 36765 2735 36836 2806
rect 36860 2735 36931 2806
rect 42422 2838 42634 3250
rect 41930 2638 42142 2788
rect 1067 2018 1138 2089
rect 1162 2018 1233 2089
rect 1271 2018 1342 2089
rect 1366 2018 1437 2089
rect 36085 2019 36156 2090
rect 36180 2019 36251 2090
rect 36289 2019 36360 2090
rect 36384 2019 36455 2090
rect 591 1677 662 1748
rect 686 1677 757 1748
rect 795 1677 866 1748
rect 890 1677 961 1748
rect 36561 1731 36632 1802
rect 36656 1731 36727 1802
rect 36765 1731 36836 1802
rect 36860 1731 36931 1802
rect 1067 1363 1138 1434
rect 1162 1363 1233 1434
rect 1271 1363 1342 1434
rect 1366 1363 1437 1434
rect 1067 1253 1138 1324
rect 1162 1253 1233 1324
rect 1271 1253 1342 1324
rect 1366 1253 1437 1324
rect 37431 2247 37495 2311
rect 37430 2135 37494 2199
rect 41930 2096 42142 2246
rect 37430 2017 37494 2081
rect 41930 1540 42142 1690
rect 1067 1014 1138 1085
rect 1162 1014 1233 1085
rect 1271 1014 1342 1085
rect 1366 1014 1437 1085
rect 36085 1015 36156 1086
rect 36180 1015 36251 1086
rect 36289 1015 36360 1086
rect 36384 1015 36455 1086
rect 591 741 662 812
rect 686 741 757 812
rect 795 741 866 812
rect 890 741 961 812
rect 36094 817 36158 881
rect 36190 817 36254 881
rect 36286 817 36350 881
rect 36382 817 36446 881
rect 36094 726 36158 790
rect 36190 726 36254 790
rect 36286 726 36350 790
rect 36382 726 36446 790
rect 36094 635 36158 699
rect 36190 635 36254 699
rect 36286 635 36350 699
rect 36382 635 36446 699
rect 36561 455 36632 526
rect 36656 455 36727 526
rect 36765 455 36836 526
rect 36860 455 36931 526
rect 42422 1080 42634 1492
rect 37427 819 37483 875
rect 37427 728 37483 784
rect 37427 637 37483 693
rect 42410 384 42648 546
<< metal3 >>
rect 41684 23656 42660 23668
rect 41684 23655 42410 23656
rect 41684 23498 41707 23655
rect 41821 23498 42410 23655
rect 41684 23494 42410 23498
rect 42648 23494 42660 23656
rect 41684 23484 42660 23494
rect 42396 23250 42660 23276
rect 42396 22838 42422 23250
rect 42634 22838 42660 23250
rect 42396 22814 42660 22838
rect 41602 22788 42164 22806
rect 41602 22638 41930 22788
rect 42142 22638 42164 22788
rect 41602 22624 42164 22638
rect 41602 22246 42164 22264
rect 41602 22096 41930 22246
rect 42142 22096 42164 22246
rect 41602 22082 42164 22096
rect 41602 21690 42164 21708
rect 41602 21540 41930 21690
rect 42142 21540 42164 21690
rect 41602 21526 42164 21540
rect 42396 21492 42660 21518
rect 42396 21080 42422 21492
rect 42634 21080 42660 21492
rect 42396 21056 42660 21080
rect 41684 20546 42660 20558
rect 41684 20545 42410 20546
rect 41684 20388 41707 20545
rect 41821 20388 42410 20545
rect 41684 20384 42410 20388
rect 42648 20384 42660 20546
rect 41684 20374 42660 20384
rect 2284 20167 2482 20168
rect 1884 20104 2176 20167
rect 1884 19946 1898 20104
rect 2160 19946 2176 20104
rect 570 19889 984 19900
rect 570 19634 587 19889
rect 969 19634 984 19889
rect 570 19620 984 19634
rect 1046 19620 1460 19900
rect 1046 19451 1460 19462
rect 1046 19196 1063 19451
rect 1445 19196 1460 19451
rect 1046 19182 1460 19196
rect 1884 19442 2176 19946
rect 5012 20104 5304 20166
rect 5012 19946 5026 20104
rect 5288 19946 5304 20104
rect 3420 19882 3790 19900
rect 3420 19638 3444 19882
rect 3770 19638 3790 19882
rect 3420 19620 3790 19638
rect 1884 19386 1904 19442
rect 1960 19386 1998 19442
rect 2054 19386 2092 19442
rect 2148 19386 2176 19442
rect 1884 19348 2176 19386
rect 1884 19292 1904 19348
rect 1960 19292 1998 19348
rect 2054 19292 2092 19348
rect 2148 19292 2176 19348
rect 1884 19254 2176 19292
rect 1884 19198 1904 19254
rect 1960 19198 1998 19254
rect 2054 19198 2092 19254
rect 2148 19198 2176 19254
rect 1884 19182 2176 19198
rect 5012 19442 5304 19946
rect 5012 19386 5032 19442
rect 5088 19386 5126 19442
rect 5182 19386 5220 19442
rect 5276 19386 5304 19442
rect 5012 19348 5304 19386
rect 5012 19292 5032 19348
rect 5088 19292 5126 19348
rect 5182 19292 5220 19348
rect 5276 19292 5304 19348
rect 5012 19254 5304 19292
rect 5012 19198 5032 19254
rect 5088 19198 5126 19254
rect 5182 19198 5220 19254
rect 5276 19198 5304 19254
rect 5012 19182 5304 19198
rect 5884 20104 6176 20166
rect 5884 19946 5898 20104
rect 6160 19946 6176 20104
rect 5884 19442 6176 19946
rect 9012 20104 9304 20166
rect 9012 19946 9026 20104
rect 9288 19946 9304 20104
rect 7420 19882 7790 19900
rect 7420 19638 7444 19882
rect 7770 19638 7790 19882
rect 7420 19620 7790 19638
rect 5884 19386 5904 19442
rect 5960 19386 5998 19442
rect 6054 19386 6092 19442
rect 6148 19386 6176 19442
rect 5884 19348 6176 19386
rect 5884 19292 5904 19348
rect 5960 19292 5998 19348
rect 6054 19292 6092 19348
rect 6148 19292 6176 19348
rect 5884 19254 6176 19292
rect 5884 19198 5904 19254
rect 5960 19198 5998 19254
rect 6054 19198 6092 19254
rect 6148 19198 6176 19254
rect 5884 19182 6176 19198
rect 9012 19442 9304 19946
rect 9012 19386 9032 19442
rect 9088 19386 9126 19442
rect 9182 19386 9220 19442
rect 9276 19386 9304 19442
rect 9012 19348 9304 19386
rect 9012 19292 9032 19348
rect 9088 19292 9126 19348
rect 9182 19292 9220 19348
rect 9276 19292 9304 19348
rect 9012 19254 9304 19292
rect 9012 19198 9032 19254
rect 9088 19198 9126 19254
rect 9182 19198 9220 19254
rect 9276 19198 9304 19254
rect 9012 19182 9304 19198
rect 9884 20104 10176 20166
rect 9884 19946 9898 20104
rect 10160 19946 10176 20104
rect 9884 19442 10176 19946
rect 13012 20104 13304 20166
rect 13012 19946 13026 20104
rect 13288 19946 13304 20104
rect 11420 19882 11790 19900
rect 11420 19638 11444 19882
rect 11770 19638 11790 19882
rect 11420 19620 11790 19638
rect 9884 19386 9904 19442
rect 9960 19386 9998 19442
rect 10054 19386 10092 19442
rect 10148 19386 10176 19442
rect 9884 19348 10176 19386
rect 9884 19292 9904 19348
rect 9960 19292 9998 19348
rect 10054 19292 10092 19348
rect 10148 19292 10176 19348
rect 9884 19254 10176 19292
rect 9884 19198 9904 19254
rect 9960 19198 9998 19254
rect 10054 19198 10092 19254
rect 10148 19198 10176 19254
rect 9884 19182 10176 19198
rect 13012 19442 13304 19946
rect 13012 19386 13032 19442
rect 13088 19386 13126 19442
rect 13182 19386 13220 19442
rect 13276 19386 13304 19442
rect 13012 19348 13304 19386
rect 13012 19292 13032 19348
rect 13088 19292 13126 19348
rect 13182 19292 13220 19348
rect 13276 19292 13304 19348
rect 13012 19254 13304 19292
rect 13012 19198 13032 19254
rect 13088 19198 13126 19254
rect 13182 19198 13220 19254
rect 13276 19198 13304 19254
rect 13012 19182 13304 19198
rect 13884 20104 14176 20166
rect 13884 19946 13898 20104
rect 14160 19946 14176 20104
rect 13884 19442 14176 19946
rect 17012 20104 17304 20166
rect 17012 19946 17026 20104
rect 17288 19946 17304 20104
rect 15420 19882 15790 19900
rect 15420 19638 15444 19882
rect 15770 19638 15790 19882
rect 15420 19620 15790 19638
rect 13884 19386 13904 19442
rect 13960 19386 13998 19442
rect 14054 19386 14092 19442
rect 14148 19386 14176 19442
rect 13884 19348 14176 19386
rect 13884 19292 13904 19348
rect 13960 19292 13998 19348
rect 14054 19292 14092 19348
rect 14148 19292 14176 19348
rect 13884 19254 14176 19292
rect 13884 19198 13904 19254
rect 13960 19198 13998 19254
rect 14054 19198 14092 19254
rect 14148 19198 14176 19254
rect 13884 19182 14176 19198
rect 17012 19442 17304 19946
rect 17012 19386 17032 19442
rect 17088 19386 17126 19442
rect 17182 19386 17220 19442
rect 17276 19386 17304 19442
rect 17012 19348 17304 19386
rect 17012 19292 17032 19348
rect 17088 19292 17126 19348
rect 17182 19292 17220 19348
rect 17276 19292 17304 19348
rect 17012 19254 17304 19292
rect 17012 19198 17032 19254
rect 17088 19198 17126 19254
rect 17182 19198 17220 19254
rect 17276 19198 17304 19254
rect 17012 19182 17304 19198
rect 17884 20104 18176 20166
rect 17884 19946 17898 20104
rect 18160 19946 18176 20104
rect 17884 19442 18176 19946
rect 21012 20104 21304 20166
rect 21012 19946 21026 20104
rect 21288 19946 21304 20104
rect 19420 19882 19790 19900
rect 19420 19638 19444 19882
rect 19770 19638 19790 19882
rect 19420 19620 19790 19638
rect 17884 19386 17904 19442
rect 17960 19386 17998 19442
rect 18054 19386 18092 19442
rect 18148 19386 18176 19442
rect 17884 19348 18176 19386
rect 17884 19292 17904 19348
rect 17960 19292 17998 19348
rect 18054 19292 18092 19348
rect 18148 19292 18176 19348
rect 17884 19254 18176 19292
rect 17884 19198 17904 19254
rect 17960 19198 17998 19254
rect 18054 19198 18092 19254
rect 18148 19198 18176 19254
rect 17884 19182 18176 19198
rect 21012 19442 21304 19946
rect 21012 19386 21032 19442
rect 21088 19386 21126 19442
rect 21182 19386 21220 19442
rect 21276 19386 21304 19442
rect 21012 19348 21304 19386
rect 21012 19292 21032 19348
rect 21088 19292 21126 19348
rect 21182 19292 21220 19348
rect 21276 19292 21304 19348
rect 21012 19254 21304 19292
rect 21012 19198 21032 19254
rect 21088 19198 21126 19254
rect 21182 19198 21220 19254
rect 21276 19198 21304 19254
rect 21012 19182 21304 19198
rect 21884 20104 22176 20166
rect 21884 19946 21898 20104
rect 22160 19946 22176 20104
rect 21884 19442 22176 19946
rect 25012 20104 25304 20166
rect 25012 19946 25026 20104
rect 25288 19946 25304 20104
rect 23420 19882 23790 19900
rect 23420 19638 23444 19882
rect 23770 19638 23790 19882
rect 23420 19620 23790 19638
rect 21884 19386 21904 19442
rect 21960 19386 21998 19442
rect 22054 19386 22092 19442
rect 22148 19386 22176 19442
rect 21884 19348 22176 19386
rect 21884 19292 21904 19348
rect 21960 19292 21998 19348
rect 22054 19292 22092 19348
rect 22148 19292 22176 19348
rect 21884 19254 22176 19292
rect 21884 19198 21904 19254
rect 21960 19198 21998 19254
rect 22054 19198 22092 19254
rect 22148 19198 22176 19254
rect 21884 19182 22176 19198
rect 25012 19442 25304 19946
rect 25012 19386 25032 19442
rect 25088 19386 25126 19442
rect 25182 19386 25220 19442
rect 25276 19386 25304 19442
rect 25012 19348 25304 19386
rect 25012 19292 25032 19348
rect 25088 19292 25126 19348
rect 25182 19292 25220 19348
rect 25276 19292 25304 19348
rect 25012 19254 25304 19292
rect 25012 19198 25032 19254
rect 25088 19198 25126 19254
rect 25182 19198 25220 19254
rect 25276 19198 25304 19254
rect 25012 19182 25304 19198
rect 25884 20104 26176 20166
rect 25884 19946 25898 20104
rect 26160 19946 26176 20104
rect 25884 19442 26176 19946
rect 29012 20104 29304 20166
rect 29012 19946 29026 20104
rect 29288 19946 29304 20104
rect 27420 19882 27790 19900
rect 27420 19638 27444 19882
rect 27770 19638 27790 19882
rect 27420 19620 27790 19638
rect 25884 19386 25904 19442
rect 25960 19386 25998 19442
rect 26054 19386 26092 19442
rect 26148 19386 26176 19442
rect 25884 19348 26176 19386
rect 25884 19292 25904 19348
rect 25960 19292 25998 19348
rect 26054 19292 26092 19348
rect 26148 19292 26176 19348
rect 25884 19254 26176 19292
rect 25884 19198 25904 19254
rect 25960 19198 25998 19254
rect 26054 19198 26092 19254
rect 26148 19198 26176 19254
rect 25884 19182 26176 19198
rect 29012 19442 29304 19946
rect 29012 19386 29032 19442
rect 29088 19386 29126 19442
rect 29182 19386 29220 19442
rect 29276 19386 29304 19442
rect 29012 19348 29304 19386
rect 29012 19292 29032 19348
rect 29088 19292 29126 19348
rect 29182 19292 29220 19348
rect 29276 19292 29304 19348
rect 29012 19254 29304 19292
rect 29012 19198 29032 19254
rect 29088 19198 29126 19254
rect 29182 19198 29220 19254
rect 29276 19198 29304 19254
rect 29012 19182 29304 19198
rect 29884 20104 30176 20166
rect 29884 19946 29898 20104
rect 30160 19946 30176 20104
rect 29884 19442 30176 19946
rect 33012 20104 33304 20166
rect 33012 19946 33026 20104
rect 33288 19946 33304 20104
rect 31420 19882 31790 19900
rect 31420 19638 31444 19882
rect 31770 19638 31790 19882
rect 31420 19620 31790 19638
rect 29884 19386 29904 19442
rect 29960 19386 29998 19442
rect 30054 19386 30092 19442
rect 30148 19386 30176 19442
rect 29884 19348 30176 19386
rect 29884 19292 29904 19348
rect 29960 19292 29998 19348
rect 30054 19292 30092 19348
rect 30148 19292 30176 19348
rect 29884 19254 30176 19292
rect 29884 19198 29904 19254
rect 29960 19198 29998 19254
rect 30054 19198 30092 19254
rect 30148 19198 30176 19254
rect 29884 19182 30176 19198
rect 33012 19442 33304 19946
rect 33012 19386 33032 19442
rect 33088 19386 33126 19442
rect 33182 19386 33220 19442
rect 33276 19386 33304 19442
rect 33012 19348 33304 19386
rect 33012 19292 33032 19348
rect 33088 19292 33126 19348
rect 33182 19292 33220 19348
rect 33276 19292 33304 19348
rect 33012 19254 33304 19292
rect 33012 19198 33032 19254
rect 33088 19198 33126 19254
rect 33182 19198 33220 19254
rect 33276 19198 33304 19254
rect 33012 19182 33304 19198
rect 33884 20104 34176 20166
rect 33884 19946 33898 20104
rect 34160 19946 34176 20104
rect 37012 20104 37304 20166
rect 37012 19980 37026 20104
rect 37288 19980 37304 20104
rect 37012 19968 37304 19980
rect 33884 19442 34176 19946
rect 36540 19885 36954 19900
rect 35396 19847 35810 19862
rect 35396 19783 35426 19847
rect 35490 19783 35522 19847
rect 35586 19783 35618 19847
rect 35682 19783 35714 19847
rect 35778 19783 35810 19847
rect 35396 19753 35810 19783
rect 35396 19689 35426 19753
rect 35490 19689 35522 19753
rect 35586 19689 35618 19753
rect 35682 19689 35714 19753
rect 35778 19689 35810 19753
rect 36540 19821 36570 19885
rect 36634 19821 36666 19885
rect 36730 19821 36762 19885
rect 36826 19821 36858 19885
rect 36922 19821 36954 19885
rect 36540 19791 36954 19821
rect 36540 19727 36570 19791
rect 36634 19727 36666 19791
rect 36730 19727 36762 19791
rect 36826 19727 36858 19791
rect 36922 19727 36954 19791
rect 36540 19692 36954 19727
rect 35396 19655 35810 19689
rect 41684 19656 42660 19668
rect 41684 19655 42410 19656
rect 33884 19386 33904 19442
rect 33960 19386 33998 19442
rect 34054 19386 34092 19442
rect 34148 19386 34176 19442
rect 33884 19348 34176 19386
rect 33884 19292 33904 19348
rect 33960 19292 33998 19348
rect 34054 19292 34092 19348
rect 34148 19292 34176 19348
rect 33884 19254 34176 19292
rect 33884 19198 33904 19254
rect 33960 19198 33998 19254
rect 34054 19198 34092 19254
rect 34148 19198 34176 19254
rect 33884 19182 34176 19198
rect 36064 19557 37512 19585
rect 36064 19493 36094 19557
rect 36158 19493 36190 19557
rect 36254 19493 36286 19557
rect 36350 19493 36382 19557
rect 36446 19555 37512 19557
rect 36446 19493 37423 19555
rect 36064 19491 37423 19493
rect 37487 19491 37512 19555
rect 36064 19466 37512 19491
rect 41684 19498 41707 19655
rect 41821 19498 42410 19655
rect 41684 19494 42410 19498
rect 42648 19494 42660 19656
rect 41684 19484 42660 19494
rect 36064 19402 36094 19466
rect 36158 19402 36190 19466
rect 36254 19402 36286 19466
rect 36350 19402 36382 19466
rect 36446 19463 37512 19466
rect 36446 19402 37423 19463
rect 36064 19399 37423 19402
rect 37487 19399 37512 19463
rect 36064 19375 37512 19399
rect 36064 19311 36094 19375
rect 36158 19311 36190 19375
rect 36254 19311 36286 19375
rect 36350 19311 36382 19375
rect 36446 19372 37512 19375
rect 36446 19311 37423 19372
rect 36064 19308 37423 19311
rect 37487 19308 37512 19372
rect 36064 19286 37512 19308
rect 36064 19281 36478 19286
rect 36064 19217 36094 19281
rect 36158 19217 36190 19281
rect 36254 19217 36286 19281
rect 36350 19217 36382 19281
rect 36446 19217 36478 19281
rect 36064 19182 36478 19217
rect 42396 19250 42660 19276
rect 36540 18870 36954 18890
rect 570 18816 984 18836
rect 570 18745 591 18816
rect 662 18745 686 18816
rect 757 18745 795 18816
rect 866 18745 890 18816
rect 961 18745 984 18816
rect 36540 18799 36561 18870
rect 36632 18799 36656 18870
rect 36727 18799 36765 18870
rect 36836 18799 36860 18870
rect 36931 18799 36954 18870
rect 42396 18838 42422 19250
rect 42634 18838 42660 19250
rect 42396 18814 42660 18838
rect 36540 18780 36954 18799
rect 41602 18788 42164 18806
rect 570 18726 984 18745
rect 41602 18638 41930 18788
rect 42142 18638 42164 18788
rect 41602 18624 42164 18638
rect 570 18502 984 18522
rect 570 18431 591 18502
rect 662 18431 686 18502
rect 757 18431 795 18502
rect 866 18431 890 18502
rect 961 18431 984 18502
rect 570 18412 984 18431
rect 1046 18363 1460 18383
rect 1046 18292 1067 18363
rect 1138 18292 1162 18363
rect 1233 18292 1271 18363
rect 1342 18292 1366 18363
rect 1437 18292 1460 18363
rect 1046 18273 1460 18292
rect 37392 18307 37542 18332
rect 37392 18243 37431 18307
rect 37495 18243 37542 18307
rect 37392 18195 37542 18243
rect 1046 18153 1460 18173
rect 1046 18082 1067 18153
rect 1138 18082 1162 18153
rect 1233 18082 1271 18153
rect 1342 18082 1366 18153
rect 1437 18082 1460 18153
rect 1046 18063 1460 18082
rect 36064 18154 36478 18174
rect 36064 18083 36085 18154
rect 36156 18083 36180 18154
rect 36251 18083 36289 18154
rect 36360 18083 36384 18154
rect 36455 18083 36478 18154
rect 36064 18064 36478 18083
rect 37392 18131 37430 18195
rect 37494 18131 37542 18195
rect 37392 18077 37542 18131
rect 41602 18246 42164 18264
rect 41602 18096 41930 18246
rect 42142 18096 42164 18246
rect 41602 18082 42164 18096
rect 37392 18013 37430 18077
rect 37494 18013 37542 18077
rect 37392 17988 37542 18013
rect 570 17866 984 17886
rect 570 17795 591 17866
rect 662 17795 686 17866
rect 757 17795 795 17866
rect 866 17795 890 17866
rect 961 17795 984 17866
rect 570 17776 984 17795
rect 36540 17866 36954 17886
rect 36540 17795 36561 17866
rect 36632 17795 36656 17866
rect 36727 17795 36765 17866
rect 36836 17795 36860 17866
rect 36931 17795 36954 17866
rect 36540 17776 36954 17795
rect 41602 17690 42164 17708
rect 41602 17540 41930 17690
rect 42142 17540 42164 17690
rect 41602 17526 42164 17540
rect 42396 17492 42660 17518
rect 1046 17150 1460 17170
rect 1046 17079 1067 17150
rect 1138 17079 1162 17150
rect 1233 17079 1271 17150
rect 1342 17079 1366 17150
rect 1437 17079 1460 17150
rect 1046 17060 1460 17079
rect 36064 17150 36478 17170
rect 36064 17079 36085 17150
rect 36156 17079 36180 17150
rect 36251 17079 36289 17150
rect 36360 17079 36384 17150
rect 36455 17079 36478 17150
rect 36064 17060 36478 17079
rect 42396 17080 42422 17492
rect 42634 17080 42660 17492
rect 42396 17056 42660 17080
rect 570 16862 984 16882
rect 570 16791 591 16862
rect 662 16791 686 16862
rect 757 16791 795 16862
rect 866 16791 890 16862
rect 961 16791 984 16862
rect 570 16772 984 16791
rect 36540 16862 36954 16882
rect 36540 16791 36561 16862
rect 36632 16791 36656 16862
rect 36727 16791 36765 16862
rect 36836 16791 36860 16862
rect 36931 16791 36954 16862
rect 36540 16772 36954 16791
rect 36064 16652 37512 16680
rect 36064 16588 36094 16652
rect 36158 16588 36190 16652
rect 36254 16588 36286 16652
rect 36350 16588 36382 16652
rect 36446 16650 37512 16652
rect 36446 16588 37423 16650
rect 36064 16586 37423 16588
rect 37487 16586 37512 16650
rect 36064 16561 37512 16586
rect 36064 16497 36094 16561
rect 36158 16497 36190 16561
rect 36254 16497 36286 16561
rect 36350 16497 36382 16561
rect 36446 16558 37512 16561
rect 36446 16497 37423 16558
rect 36064 16494 37423 16497
rect 37487 16494 37512 16558
rect 36064 16470 37512 16494
rect 36064 16406 36094 16470
rect 36158 16406 36190 16470
rect 36254 16406 36286 16470
rect 36350 16406 36382 16470
rect 36446 16467 37512 16470
rect 36446 16406 37423 16467
rect 36064 16403 37423 16406
rect 37487 16403 37512 16467
rect 36064 16381 37512 16403
rect 41684 16546 42660 16558
rect 41684 16545 42410 16546
rect 41684 16388 41707 16545
rect 41821 16388 42410 16545
rect 41684 16384 42410 16388
rect 42648 16384 42660 16546
rect 41684 16374 42660 16384
rect 1046 16145 1460 16165
rect 1046 16074 1067 16145
rect 1138 16074 1162 16145
rect 1233 16074 1271 16145
rect 1342 16074 1366 16145
rect 1437 16074 1460 16145
rect 1046 16055 1460 16074
rect 36064 16146 36478 16166
rect 36064 16075 36085 16146
rect 36156 16075 36180 16146
rect 36251 16075 36289 16146
rect 36360 16075 36384 16146
rect 36455 16075 36478 16146
rect 36064 16056 36478 16075
rect 570 15858 984 15878
rect 570 15787 591 15858
rect 662 15787 686 15858
rect 757 15787 795 15858
rect 866 15787 890 15858
rect 961 15787 984 15858
rect 570 15768 984 15787
rect 36540 15858 36954 15878
rect 36540 15787 36561 15858
rect 36632 15787 36656 15858
rect 36727 15787 36765 15858
rect 36836 15787 36860 15858
rect 36931 15787 36954 15858
rect 36540 15768 36954 15787
rect 41684 15656 42660 15668
rect 41684 15655 42410 15656
rect 41684 15498 41707 15655
rect 41821 15498 42410 15655
rect 41684 15494 42410 15498
rect 42648 15494 42660 15656
rect 41684 15484 42660 15494
rect 42396 15250 42660 15276
rect 1046 15142 1460 15162
rect 1046 15071 1067 15142
rect 1138 15071 1162 15142
rect 1233 15071 1271 15142
rect 1342 15071 1366 15142
rect 1437 15071 1460 15142
rect 1046 15052 1460 15071
rect 36064 15142 36478 15162
rect 36064 15071 36085 15142
rect 36156 15071 36180 15142
rect 36251 15071 36289 15142
rect 36360 15071 36384 15142
rect 36455 15071 36478 15142
rect 36064 15052 36478 15071
rect 570 14854 984 14874
rect 570 14783 591 14854
rect 662 14783 686 14854
rect 757 14783 795 14854
rect 866 14783 890 14854
rect 961 14783 984 14854
rect 570 14764 984 14783
rect 36540 14854 36954 14874
rect 36540 14783 36561 14854
rect 36632 14783 36656 14854
rect 36727 14783 36765 14854
rect 36836 14783 36860 14854
rect 36931 14783 36954 14854
rect 42396 14838 42422 15250
rect 42634 14838 42660 15250
rect 42396 14814 42660 14838
rect 36540 14764 36954 14783
rect 41602 14788 42164 14806
rect 41602 14638 41930 14788
rect 42142 14638 42164 14788
rect 41602 14624 42164 14638
rect 37392 14307 37542 14332
rect 37392 14243 37431 14307
rect 37495 14243 37542 14307
rect 37392 14195 37542 14243
rect 1046 14138 1460 14158
rect 1046 14067 1067 14138
rect 1138 14067 1162 14138
rect 1233 14067 1271 14138
rect 1342 14067 1366 14138
rect 1437 14067 1460 14138
rect 1046 14048 1460 14067
rect 36064 14138 36478 14158
rect 36064 14067 36085 14138
rect 36156 14067 36180 14138
rect 36251 14067 36289 14138
rect 36360 14067 36384 14138
rect 36455 14067 36478 14138
rect 36064 14048 36478 14067
rect 37392 14131 37430 14195
rect 37494 14131 37542 14195
rect 37392 14077 37542 14131
rect 41602 14246 42164 14264
rect 41602 14096 41930 14246
rect 42142 14096 42164 14246
rect 41602 14082 42164 14096
rect 37392 14013 37430 14077
rect 37494 14013 37542 14077
rect 37392 13988 37542 14013
rect 570 13850 984 13870
rect 570 13779 591 13850
rect 662 13779 686 13850
rect 757 13779 795 13850
rect 866 13779 890 13850
rect 961 13779 984 13850
rect 570 13760 984 13779
rect 36540 13850 36954 13870
rect 36540 13779 36561 13850
rect 36632 13779 36656 13850
rect 36727 13779 36765 13850
rect 36836 13779 36860 13850
rect 36931 13779 36954 13850
rect 36540 13760 36954 13779
rect 41602 13690 42164 13708
rect 41602 13540 41930 13690
rect 42142 13540 42164 13690
rect 41602 13526 42164 13540
rect 42396 13492 42660 13518
rect 1046 13134 1460 13154
rect 1046 13063 1067 13134
rect 1138 13063 1162 13134
rect 1233 13063 1271 13134
rect 1342 13063 1366 13134
rect 1437 13063 1460 13134
rect 1046 13044 1460 13063
rect 36064 13134 36478 13154
rect 36064 13063 36085 13134
rect 36156 13063 36180 13134
rect 36251 13063 36289 13134
rect 36360 13063 36384 13134
rect 36455 13063 36478 13134
rect 36064 13044 36478 13063
rect 42396 13080 42422 13492
rect 42634 13080 42660 13492
rect 42396 13056 42660 13080
rect 570 12846 984 12866
rect 570 12775 591 12846
rect 662 12775 686 12846
rect 757 12775 795 12846
rect 866 12775 890 12846
rect 961 12775 984 12846
rect 570 12756 984 12775
rect 36540 12846 36954 12866
rect 36540 12775 36561 12846
rect 36632 12775 36656 12846
rect 36727 12775 36765 12846
rect 36836 12775 36860 12846
rect 36931 12775 36954 12846
rect 36540 12756 36954 12775
rect 36064 12594 37512 12622
rect 36064 12530 36094 12594
rect 36158 12530 36190 12594
rect 36254 12530 36286 12594
rect 36350 12530 36382 12594
rect 36446 12592 37512 12594
rect 36446 12530 37423 12592
rect 36064 12528 37423 12530
rect 37487 12528 37512 12592
rect 36064 12503 37512 12528
rect 36064 12439 36094 12503
rect 36158 12439 36190 12503
rect 36254 12439 36286 12503
rect 36350 12439 36382 12503
rect 36446 12500 37512 12503
rect 36446 12439 37423 12500
rect 36064 12436 37423 12439
rect 37487 12436 37512 12500
rect 36064 12412 37512 12436
rect 36064 12348 36094 12412
rect 36158 12348 36190 12412
rect 36254 12348 36286 12412
rect 36350 12348 36382 12412
rect 36446 12409 37512 12412
rect 36446 12348 37423 12409
rect 36064 12345 37423 12348
rect 37487 12345 37512 12409
rect 41684 12546 42660 12558
rect 41684 12545 42410 12546
rect 41684 12388 41707 12545
rect 41821 12388 42410 12545
rect 41684 12384 42410 12388
rect 42648 12384 42660 12546
rect 41684 12374 42660 12384
rect 36064 12323 37512 12345
rect 1046 12130 1460 12150
rect 1046 12059 1067 12130
rect 1138 12059 1162 12130
rect 1233 12059 1271 12130
rect 1342 12059 1366 12130
rect 1437 12059 1460 12130
rect 1046 12040 1460 12059
rect 36064 12130 36478 12150
rect 36064 12059 36085 12130
rect 36156 12059 36180 12130
rect 36251 12059 36289 12130
rect 36360 12059 36384 12130
rect 36455 12059 36478 12130
rect 36064 12040 36478 12059
rect 570 11842 984 11862
rect 570 11771 591 11842
rect 662 11771 686 11842
rect 757 11771 795 11842
rect 866 11771 890 11842
rect 961 11771 984 11842
rect 570 11752 984 11771
rect 36540 11842 36954 11862
rect 36540 11771 36561 11842
rect 36632 11771 36656 11842
rect 36727 11771 36765 11842
rect 36836 11771 36860 11842
rect 36931 11771 36954 11842
rect 36540 11752 36954 11771
rect 41684 11656 42660 11668
rect 41684 11655 42410 11656
rect 41684 11498 41707 11655
rect 41821 11498 42410 11655
rect 41684 11494 42410 11498
rect 42648 11494 42660 11656
rect 41684 11484 42660 11494
rect 42396 11250 42660 11276
rect 1046 11126 1460 11146
rect 1046 11055 1067 11126
rect 1138 11055 1162 11126
rect 1233 11055 1271 11126
rect 1342 11055 1366 11126
rect 1437 11055 1460 11126
rect 1046 11036 1460 11055
rect 36064 11126 36478 11146
rect 36064 11055 36085 11126
rect 36156 11055 36180 11126
rect 36251 11055 36289 11126
rect 36360 11055 36384 11126
rect 36455 11055 36478 11126
rect 36064 11036 36478 11055
rect 570 10838 984 10858
rect 570 10767 591 10838
rect 662 10767 686 10838
rect 757 10767 795 10838
rect 866 10767 890 10838
rect 961 10767 984 10838
rect 570 10748 984 10767
rect 36540 10838 36954 10858
rect 36540 10767 36561 10838
rect 36632 10767 36656 10838
rect 36727 10767 36765 10838
rect 36836 10767 36860 10838
rect 36931 10767 36954 10838
rect 42396 10838 42422 11250
rect 42634 10838 42660 11250
rect 42396 10814 42660 10838
rect 36540 10748 36954 10767
rect 41602 10788 42164 10806
rect 41602 10638 41930 10788
rect 42142 10638 42164 10788
rect 41602 10624 42164 10638
rect 37392 10307 37542 10332
rect 37392 10243 37431 10307
rect 37495 10243 37542 10307
rect 37392 10195 37542 10243
rect 1046 10122 1460 10142
rect 1046 10051 1067 10122
rect 1138 10051 1162 10122
rect 1233 10051 1271 10122
rect 1342 10051 1366 10122
rect 1437 10051 1460 10122
rect 1046 10032 1460 10051
rect 36064 10122 36478 10142
rect 36064 10051 36085 10122
rect 36156 10051 36180 10122
rect 36251 10051 36289 10122
rect 36360 10051 36384 10122
rect 36455 10051 36478 10122
rect 36064 10032 36478 10051
rect 37392 10131 37430 10195
rect 37494 10131 37542 10195
rect 37392 10077 37542 10131
rect 41602 10246 42164 10264
rect 41602 10096 41930 10246
rect 42142 10096 42164 10246
rect 41602 10082 42164 10096
rect 37392 10013 37430 10077
rect 37494 10013 37542 10077
rect 37392 9988 37542 10013
rect 570 9834 984 9854
rect 570 9763 591 9834
rect 662 9763 686 9834
rect 757 9763 795 9834
rect 866 9763 890 9834
rect 961 9763 984 9834
rect 570 9744 984 9763
rect 36540 9834 36954 9854
rect 36540 9763 36561 9834
rect 36632 9763 36656 9834
rect 36727 9763 36765 9834
rect 36836 9763 36860 9834
rect 36931 9763 36954 9834
rect 36540 9744 36954 9763
rect 41602 9690 42164 9708
rect 41602 9540 41930 9690
rect 42142 9540 42164 9690
rect 41602 9526 42164 9540
rect 42396 9492 42660 9518
rect 1046 9118 1460 9138
rect 1046 9047 1067 9118
rect 1138 9047 1162 9118
rect 1233 9047 1271 9118
rect 1342 9047 1366 9118
rect 1437 9047 1460 9118
rect 1046 9028 1460 9047
rect 36064 9118 36478 9138
rect 36064 9047 36085 9118
rect 36156 9047 36180 9118
rect 36251 9047 36289 9118
rect 36360 9047 36384 9118
rect 36455 9047 36478 9118
rect 42396 9080 42422 9492
rect 42634 9080 42660 9492
rect 42396 9056 42660 9080
rect 36064 9028 36478 9047
rect 570 8830 984 8850
rect 570 8759 591 8830
rect 662 8759 686 8830
rect 757 8759 795 8830
rect 866 8759 890 8830
rect 961 8759 984 8830
rect 570 8740 984 8759
rect 36540 8830 36954 8850
rect 36540 8759 36561 8830
rect 36632 8759 36656 8830
rect 36727 8759 36765 8830
rect 36836 8759 36860 8830
rect 36931 8759 36954 8830
rect 36540 8740 36954 8759
rect 41684 8546 42660 8558
rect 41684 8545 42410 8546
rect 36064 8501 37512 8529
rect 36064 8437 36094 8501
rect 36158 8437 36190 8501
rect 36254 8437 36286 8501
rect 36350 8437 36382 8501
rect 36446 8499 37512 8501
rect 36446 8437 37423 8499
rect 36064 8435 37423 8437
rect 37487 8435 37512 8499
rect 36064 8410 37512 8435
rect 36064 8346 36094 8410
rect 36158 8346 36190 8410
rect 36254 8346 36286 8410
rect 36350 8346 36382 8410
rect 36446 8407 37512 8410
rect 36446 8346 37423 8407
rect 36064 8343 37423 8346
rect 37487 8343 37512 8407
rect 41684 8388 41707 8545
rect 41821 8388 42410 8545
rect 41684 8384 42410 8388
rect 42648 8384 42660 8546
rect 41684 8374 42660 8384
rect 36064 8319 37512 8343
rect 36064 8255 36094 8319
rect 36158 8255 36190 8319
rect 36254 8255 36286 8319
rect 36350 8255 36382 8319
rect 36446 8316 37512 8319
rect 36446 8255 37423 8316
rect 36064 8252 37423 8255
rect 37487 8252 37512 8316
rect 36064 8230 37512 8252
rect 1046 8114 1460 8134
rect 1046 8043 1067 8114
rect 1138 8043 1162 8114
rect 1233 8043 1271 8114
rect 1342 8043 1366 8114
rect 1437 8043 1460 8114
rect 1046 8024 1460 8043
rect 36064 8114 36478 8134
rect 36064 8043 36085 8114
rect 36156 8043 36180 8114
rect 36251 8043 36289 8114
rect 36360 8043 36384 8114
rect 36455 8043 36478 8114
rect 36064 8024 36478 8043
rect 570 7826 984 7846
rect 570 7755 591 7826
rect 662 7755 686 7826
rect 757 7755 795 7826
rect 866 7755 890 7826
rect 961 7755 984 7826
rect 570 7736 984 7755
rect 36540 7826 36954 7846
rect 36540 7755 36561 7826
rect 36632 7755 36656 7826
rect 36727 7755 36765 7826
rect 36836 7755 36860 7826
rect 36931 7755 36954 7826
rect 36540 7736 36954 7755
rect 41684 7656 42660 7668
rect 41684 7655 42410 7656
rect 41684 7498 41707 7655
rect 41821 7498 42410 7655
rect 41684 7494 42410 7498
rect 42648 7494 42660 7656
rect 41684 7484 42660 7494
rect 42396 7250 42660 7276
rect 1046 7110 1460 7130
rect 1046 7039 1067 7110
rect 1138 7039 1162 7110
rect 1233 7039 1271 7110
rect 1342 7039 1366 7110
rect 1437 7039 1460 7110
rect 1046 7020 1460 7039
rect 36064 7110 36478 7130
rect 36064 7039 36085 7110
rect 36156 7039 36180 7110
rect 36251 7039 36289 7110
rect 36360 7039 36384 7110
rect 36455 7039 36478 7110
rect 36064 7020 36478 7039
rect 570 6822 984 6842
rect 570 6751 591 6822
rect 662 6751 686 6822
rect 757 6751 795 6822
rect 866 6751 890 6822
rect 961 6751 984 6822
rect 570 6732 984 6751
rect 36540 6822 36954 6842
rect 36540 6751 36561 6822
rect 36632 6751 36656 6822
rect 36727 6751 36765 6822
rect 36836 6751 36860 6822
rect 36931 6751 36954 6822
rect 42396 6838 42422 7250
rect 42634 6838 42660 7250
rect 42396 6814 42660 6838
rect 36540 6732 36954 6751
rect 41602 6788 42164 6806
rect 41602 6638 41930 6788
rect 42142 6638 42164 6788
rect 41602 6624 42164 6638
rect 37392 6305 37542 6330
rect 37392 6241 37431 6305
rect 37495 6241 37542 6305
rect 37392 6193 37542 6241
rect 37392 6129 37430 6193
rect 37494 6129 37542 6193
rect 1046 6106 1460 6126
rect 1046 6035 1067 6106
rect 1138 6035 1162 6106
rect 1233 6035 1271 6106
rect 1342 6035 1366 6106
rect 1437 6035 1460 6106
rect 1046 6016 1460 6035
rect 36064 6106 36478 6126
rect 36064 6035 36085 6106
rect 36156 6035 36180 6106
rect 36251 6035 36289 6106
rect 36360 6035 36384 6106
rect 36455 6035 36478 6106
rect 36064 6016 36478 6035
rect 37392 6075 37542 6129
rect 41602 6246 42164 6264
rect 41602 6096 41930 6246
rect 42142 6096 42164 6246
rect 41602 6082 42164 6096
rect 37392 6011 37430 6075
rect 37494 6011 37542 6075
rect 37392 5986 37542 6011
rect 570 5818 984 5838
rect 570 5747 591 5818
rect 662 5747 686 5818
rect 757 5747 795 5818
rect 866 5747 890 5818
rect 961 5747 984 5818
rect 570 5728 984 5747
rect 36540 5818 36954 5838
rect 36540 5747 36561 5818
rect 36632 5747 36656 5818
rect 36727 5747 36765 5818
rect 36836 5747 36860 5818
rect 36931 5747 36954 5818
rect 36540 5728 36954 5747
rect 41602 5690 42164 5708
rect 41602 5540 41930 5690
rect 42142 5540 42164 5690
rect 41602 5526 42164 5540
rect 42396 5492 42660 5518
rect 1046 5102 1460 5122
rect 1046 5031 1067 5102
rect 1138 5031 1162 5102
rect 1233 5031 1271 5102
rect 1342 5031 1366 5102
rect 1437 5031 1460 5102
rect 1046 5012 1460 5031
rect 36064 5102 36478 5122
rect 36064 5031 36085 5102
rect 36156 5031 36180 5102
rect 36251 5031 36289 5102
rect 36360 5031 36384 5102
rect 36455 5031 36478 5102
rect 42396 5080 42422 5492
rect 42634 5080 42660 5492
rect 42396 5056 42660 5080
rect 36064 5012 36478 5031
rect 570 4814 984 4834
rect 570 4743 591 4814
rect 662 4743 686 4814
rect 757 4743 795 4814
rect 866 4743 890 4814
rect 961 4743 984 4814
rect 570 4724 984 4743
rect 36540 4814 36954 4834
rect 36540 4743 36561 4814
rect 36632 4743 36656 4814
rect 36727 4743 36765 4814
rect 36836 4743 36860 4814
rect 36931 4743 36954 4814
rect 36540 4724 36954 4743
rect 41684 4546 42660 4558
rect 41684 4545 42410 4546
rect 41684 4388 41707 4545
rect 41821 4388 42410 4545
rect 41684 4384 42410 4388
rect 42648 4384 42660 4546
rect 41684 4374 42660 4384
rect 1046 4098 1460 4118
rect 1046 4027 1067 4098
rect 1138 4027 1162 4098
rect 1233 4027 1271 4098
rect 1342 4027 1366 4098
rect 1437 4027 1460 4098
rect 1046 4008 1460 4027
rect 36064 4098 36478 4118
rect 36064 4027 36085 4098
rect 36156 4027 36180 4098
rect 36251 4027 36289 4098
rect 36360 4027 36384 4098
rect 36455 4027 36478 4098
rect 36064 4008 36478 4027
rect 570 3810 984 3830
rect 570 3739 591 3810
rect 662 3739 686 3810
rect 757 3739 795 3810
rect 866 3739 890 3810
rect 961 3739 984 3810
rect 570 3720 984 3739
rect 36540 3810 36954 3830
rect 36540 3739 36561 3810
rect 36632 3739 36656 3810
rect 36727 3739 36765 3810
rect 36836 3739 36860 3810
rect 36931 3739 36954 3810
rect 36540 3720 36954 3739
rect 41684 3656 42660 3668
rect 41684 3655 42410 3656
rect 36064 3589 37512 3617
rect 36064 3525 36094 3589
rect 36158 3525 36190 3589
rect 36254 3525 36286 3589
rect 36350 3525 36382 3589
rect 36446 3587 37512 3589
rect 36446 3525 37423 3587
rect 36064 3523 37423 3525
rect 37487 3523 37512 3587
rect 36064 3498 37512 3523
rect 36064 3434 36094 3498
rect 36158 3434 36190 3498
rect 36254 3434 36286 3498
rect 36350 3434 36382 3498
rect 36446 3495 37512 3498
rect 36446 3434 37423 3495
rect 36064 3431 37423 3434
rect 37487 3431 37512 3495
rect 41684 3498 41707 3655
rect 41821 3498 42410 3655
rect 41684 3494 42410 3498
rect 42648 3494 42660 3656
rect 41684 3484 42660 3494
rect 36064 3407 37512 3431
rect 36064 3343 36094 3407
rect 36158 3343 36190 3407
rect 36254 3343 36286 3407
rect 36350 3343 36382 3407
rect 36446 3404 37512 3407
rect 36446 3343 37423 3404
rect 36064 3340 37423 3343
rect 37487 3340 37512 3404
rect 36064 3318 37512 3340
rect 42396 3250 42660 3276
rect 1046 3092 1460 3112
rect 1046 3021 1067 3092
rect 1138 3021 1162 3092
rect 1233 3021 1271 3092
rect 1342 3021 1366 3092
rect 1437 3021 1460 3092
rect 1046 3002 1460 3021
rect 36064 3094 36478 3114
rect 36064 3023 36085 3094
rect 36156 3023 36180 3094
rect 36251 3023 36289 3094
rect 36360 3023 36384 3094
rect 36455 3023 36478 3094
rect 36064 3004 36478 3023
rect 42396 2838 42422 3250
rect 42634 2838 42660 3250
rect 570 2806 984 2826
rect 570 2735 591 2806
rect 662 2735 686 2806
rect 757 2735 795 2806
rect 866 2735 890 2806
rect 961 2735 984 2806
rect 570 2716 984 2735
rect 36540 2806 36954 2826
rect 42396 2814 42660 2838
rect 36540 2735 36561 2806
rect 36632 2735 36656 2806
rect 36727 2735 36765 2806
rect 36836 2735 36860 2806
rect 36931 2735 36954 2806
rect 36540 2716 36954 2735
rect 41602 2788 42164 2806
rect 41602 2638 41930 2788
rect 42142 2638 42164 2788
rect 41602 2624 42164 2638
rect 37392 2311 37542 2336
rect 37392 2247 37431 2311
rect 37495 2247 37542 2311
rect 37392 2199 37542 2247
rect 37392 2135 37430 2199
rect 37494 2135 37542 2199
rect 1046 2089 1460 2109
rect 1046 2018 1067 2089
rect 1138 2018 1162 2089
rect 1233 2018 1271 2089
rect 1342 2018 1366 2089
rect 1437 2018 1460 2089
rect 1046 1999 1460 2018
rect 36064 2090 36478 2110
rect 36064 2019 36085 2090
rect 36156 2019 36180 2090
rect 36251 2019 36289 2090
rect 36360 2019 36384 2090
rect 36455 2019 36478 2090
rect 36064 2000 36478 2019
rect 37392 2081 37542 2135
rect 41602 2246 42164 2264
rect 41602 2096 41930 2246
rect 42142 2096 42164 2246
rect 41602 2082 42164 2096
rect 37392 2017 37430 2081
rect 37494 2017 37542 2081
rect 37392 1992 37542 2017
rect 36540 1802 36954 1822
rect 570 1748 984 1768
rect 570 1677 591 1748
rect 662 1677 686 1748
rect 757 1677 795 1748
rect 866 1677 890 1748
rect 961 1677 984 1748
rect 36540 1731 36561 1802
rect 36632 1731 36656 1802
rect 36727 1731 36765 1802
rect 36836 1731 36860 1802
rect 36931 1731 36954 1802
rect 36540 1712 36954 1731
rect 570 1658 984 1677
rect 41602 1690 42164 1708
rect 41602 1540 41930 1690
rect 42142 1540 42164 1690
rect 41602 1526 42164 1540
rect 42396 1492 42660 1518
rect 1046 1434 1460 1454
rect 1046 1363 1067 1434
rect 1138 1363 1162 1434
rect 1233 1363 1271 1434
rect 1342 1363 1366 1434
rect 1437 1363 1460 1434
rect 1046 1324 1460 1363
rect 1046 1253 1067 1324
rect 1138 1253 1162 1324
rect 1233 1253 1271 1324
rect 1342 1253 1366 1324
rect 1437 1253 1460 1324
rect 1046 1234 1460 1253
rect 1046 1085 1460 1105
rect 1046 1014 1067 1085
rect 1138 1014 1162 1085
rect 1233 1014 1271 1085
rect 1342 1014 1366 1085
rect 1437 1014 1460 1085
rect 1046 995 1460 1014
rect 36064 1086 36478 1106
rect 36064 1015 36085 1086
rect 36156 1015 36180 1086
rect 36251 1015 36289 1086
rect 36360 1015 36384 1086
rect 36455 1015 36478 1086
rect 42396 1080 42422 1492
rect 42634 1080 42660 1492
rect 42396 1056 42660 1080
rect 36064 996 36478 1015
rect 36064 881 37512 909
rect 570 812 984 832
rect 570 741 591 812
rect 662 741 686 812
rect 757 741 795 812
rect 866 741 890 812
rect 961 772 984 812
rect 36064 817 36094 881
rect 36158 817 36190 881
rect 36254 817 36286 881
rect 36350 817 36382 881
rect 36446 879 37512 881
rect 36446 817 37423 879
rect 36064 815 37423 817
rect 37487 815 37512 879
rect 36064 790 37512 815
rect 961 741 983 772
rect 570 722 983 741
rect 36064 726 36094 790
rect 36158 726 36190 790
rect 36254 726 36286 790
rect 36350 726 36382 790
rect 36446 787 37512 790
rect 36446 726 37423 787
rect 36064 723 37423 726
rect 37487 723 37512 787
rect 36064 699 37512 723
rect 36064 635 36094 699
rect 36158 635 36190 699
rect 36254 635 36286 699
rect 36350 635 36382 699
rect 36446 696 37512 699
rect 36446 635 37423 696
rect 36064 632 37423 635
rect 37487 632 37512 696
rect 36064 610 37512 632
rect 41847 557 42660 558
rect 41684 546 42660 557
rect 36540 526 36954 546
rect 36540 455 36561 526
rect 36632 455 36656 526
rect 36727 455 36765 526
rect 36836 455 36860 526
rect 36931 455 36954 526
rect 36540 436 36954 455
rect 41684 544 42410 546
rect 41684 387 41707 544
rect 41821 387 42410 544
rect 41684 384 42410 387
rect 42648 384 42660 546
rect 41684 374 42660 384
rect 41684 373 41847 374
<< via3 >>
rect 41707 23498 41821 23655
rect 42410 23494 42648 23656
rect 42422 22838 42634 23250
rect 41930 22638 42142 22788
rect 41930 22096 42142 22246
rect 41930 21540 42142 21690
rect 42422 21080 42634 21492
rect 41707 20388 41821 20545
rect 42410 20384 42648 20546
rect 587 19634 969 19889
rect 1063 19196 1445 19451
rect 3444 19638 3770 19882
rect 7444 19638 7770 19882
rect 11444 19638 11770 19882
rect 15444 19638 15770 19882
rect 19444 19638 19770 19882
rect 23444 19638 23770 19882
rect 27444 19638 27770 19882
rect 31444 19638 31770 19882
rect 35426 19783 35490 19847
rect 35522 19783 35586 19847
rect 35618 19783 35682 19847
rect 35714 19783 35778 19847
rect 35426 19689 35490 19753
rect 35522 19689 35586 19753
rect 35618 19689 35682 19753
rect 35714 19689 35778 19753
rect 36570 19821 36634 19885
rect 36666 19821 36730 19885
rect 36762 19821 36826 19885
rect 36858 19821 36922 19885
rect 36570 19727 36634 19791
rect 36666 19727 36730 19791
rect 36762 19727 36826 19791
rect 36858 19727 36922 19791
rect 36094 19493 36158 19557
rect 36190 19493 36254 19557
rect 36286 19493 36350 19557
rect 36382 19493 36446 19557
rect 37423 19551 37487 19555
rect 37423 19495 37427 19551
rect 37427 19495 37483 19551
rect 37483 19495 37487 19551
rect 37423 19491 37487 19495
rect 41707 19498 41821 19655
rect 42410 19494 42648 19656
rect 36094 19402 36158 19466
rect 36190 19402 36254 19466
rect 36286 19402 36350 19466
rect 36382 19402 36446 19466
rect 37423 19460 37487 19463
rect 37423 19404 37427 19460
rect 37427 19404 37483 19460
rect 37483 19404 37487 19460
rect 37423 19399 37487 19404
rect 36094 19311 36158 19375
rect 36190 19311 36254 19375
rect 36286 19311 36350 19375
rect 36382 19311 36446 19375
rect 37423 19369 37487 19372
rect 37423 19313 37427 19369
rect 37427 19313 37483 19369
rect 37483 19313 37487 19369
rect 37423 19308 37487 19313
rect 36094 19217 36158 19281
rect 36190 19217 36254 19281
rect 36286 19217 36350 19281
rect 36382 19217 36446 19281
rect 591 18745 662 18816
rect 686 18745 757 18816
rect 795 18745 866 18816
rect 890 18745 961 18816
rect 36561 18799 36632 18870
rect 36656 18799 36727 18870
rect 36765 18799 36836 18870
rect 36860 18799 36931 18870
rect 42422 18838 42634 19250
rect 41930 18638 42142 18788
rect 591 18431 662 18502
rect 686 18431 757 18502
rect 795 18431 866 18502
rect 890 18431 961 18502
rect 1067 18292 1138 18363
rect 1162 18292 1233 18363
rect 1271 18292 1342 18363
rect 1366 18292 1437 18363
rect 37431 18243 37495 18307
rect 1067 18082 1138 18153
rect 1162 18082 1233 18153
rect 1271 18082 1342 18153
rect 1366 18082 1437 18153
rect 36085 18083 36156 18154
rect 36180 18083 36251 18154
rect 36289 18083 36360 18154
rect 36384 18083 36455 18154
rect 37430 18131 37494 18195
rect 41930 18096 42142 18246
rect 37430 18013 37494 18077
rect 591 17795 662 17866
rect 686 17795 757 17866
rect 795 17795 866 17866
rect 890 17795 961 17866
rect 36561 17795 36632 17866
rect 36656 17795 36727 17866
rect 36765 17795 36836 17866
rect 36860 17795 36931 17866
rect 41930 17540 42142 17690
rect 1067 17079 1138 17150
rect 1162 17079 1233 17150
rect 1271 17079 1342 17150
rect 1366 17079 1437 17150
rect 36085 17079 36156 17150
rect 36180 17079 36251 17150
rect 36289 17079 36360 17150
rect 36384 17079 36455 17150
rect 42422 17080 42634 17492
rect 591 16791 662 16862
rect 686 16791 757 16862
rect 795 16791 866 16862
rect 890 16791 961 16862
rect 36561 16791 36632 16862
rect 36656 16791 36727 16862
rect 36765 16791 36836 16862
rect 36860 16791 36931 16862
rect 36094 16588 36158 16652
rect 36190 16588 36254 16652
rect 36286 16588 36350 16652
rect 36382 16588 36446 16652
rect 37423 16646 37487 16650
rect 37423 16590 37427 16646
rect 37427 16590 37483 16646
rect 37483 16590 37487 16646
rect 37423 16586 37487 16590
rect 36094 16497 36158 16561
rect 36190 16497 36254 16561
rect 36286 16497 36350 16561
rect 36382 16497 36446 16561
rect 37423 16555 37487 16558
rect 37423 16499 37427 16555
rect 37427 16499 37483 16555
rect 37483 16499 37487 16555
rect 37423 16494 37487 16499
rect 36094 16406 36158 16470
rect 36190 16406 36254 16470
rect 36286 16406 36350 16470
rect 36382 16406 36446 16470
rect 37423 16464 37487 16467
rect 37423 16408 37427 16464
rect 37427 16408 37483 16464
rect 37483 16408 37487 16464
rect 37423 16403 37487 16408
rect 41707 16388 41821 16545
rect 42410 16384 42648 16546
rect 1067 16074 1138 16145
rect 1162 16074 1233 16145
rect 1271 16074 1342 16145
rect 1366 16074 1437 16145
rect 36085 16075 36156 16146
rect 36180 16075 36251 16146
rect 36289 16075 36360 16146
rect 36384 16075 36455 16146
rect 591 15787 662 15858
rect 686 15787 757 15858
rect 795 15787 866 15858
rect 890 15787 961 15858
rect 36561 15787 36632 15858
rect 36656 15787 36727 15858
rect 36765 15787 36836 15858
rect 36860 15787 36931 15858
rect 41707 15498 41821 15655
rect 42410 15494 42648 15656
rect 1067 15071 1138 15142
rect 1162 15071 1233 15142
rect 1271 15071 1342 15142
rect 1366 15071 1437 15142
rect 36085 15071 36156 15142
rect 36180 15071 36251 15142
rect 36289 15071 36360 15142
rect 36384 15071 36455 15142
rect 591 14783 662 14854
rect 686 14783 757 14854
rect 795 14783 866 14854
rect 890 14783 961 14854
rect 36561 14783 36632 14854
rect 36656 14783 36727 14854
rect 36765 14783 36836 14854
rect 36860 14783 36931 14854
rect 42422 14838 42634 15250
rect 41930 14638 42142 14788
rect 37431 14243 37495 14307
rect 1067 14067 1138 14138
rect 1162 14067 1233 14138
rect 1271 14067 1342 14138
rect 1366 14067 1437 14138
rect 36085 14067 36156 14138
rect 36180 14067 36251 14138
rect 36289 14067 36360 14138
rect 36384 14067 36455 14138
rect 37430 14131 37494 14195
rect 41930 14096 42142 14246
rect 37430 14013 37494 14077
rect 591 13779 662 13850
rect 686 13779 757 13850
rect 795 13779 866 13850
rect 890 13779 961 13850
rect 36561 13779 36632 13850
rect 36656 13779 36727 13850
rect 36765 13779 36836 13850
rect 36860 13779 36931 13850
rect 41930 13540 42142 13690
rect 1067 13063 1138 13134
rect 1162 13063 1233 13134
rect 1271 13063 1342 13134
rect 1366 13063 1437 13134
rect 36085 13063 36156 13134
rect 36180 13063 36251 13134
rect 36289 13063 36360 13134
rect 36384 13063 36455 13134
rect 42422 13080 42634 13492
rect 591 12775 662 12846
rect 686 12775 757 12846
rect 795 12775 866 12846
rect 890 12775 961 12846
rect 36561 12775 36632 12846
rect 36656 12775 36727 12846
rect 36765 12775 36836 12846
rect 36860 12775 36931 12846
rect 36094 12530 36158 12594
rect 36190 12530 36254 12594
rect 36286 12530 36350 12594
rect 36382 12530 36446 12594
rect 37423 12588 37487 12592
rect 37423 12532 37427 12588
rect 37427 12532 37483 12588
rect 37483 12532 37487 12588
rect 37423 12528 37487 12532
rect 36094 12439 36158 12503
rect 36190 12439 36254 12503
rect 36286 12439 36350 12503
rect 36382 12439 36446 12503
rect 37423 12497 37487 12500
rect 37423 12441 37427 12497
rect 37427 12441 37483 12497
rect 37483 12441 37487 12497
rect 37423 12436 37487 12441
rect 36094 12348 36158 12412
rect 36190 12348 36254 12412
rect 36286 12348 36350 12412
rect 36382 12348 36446 12412
rect 37423 12406 37487 12409
rect 37423 12350 37427 12406
rect 37427 12350 37483 12406
rect 37483 12350 37487 12406
rect 37423 12345 37487 12350
rect 41707 12388 41821 12545
rect 42410 12384 42648 12546
rect 1067 12059 1138 12130
rect 1162 12059 1233 12130
rect 1271 12059 1342 12130
rect 1366 12059 1437 12130
rect 36085 12059 36156 12130
rect 36180 12059 36251 12130
rect 36289 12059 36360 12130
rect 36384 12059 36455 12130
rect 591 11771 662 11842
rect 686 11771 757 11842
rect 795 11771 866 11842
rect 890 11771 961 11842
rect 36561 11771 36632 11842
rect 36656 11771 36727 11842
rect 36765 11771 36836 11842
rect 36860 11771 36931 11842
rect 41707 11498 41821 11655
rect 42410 11494 42648 11656
rect 1067 11055 1138 11126
rect 1162 11055 1233 11126
rect 1271 11055 1342 11126
rect 1366 11055 1437 11126
rect 36085 11055 36156 11126
rect 36180 11055 36251 11126
rect 36289 11055 36360 11126
rect 36384 11055 36455 11126
rect 591 10767 662 10838
rect 686 10767 757 10838
rect 795 10767 866 10838
rect 890 10767 961 10838
rect 36561 10767 36632 10838
rect 36656 10767 36727 10838
rect 36765 10767 36836 10838
rect 36860 10767 36931 10838
rect 42422 10838 42634 11250
rect 41930 10638 42142 10788
rect 37431 10243 37495 10307
rect 1067 10051 1138 10122
rect 1162 10051 1233 10122
rect 1271 10051 1342 10122
rect 1366 10051 1437 10122
rect 36085 10051 36156 10122
rect 36180 10051 36251 10122
rect 36289 10051 36360 10122
rect 36384 10051 36455 10122
rect 37430 10131 37494 10195
rect 41930 10096 42142 10246
rect 37430 10013 37494 10077
rect 591 9763 662 9834
rect 686 9763 757 9834
rect 795 9763 866 9834
rect 890 9763 961 9834
rect 36561 9763 36632 9834
rect 36656 9763 36727 9834
rect 36765 9763 36836 9834
rect 36860 9763 36931 9834
rect 41930 9540 42142 9690
rect 1067 9047 1138 9118
rect 1162 9047 1233 9118
rect 1271 9047 1342 9118
rect 1366 9047 1437 9118
rect 36085 9047 36156 9118
rect 36180 9047 36251 9118
rect 36289 9047 36360 9118
rect 36384 9047 36455 9118
rect 42422 9080 42634 9492
rect 591 8759 662 8830
rect 686 8759 757 8830
rect 795 8759 866 8830
rect 890 8759 961 8830
rect 36561 8759 36632 8830
rect 36656 8759 36727 8830
rect 36765 8759 36836 8830
rect 36860 8759 36931 8830
rect 36094 8437 36158 8501
rect 36190 8437 36254 8501
rect 36286 8437 36350 8501
rect 36382 8437 36446 8501
rect 37423 8495 37487 8499
rect 37423 8439 37427 8495
rect 37427 8439 37483 8495
rect 37483 8439 37487 8495
rect 37423 8435 37487 8439
rect 36094 8346 36158 8410
rect 36190 8346 36254 8410
rect 36286 8346 36350 8410
rect 36382 8346 36446 8410
rect 37423 8404 37487 8407
rect 37423 8348 37427 8404
rect 37427 8348 37483 8404
rect 37483 8348 37487 8404
rect 37423 8343 37487 8348
rect 41707 8388 41821 8545
rect 42410 8384 42648 8546
rect 36094 8255 36158 8319
rect 36190 8255 36254 8319
rect 36286 8255 36350 8319
rect 36382 8255 36446 8319
rect 37423 8313 37487 8316
rect 37423 8257 37427 8313
rect 37427 8257 37483 8313
rect 37483 8257 37487 8313
rect 37423 8252 37487 8257
rect 1067 8043 1138 8114
rect 1162 8043 1233 8114
rect 1271 8043 1342 8114
rect 1366 8043 1437 8114
rect 36085 8043 36156 8114
rect 36180 8043 36251 8114
rect 36289 8043 36360 8114
rect 36384 8043 36455 8114
rect 591 7755 662 7826
rect 686 7755 757 7826
rect 795 7755 866 7826
rect 890 7755 961 7826
rect 36561 7755 36632 7826
rect 36656 7755 36727 7826
rect 36765 7755 36836 7826
rect 36860 7755 36931 7826
rect 41707 7498 41821 7655
rect 42410 7494 42648 7656
rect 1067 7039 1138 7110
rect 1162 7039 1233 7110
rect 1271 7039 1342 7110
rect 1366 7039 1437 7110
rect 36085 7039 36156 7110
rect 36180 7039 36251 7110
rect 36289 7039 36360 7110
rect 36384 7039 36455 7110
rect 591 6751 662 6822
rect 686 6751 757 6822
rect 795 6751 866 6822
rect 890 6751 961 6822
rect 36561 6751 36632 6822
rect 36656 6751 36727 6822
rect 36765 6751 36836 6822
rect 36860 6751 36931 6822
rect 42422 6838 42634 7250
rect 41930 6638 42142 6788
rect 37431 6241 37495 6305
rect 37430 6129 37494 6193
rect 1067 6035 1138 6106
rect 1162 6035 1233 6106
rect 1271 6035 1342 6106
rect 1366 6035 1437 6106
rect 36085 6035 36156 6106
rect 36180 6035 36251 6106
rect 36289 6035 36360 6106
rect 36384 6035 36455 6106
rect 41930 6096 42142 6246
rect 37430 6011 37494 6075
rect 591 5747 662 5818
rect 686 5747 757 5818
rect 795 5747 866 5818
rect 890 5747 961 5818
rect 36561 5747 36632 5818
rect 36656 5747 36727 5818
rect 36765 5747 36836 5818
rect 36860 5747 36931 5818
rect 41930 5540 42142 5690
rect 1067 5031 1138 5102
rect 1162 5031 1233 5102
rect 1271 5031 1342 5102
rect 1366 5031 1437 5102
rect 36085 5031 36156 5102
rect 36180 5031 36251 5102
rect 36289 5031 36360 5102
rect 36384 5031 36455 5102
rect 42422 5080 42634 5492
rect 591 4743 662 4814
rect 686 4743 757 4814
rect 795 4743 866 4814
rect 890 4743 961 4814
rect 36561 4743 36632 4814
rect 36656 4743 36727 4814
rect 36765 4743 36836 4814
rect 36860 4743 36931 4814
rect 41707 4388 41821 4545
rect 42410 4384 42648 4546
rect 1067 4027 1138 4098
rect 1162 4027 1233 4098
rect 1271 4027 1342 4098
rect 1366 4027 1437 4098
rect 36085 4027 36156 4098
rect 36180 4027 36251 4098
rect 36289 4027 36360 4098
rect 36384 4027 36455 4098
rect 591 3739 662 3810
rect 686 3739 757 3810
rect 795 3739 866 3810
rect 890 3739 961 3810
rect 36561 3739 36632 3810
rect 36656 3739 36727 3810
rect 36765 3739 36836 3810
rect 36860 3739 36931 3810
rect 36094 3525 36158 3589
rect 36190 3525 36254 3589
rect 36286 3525 36350 3589
rect 36382 3525 36446 3589
rect 37423 3583 37487 3587
rect 37423 3527 37427 3583
rect 37427 3527 37483 3583
rect 37483 3527 37487 3583
rect 37423 3523 37487 3527
rect 36094 3434 36158 3498
rect 36190 3434 36254 3498
rect 36286 3434 36350 3498
rect 36382 3434 36446 3498
rect 37423 3492 37487 3495
rect 37423 3436 37427 3492
rect 37427 3436 37483 3492
rect 37483 3436 37487 3492
rect 37423 3431 37487 3436
rect 41707 3498 41821 3655
rect 42410 3494 42648 3656
rect 36094 3343 36158 3407
rect 36190 3343 36254 3407
rect 36286 3343 36350 3407
rect 36382 3343 36446 3407
rect 37423 3401 37487 3404
rect 37423 3345 37427 3401
rect 37427 3345 37483 3401
rect 37483 3345 37487 3401
rect 37423 3340 37487 3345
rect 1067 3021 1138 3092
rect 1162 3021 1233 3092
rect 1271 3021 1342 3092
rect 1366 3021 1437 3092
rect 36085 3023 36156 3094
rect 36180 3023 36251 3094
rect 36289 3023 36360 3094
rect 36384 3023 36455 3094
rect 42422 2838 42634 3250
rect 591 2735 662 2806
rect 686 2735 757 2806
rect 795 2735 866 2806
rect 890 2735 961 2806
rect 36561 2735 36632 2806
rect 36656 2735 36727 2806
rect 36765 2735 36836 2806
rect 36860 2735 36931 2806
rect 41930 2638 42142 2788
rect 37431 2247 37495 2311
rect 37430 2135 37494 2199
rect 1067 2018 1138 2089
rect 1162 2018 1233 2089
rect 1271 2018 1342 2089
rect 1366 2018 1437 2089
rect 36085 2019 36156 2090
rect 36180 2019 36251 2090
rect 36289 2019 36360 2090
rect 36384 2019 36455 2090
rect 41930 2096 42142 2246
rect 37430 2017 37494 2081
rect 591 1677 662 1748
rect 686 1677 757 1748
rect 795 1677 866 1748
rect 890 1677 961 1748
rect 36561 1731 36632 1802
rect 36656 1731 36727 1802
rect 36765 1731 36836 1802
rect 36860 1731 36931 1802
rect 41930 1540 42142 1690
rect 1067 1363 1138 1434
rect 1162 1363 1233 1434
rect 1271 1363 1342 1434
rect 1366 1363 1437 1434
rect 1067 1253 1138 1324
rect 1162 1253 1233 1324
rect 1271 1253 1342 1324
rect 1366 1253 1437 1324
rect 1067 1014 1138 1085
rect 1162 1014 1233 1085
rect 1271 1014 1342 1085
rect 1366 1014 1437 1085
rect 36085 1015 36156 1086
rect 36180 1015 36251 1086
rect 36289 1015 36360 1086
rect 36384 1015 36455 1086
rect 42422 1080 42634 1492
rect 591 741 662 812
rect 686 741 757 812
rect 795 741 866 812
rect 890 741 961 812
rect 36094 817 36158 881
rect 36190 817 36254 881
rect 36286 817 36350 881
rect 36382 817 36446 881
rect 37423 875 37487 879
rect 37423 819 37427 875
rect 37427 819 37483 875
rect 37483 819 37487 875
rect 37423 815 37487 819
rect 36094 726 36158 790
rect 36190 726 36254 790
rect 36286 726 36350 790
rect 36382 726 36446 790
rect 37423 784 37487 787
rect 37423 728 37427 784
rect 37427 728 37483 784
rect 37483 728 37487 784
rect 37423 723 37487 728
rect 36094 635 36158 699
rect 36190 635 36254 699
rect 36286 635 36350 699
rect 36382 635 36446 699
rect 37423 693 37487 696
rect 37423 637 37427 693
rect 37427 637 37483 693
rect 37483 637 37487 693
rect 37423 632 37487 637
rect 36561 455 36632 526
rect 36656 455 36727 526
rect 36765 455 36836 526
rect 36860 455 36931 526
rect 41707 387 41821 544
rect 42410 384 42648 546
<< metal4 >>
rect 570 19889 984 24166
rect 570 19634 587 19889
rect 969 19634 984 19889
rect 570 18816 984 19634
rect 570 18745 591 18816
rect 662 18745 686 18816
rect 757 18745 795 18816
rect 866 18745 890 18816
rect 961 18745 984 18816
rect 570 18502 984 18745
rect 570 18431 591 18502
rect 662 18431 686 18502
rect 757 18431 795 18502
rect 866 18431 890 18502
rect 961 18431 984 18502
rect 570 17866 984 18431
rect 570 17795 591 17866
rect 662 17795 686 17866
rect 757 17795 795 17866
rect 866 17795 890 17866
rect 961 17795 984 17866
rect 570 16862 984 17795
rect 570 16791 591 16862
rect 662 16791 686 16862
rect 757 16791 795 16862
rect 866 16791 890 16862
rect 961 16791 984 16862
rect 570 15858 984 16791
rect 570 15787 591 15858
rect 662 15787 686 15858
rect 757 15787 795 15858
rect 866 15787 890 15858
rect 961 15787 984 15858
rect 570 14854 984 15787
rect 570 14783 591 14854
rect 662 14783 686 14854
rect 757 14783 795 14854
rect 866 14783 890 14854
rect 961 14783 984 14854
rect 570 13850 984 14783
rect 570 13779 591 13850
rect 662 13779 686 13850
rect 757 13779 795 13850
rect 866 13779 890 13850
rect 961 13779 984 13850
rect 570 12846 984 13779
rect 570 12775 591 12846
rect 662 12775 686 12846
rect 757 12775 795 12846
rect 866 12775 890 12846
rect 961 12775 984 12846
rect 570 11842 984 12775
rect 570 11771 591 11842
rect 662 11771 686 11842
rect 757 11771 795 11842
rect 866 11771 890 11842
rect 961 11771 984 11842
rect 570 10838 984 11771
rect 570 10767 591 10838
rect 662 10767 686 10838
rect 757 10767 795 10838
rect 866 10767 890 10838
rect 961 10767 984 10838
rect 570 9834 984 10767
rect 570 9763 591 9834
rect 662 9763 686 9834
rect 757 9763 795 9834
rect 866 9763 890 9834
rect 961 9763 984 9834
rect 570 8830 984 9763
rect 570 8759 591 8830
rect 662 8759 686 8830
rect 757 8759 795 8830
rect 866 8759 890 8830
rect 961 8759 984 8830
rect 570 7826 984 8759
rect 570 7755 591 7826
rect 662 7755 686 7826
rect 757 7755 795 7826
rect 866 7755 890 7826
rect 961 7755 984 7826
rect 570 6822 984 7755
rect 570 6751 591 6822
rect 662 6751 686 6822
rect 757 6751 795 6822
rect 866 6751 890 6822
rect 961 6751 984 6822
rect 570 5818 984 6751
rect 570 5747 591 5818
rect 662 5747 686 5818
rect 757 5747 795 5818
rect 866 5747 890 5818
rect 961 5747 984 5818
rect 570 4814 984 5747
rect 570 4743 591 4814
rect 662 4743 686 4814
rect 757 4743 795 4814
rect 866 4743 890 4814
rect 961 4743 984 4814
rect 570 3810 984 4743
rect 570 3739 591 3810
rect 662 3739 686 3810
rect 757 3739 795 3810
rect 866 3739 890 3810
rect 961 3739 984 3810
rect 570 2806 984 3739
rect 570 2735 591 2806
rect 662 2735 686 2806
rect 757 2735 795 2806
rect 866 2735 890 2806
rect 961 2735 984 2806
rect 570 1748 984 2735
rect 570 1677 591 1748
rect 662 1677 686 1748
rect 757 1677 795 1748
rect 866 1677 890 1748
rect 961 1677 984 1748
rect 570 812 984 1677
rect 570 741 591 812
rect 662 741 686 812
rect 757 741 795 812
rect 866 741 890 812
rect 961 741 984 812
rect 570 42 984 741
rect 1046 19451 1460 24166
rect 41602 23655 41847 23668
rect 41602 23498 41707 23655
rect 41821 23498 41847 23655
rect 41602 23484 41847 23498
rect 41908 22806 42322 24166
rect 41602 22788 42322 22806
rect 41602 22638 41930 22788
rect 42142 22638 42322 22788
rect 41602 22624 42322 22638
rect 41908 22264 42322 22624
rect 41602 22246 42322 22264
rect 41602 22096 41930 22246
rect 42142 22096 42322 22246
rect 41602 22082 42322 22096
rect 41908 21708 42322 22082
rect 41602 21690 42322 21708
rect 41602 21540 41930 21690
rect 42142 21540 42322 21690
rect 41602 21526 42322 21540
rect 41602 20545 41847 20558
rect 41602 20388 41707 20545
rect 41821 20388 41847 20545
rect 41602 20374 41847 20388
rect 3420 19882 3790 20166
rect 3420 19638 3444 19882
rect 3770 19638 3790 19882
rect 3420 19620 3790 19638
rect 7420 19882 7790 20166
rect 7420 19638 7444 19882
rect 7770 19638 7790 19882
rect 7420 19620 7790 19638
rect 11420 19882 11790 20166
rect 11420 19638 11444 19882
rect 11770 19638 11790 19882
rect 11420 19620 11790 19638
rect 15420 19882 15790 20166
rect 15420 19638 15444 19882
rect 15770 19638 15790 19882
rect 15420 19620 15790 19638
rect 19420 19882 19790 20166
rect 19420 19638 19444 19882
rect 19770 19638 19790 19882
rect 19420 19620 19790 19638
rect 23420 19882 23790 20166
rect 23420 19638 23444 19882
rect 23770 19638 23790 19882
rect 23420 19620 23790 19638
rect 27420 19882 27790 20166
rect 27420 19638 27444 19882
rect 27770 19638 27790 19882
rect 27420 19620 27790 19638
rect 31420 19882 31790 20166
rect 35412 19900 35782 20166
rect 31420 19638 31444 19882
rect 31770 19638 31790 19882
rect 31420 19620 31790 19638
rect 35396 19847 35810 19900
rect 35396 19783 35426 19847
rect 35490 19783 35522 19847
rect 35586 19783 35618 19847
rect 35682 19783 35714 19847
rect 35778 19783 35810 19847
rect 35396 19753 35810 19783
rect 35396 19689 35426 19753
rect 35490 19689 35522 19753
rect 35586 19689 35618 19753
rect 35682 19689 35714 19753
rect 35778 19689 35810 19753
rect 35396 19620 35810 19689
rect 1046 19196 1063 19451
rect 1445 19196 1460 19451
rect 1046 18363 1460 19196
rect 1046 18292 1067 18363
rect 1138 18292 1162 18363
rect 1233 18292 1271 18363
rect 1342 18292 1366 18363
rect 1437 18292 1460 18363
rect 1046 18153 1460 18292
rect 1046 18082 1067 18153
rect 1138 18082 1162 18153
rect 1233 18082 1271 18153
rect 1342 18082 1366 18153
rect 1437 18082 1460 18153
rect 1046 17150 1460 18082
rect 36064 19557 36478 19902
rect 36064 19493 36094 19557
rect 36158 19493 36190 19557
rect 36254 19493 36286 19557
rect 36350 19493 36382 19557
rect 36446 19493 36478 19557
rect 36064 19466 36478 19493
rect 36064 19402 36094 19466
rect 36158 19402 36190 19466
rect 36254 19402 36286 19466
rect 36350 19402 36382 19466
rect 36446 19402 36478 19466
rect 36064 19375 36478 19402
rect 36064 19311 36094 19375
rect 36158 19311 36190 19375
rect 36254 19311 36286 19375
rect 36350 19311 36382 19375
rect 36446 19311 36478 19375
rect 36064 19281 36478 19311
rect 36064 19217 36094 19281
rect 36158 19217 36190 19281
rect 36254 19217 36286 19281
rect 36350 19217 36382 19281
rect 36446 19217 36478 19281
rect 36064 18662 36478 19217
rect 36540 19885 36954 19902
rect 36540 19821 36570 19885
rect 36634 19821 36666 19885
rect 36730 19821 36762 19885
rect 36826 19821 36858 19885
rect 36922 19821 36954 19885
rect 36540 19791 36954 19821
rect 36540 19727 36570 19791
rect 36634 19727 36666 19791
rect 36730 19727 36762 19791
rect 36826 19727 36858 19791
rect 36922 19727 36954 19791
rect 36540 18870 36954 19727
rect 41602 19655 41847 19668
rect 37394 19555 37602 19585
rect 37394 19491 37423 19555
rect 37487 19491 37602 19555
rect 37394 19463 37602 19491
rect 41602 19498 41707 19655
rect 41821 19498 41847 19655
rect 41602 19484 41847 19498
rect 37394 19399 37423 19463
rect 37487 19399 37602 19463
rect 37394 19372 37602 19399
rect 37394 19308 37423 19372
rect 37487 19308 37602 19372
rect 37394 19286 37602 19308
rect 36540 18799 36561 18870
rect 36632 18799 36656 18870
rect 36727 18799 36765 18870
rect 36836 18799 36860 18870
rect 36931 18799 36954 18870
rect 41908 18806 42322 21526
rect 36064 18380 36480 18662
rect 36064 18154 36478 18380
rect 36064 18083 36085 18154
rect 36156 18083 36180 18154
rect 36251 18083 36289 18154
rect 36360 18083 36384 18154
rect 36455 18083 36478 18154
rect 2888 17912 2948 17946
rect 3464 17912 3524 17946
rect 3892 17912 3952 17946
rect 4468 17912 4528 17946
rect 4896 17912 4956 17946
rect 5472 17912 5532 17946
rect 5900 17912 5960 17946
rect 6476 17912 6536 17946
rect 6904 17912 6964 17946
rect 7480 17912 7540 17946
rect 7908 17912 7968 17946
rect 8484 17912 8544 17946
rect 8912 17912 8972 17946
rect 9488 17912 9548 17946
rect 9916 17912 9976 17946
rect 10492 17912 10552 17946
rect 10920 17912 10980 17946
rect 11496 17912 11556 17946
rect 11924 17912 11984 17946
rect 12500 17912 12560 17946
rect 12928 17912 12988 17946
rect 13504 17912 13564 17946
rect 13932 17912 13992 17946
rect 14508 17912 14568 17946
rect 14936 17912 14996 17946
rect 15512 17912 15572 17946
rect 15940 17912 16000 17946
rect 16516 17912 16576 17946
rect 16944 17912 17004 17946
rect 17520 17912 17580 17946
rect 17948 17912 18008 17946
rect 18524 17912 18584 17946
rect 18952 17912 19012 17946
rect 19528 17912 19588 17946
rect 19956 17912 20016 17946
rect 20532 17912 20592 17946
rect 20960 17912 21020 17946
rect 21536 17912 21596 17946
rect 21964 17912 22024 17946
rect 22540 17912 22600 17946
rect 22968 17912 23028 17946
rect 23544 17912 23604 17946
rect 23972 17912 24032 17946
rect 24548 17912 24608 17946
rect 24976 17912 25036 17946
rect 25552 17912 25612 17946
rect 25980 17912 26040 17946
rect 26556 17912 26616 17946
rect 26984 17912 27044 17946
rect 27560 17912 27620 17946
rect 27988 17912 28048 17946
rect 28564 17912 28624 17946
rect 28992 17912 29052 17946
rect 29568 17912 29628 17946
rect 29996 17912 30056 17946
rect 30572 17912 30632 17946
rect 31000 17912 31060 17946
rect 31576 17912 31636 17946
rect 32004 17912 32064 17946
rect 32580 17912 32640 17946
rect 33008 17912 33068 17946
rect 33584 17912 33644 17946
rect 34012 17912 34072 17946
rect 34588 17912 34648 17946
rect 2736 17738 2774 17798
rect 3638 17738 3778 17798
rect 4642 17738 4782 17798
rect 5646 17738 5786 17798
rect 6650 17738 6790 17798
rect 7654 17738 7794 17798
rect 8658 17738 8798 17798
rect 9662 17738 9802 17798
rect 10666 17738 10806 17798
rect 11670 17738 11810 17798
rect 12674 17738 12814 17798
rect 13678 17738 13818 17798
rect 14682 17738 14822 17798
rect 15686 17738 15826 17798
rect 16690 17738 16830 17798
rect 17694 17738 17834 17798
rect 18698 17738 18838 17798
rect 19702 17738 19842 17798
rect 20706 17738 20846 17798
rect 21710 17738 21850 17798
rect 22714 17738 22854 17798
rect 23718 17738 23858 17798
rect 24722 17738 24862 17798
rect 25726 17738 25866 17798
rect 26730 17738 26870 17798
rect 27734 17738 27874 17798
rect 28738 17738 28878 17798
rect 29742 17738 29882 17798
rect 30746 17738 30886 17798
rect 31750 17738 31890 17798
rect 32754 17738 32894 17798
rect 33758 17738 33898 17798
rect 34762 17738 34796 17798
rect 2736 17162 2774 17222
rect 3638 17162 3778 17222
rect 4642 17162 4782 17222
rect 5646 17162 5786 17222
rect 6650 17162 6790 17222
rect 7654 17162 7794 17222
rect 8658 17162 8798 17222
rect 9662 17162 9802 17222
rect 10666 17162 10806 17222
rect 11670 17162 11810 17222
rect 12674 17162 12814 17222
rect 13678 17162 13818 17222
rect 14682 17162 14822 17222
rect 15686 17162 15826 17222
rect 16690 17162 16830 17222
rect 17694 17162 17834 17222
rect 18698 17162 18838 17222
rect 19702 17162 19842 17222
rect 20706 17162 20846 17222
rect 21710 17162 21850 17222
rect 22714 17162 22854 17222
rect 23718 17162 23858 17222
rect 24722 17162 24862 17222
rect 25726 17162 25866 17222
rect 26730 17162 26870 17222
rect 27734 17162 27874 17222
rect 28738 17162 28878 17222
rect 29742 17162 29882 17222
rect 30746 17162 30886 17222
rect 31750 17162 31890 17222
rect 32754 17162 32894 17222
rect 33758 17162 33898 17222
rect 34762 17162 34796 17222
rect 1046 17079 1067 17150
rect 1138 17079 1162 17150
rect 1233 17079 1271 17150
rect 1342 17079 1366 17150
rect 1437 17079 1460 17150
rect 1046 16145 1460 17079
rect 36064 17150 36478 18083
rect 36064 17079 36085 17150
rect 36156 17079 36180 17150
rect 36251 17079 36289 17150
rect 36360 17079 36384 17150
rect 36455 17079 36478 17150
rect 2888 16908 2948 17048
rect 3464 16908 3524 17048
rect 3892 16908 3952 17048
rect 4468 16908 4528 17048
rect 4896 16908 4956 17048
rect 5472 16908 5532 17048
rect 5900 16908 5960 17048
rect 6476 16908 6536 17048
rect 6904 16908 6964 17048
rect 7480 16908 7540 17048
rect 7908 16908 7968 17048
rect 8484 16908 8544 17048
rect 8912 16908 8972 17048
rect 9488 16908 9548 17048
rect 9916 16908 9976 17048
rect 10492 16908 10552 17048
rect 10920 16908 10980 17048
rect 11496 16908 11556 17048
rect 11924 16908 11984 17048
rect 12500 16908 12560 17048
rect 12928 16908 12988 17048
rect 13504 16908 13564 17048
rect 13932 16908 13992 17048
rect 14508 16908 14568 17048
rect 14936 16908 14996 17048
rect 15512 16908 15572 17048
rect 15940 16908 16000 17048
rect 16516 16908 16576 17048
rect 16944 16908 17004 17048
rect 17520 16908 17580 17048
rect 17948 16908 18008 17048
rect 18524 16908 18584 17048
rect 18952 16908 19012 17048
rect 19528 16908 19588 17048
rect 19956 16908 20016 17048
rect 20532 16908 20592 17048
rect 20960 16908 21020 17048
rect 21536 16908 21596 17048
rect 21964 16908 22024 17048
rect 22540 16908 22600 17048
rect 22968 16908 23028 17048
rect 23544 16908 23604 17048
rect 23972 16908 24032 17048
rect 24548 16908 24608 17048
rect 24976 16908 25036 17048
rect 25552 16908 25612 17048
rect 25980 16908 26040 17048
rect 26556 16908 26616 17048
rect 26984 16908 27044 17048
rect 27560 16908 27620 17048
rect 27988 16908 28048 17048
rect 28564 16908 28624 17048
rect 28992 16908 29052 17048
rect 29568 16908 29628 17048
rect 29996 16908 30056 17048
rect 30572 16908 30632 17048
rect 31000 16908 31060 17048
rect 31576 16908 31636 17048
rect 32004 16908 32064 17048
rect 32580 16908 32640 17048
rect 33008 16908 33068 17048
rect 33584 16908 33644 17048
rect 34012 16908 34072 17048
rect 34588 16908 34648 17048
rect 2736 16734 2774 16794
rect 3638 16734 3778 16794
rect 4642 16734 4782 16794
rect 5646 16734 5786 16794
rect 6650 16734 6790 16794
rect 7654 16734 7794 16794
rect 8658 16734 8798 16794
rect 9662 16734 9802 16794
rect 10666 16734 10806 16794
rect 11670 16734 11810 16794
rect 12674 16734 12814 16794
rect 13678 16734 13818 16794
rect 14682 16734 14822 16794
rect 15686 16734 15826 16794
rect 16690 16734 16830 16794
rect 17694 16734 17834 16794
rect 18698 16734 18838 16794
rect 19702 16734 19842 16794
rect 20706 16734 20846 16794
rect 21710 16734 21850 16794
rect 22714 16734 22854 16794
rect 23718 16734 23858 16794
rect 24722 16734 24862 16794
rect 25726 16734 25866 16794
rect 26730 16734 26870 16794
rect 27734 16734 27874 16794
rect 28738 16734 28878 16794
rect 29742 16734 29882 16794
rect 30746 16734 30886 16794
rect 31750 16734 31890 16794
rect 32754 16734 32894 16794
rect 33758 16734 33898 16794
rect 34762 16734 34796 16794
rect 36064 16652 36478 17079
rect 36064 16588 36094 16652
rect 36158 16588 36190 16652
rect 36254 16588 36286 16652
rect 36350 16588 36382 16652
rect 36446 16588 36478 16652
rect 36064 16561 36478 16588
rect 36064 16497 36094 16561
rect 36158 16497 36190 16561
rect 36254 16497 36286 16561
rect 36350 16497 36382 16561
rect 36446 16497 36478 16561
rect 36064 16470 36478 16497
rect 36064 16406 36094 16470
rect 36158 16406 36190 16470
rect 36254 16406 36286 16470
rect 36350 16406 36382 16470
rect 36446 16406 36478 16470
rect 2736 16158 2774 16218
rect 3638 16158 3778 16218
rect 4642 16158 4782 16218
rect 5646 16158 5786 16218
rect 6650 16158 6790 16218
rect 7654 16158 7794 16218
rect 8658 16158 8798 16218
rect 9662 16158 9802 16218
rect 10666 16158 10806 16218
rect 11670 16158 11810 16218
rect 12674 16158 12814 16218
rect 13678 16158 13818 16218
rect 14682 16158 14822 16218
rect 15686 16158 15826 16218
rect 16690 16158 16830 16218
rect 17694 16158 17834 16218
rect 18698 16158 18838 16218
rect 19702 16158 19842 16218
rect 20706 16158 20846 16218
rect 21710 16158 21850 16218
rect 22714 16158 22854 16218
rect 23718 16158 23858 16218
rect 24722 16158 24862 16218
rect 25726 16158 25866 16218
rect 26730 16158 26870 16218
rect 27734 16158 27874 16218
rect 28738 16158 28878 16218
rect 29742 16158 29882 16218
rect 30746 16158 30886 16218
rect 31750 16158 31890 16218
rect 32754 16158 32894 16218
rect 33758 16158 33898 16218
rect 34762 16158 34796 16218
rect 1046 16074 1067 16145
rect 1138 16074 1162 16145
rect 1233 16074 1271 16145
rect 1342 16074 1366 16145
rect 1437 16074 1460 16145
rect 1046 15142 1460 16074
rect 36064 16146 36478 16406
rect 36064 16075 36085 16146
rect 36156 16075 36180 16146
rect 36251 16075 36289 16146
rect 36360 16075 36384 16146
rect 36455 16075 36478 16146
rect 2888 15904 2948 16044
rect 3464 15904 3524 16044
rect 3892 15904 3952 16044
rect 4468 15904 4528 16044
rect 4896 15904 4956 16044
rect 5472 15904 5532 16044
rect 5900 15904 5960 16044
rect 6476 15904 6536 16044
rect 6904 15904 6964 16044
rect 7480 15904 7540 16044
rect 7908 15904 7968 16044
rect 8484 15904 8544 16044
rect 8912 15904 8972 16044
rect 9488 15904 9548 16044
rect 9916 15904 9976 16044
rect 10492 15904 10552 16044
rect 10920 15904 10980 16044
rect 11496 15904 11556 16044
rect 11924 15904 11984 16044
rect 12500 15904 12560 16044
rect 12928 15904 12988 16044
rect 13504 15904 13564 16044
rect 13932 15904 13992 16044
rect 14508 15904 14568 16044
rect 14936 15904 14996 16044
rect 15512 15904 15572 16044
rect 15940 15904 16000 16044
rect 16516 15904 16576 16044
rect 16944 15904 17004 16044
rect 17520 15904 17580 16044
rect 17948 15904 18008 16044
rect 18524 15904 18584 16044
rect 18952 15904 19012 16044
rect 19528 15904 19588 16044
rect 19956 15904 20016 16044
rect 20532 15904 20592 16044
rect 20960 15904 21020 16044
rect 21536 15904 21596 16044
rect 21964 15904 22024 16044
rect 22540 15904 22600 16044
rect 22968 15904 23028 16044
rect 23544 15904 23604 16044
rect 23972 15904 24032 16044
rect 24548 15904 24608 16044
rect 24976 15904 25036 16044
rect 25552 15904 25612 16044
rect 25980 15904 26040 16044
rect 26556 15904 26616 16044
rect 26984 15904 27044 16044
rect 27560 15904 27620 16044
rect 27988 15904 28048 16044
rect 28564 15904 28624 16044
rect 28992 15904 29052 16044
rect 29568 15904 29628 16044
rect 29996 15904 30056 16044
rect 30572 15904 30632 16044
rect 31000 15904 31060 16044
rect 31576 15904 31636 16044
rect 32004 15904 32064 16044
rect 32580 15904 32640 16044
rect 33008 15904 33068 16044
rect 33584 15904 33644 16044
rect 34012 15904 34072 16044
rect 34588 15904 34648 16044
rect 2736 15730 2774 15790
rect 3638 15730 3778 15790
rect 4642 15730 4782 15790
rect 5646 15730 5786 15790
rect 6650 15730 6790 15790
rect 7654 15730 7794 15790
rect 8658 15730 8798 15790
rect 9662 15730 9802 15790
rect 10666 15730 10806 15790
rect 11670 15730 11810 15790
rect 12674 15730 12814 15790
rect 13678 15730 13818 15790
rect 14682 15730 14822 15790
rect 15686 15730 15826 15790
rect 16690 15730 16830 15790
rect 17694 15730 17834 15790
rect 18698 15730 18838 15790
rect 19702 15730 19842 15790
rect 20706 15730 20846 15790
rect 21710 15730 21850 15790
rect 22714 15730 22854 15790
rect 23718 15730 23858 15790
rect 24722 15730 24862 15790
rect 25726 15730 25866 15790
rect 26730 15730 26870 15790
rect 27734 15730 27874 15790
rect 28738 15730 28878 15790
rect 29742 15730 29882 15790
rect 30746 15730 30886 15790
rect 31750 15730 31890 15790
rect 32754 15730 32894 15790
rect 33758 15730 33898 15790
rect 34762 15730 34796 15790
rect 2736 15154 2774 15214
rect 3638 15154 3778 15214
rect 4642 15154 4782 15214
rect 5646 15154 5786 15214
rect 6650 15154 6790 15214
rect 7654 15154 7794 15214
rect 8658 15154 8798 15214
rect 9662 15154 9802 15214
rect 10666 15154 10806 15214
rect 11670 15154 11810 15214
rect 12674 15154 12814 15214
rect 13678 15154 13818 15214
rect 14682 15154 14822 15214
rect 15686 15154 15826 15214
rect 16690 15154 16830 15214
rect 17694 15154 17834 15214
rect 18698 15154 18838 15214
rect 19702 15154 19842 15214
rect 20706 15154 20846 15214
rect 21710 15154 21850 15214
rect 22714 15154 22854 15214
rect 23718 15154 23858 15214
rect 24722 15154 24862 15214
rect 25726 15154 25866 15214
rect 26730 15154 26870 15214
rect 27734 15154 27874 15214
rect 28738 15154 28878 15214
rect 29742 15154 29882 15214
rect 30746 15154 30886 15214
rect 31750 15154 31890 15214
rect 32754 15154 32894 15214
rect 33758 15154 33898 15214
rect 34762 15154 34796 15214
rect 1046 15071 1067 15142
rect 1138 15071 1162 15142
rect 1233 15071 1271 15142
rect 1342 15071 1366 15142
rect 1437 15071 1460 15142
rect 1046 14138 1460 15071
rect 36064 15142 36478 16075
rect 36064 15071 36085 15142
rect 36156 15071 36180 15142
rect 36251 15071 36289 15142
rect 36360 15071 36384 15142
rect 36455 15071 36478 15142
rect 2888 14900 2948 15040
rect 3464 14900 3524 15040
rect 3892 14900 3952 15040
rect 4468 14900 4528 15040
rect 4896 14900 4956 15040
rect 5472 14900 5532 15040
rect 5900 14900 5960 15040
rect 6476 14900 6536 15040
rect 6904 14900 6964 15040
rect 7480 14900 7540 15040
rect 7908 14900 7968 15040
rect 8484 14900 8544 15040
rect 8912 14900 8972 15040
rect 9488 14900 9548 15040
rect 9916 14900 9976 15040
rect 10492 14900 10552 15040
rect 10920 14900 10980 15040
rect 11496 14900 11556 15040
rect 11924 14900 11984 15040
rect 12500 14900 12560 15040
rect 12928 14900 12988 15040
rect 13504 14900 13564 15040
rect 13932 14900 13992 15040
rect 14508 14900 14568 15040
rect 14936 14900 14996 15040
rect 15512 14900 15572 15040
rect 15940 14900 16000 15040
rect 16516 14900 16576 15040
rect 16944 14900 17004 15040
rect 17520 14900 17580 15040
rect 17948 14900 18008 15040
rect 18524 14900 18584 15040
rect 18952 14900 19012 15040
rect 19528 14900 19588 15040
rect 19956 14900 20016 15040
rect 20532 14900 20592 15040
rect 20960 14900 21020 15040
rect 21536 14900 21596 15040
rect 21964 14900 22024 15040
rect 22540 14900 22600 15040
rect 22968 14900 23028 15040
rect 23544 14900 23604 15040
rect 23972 14900 24032 15040
rect 24548 14900 24608 15040
rect 24976 14900 25036 15040
rect 25552 14900 25612 15040
rect 25980 14900 26040 15040
rect 26556 14900 26616 15040
rect 26984 14900 27044 15040
rect 27560 14900 27620 15040
rect 27988 14900 28048 15040
rect 28564 14900 28624 15040
rect 28992 14900 29052 15040
rect 29568 14900 29628 15040
rect 29996 14900 30056 15040
rect 30572 14900 30632 15040
rect 31000 14900 31060 15040
rect 31576 14900 31636 15040
rect 32004 14900 32064 15040
rect 32580 14900 32640 15040
rect 33008 14900 33068 15040
rect 33584 14900 33644 15040
rect 34012 14900 34072 15040
rect 34588 14900 34648 15040
rect 2736 14726 2774 14786
rect 3638 14726 3778 14786
rect 4642 14726 4782 14786
rect 5646 14726 5786 14786
rect 6650 14726 6790 14786
rect 7654 14726 7794 14786
rect 8658 14726 8798 14786
rect 9662 14726 9802 14786
rect 10666 14726 10806 14786
rect 11670 14726 11810 14786
rect 12674 14726 12814 14786
rect 13678 14726 13818 14786
rect 14682 14726 14822 14786
rect 15686 14726 15826 14786
rect 16690 14726 16830 14786
rect 17694 14726 17834 14786
rect 18698 14726 18838 14786
rect 19702 14726 19842 14786
rect 20706 14726 20846 14786
rect 21710 14726 21850 14786
rect 22714 14726 22854 14786
rect 23718 14726 23858 14786
rect 24722 14726 24862 14786
rect 25726 14726 25866 14786
rect 26730 14726 26870 14786
rect 27734 14726 27874 14786
rect 28738 14726 28878 14786
rect 29742 14726 29882 14786
rect 30746 14726 30886 14786
rect 31750 14726 31890 14786
rect 32754 14726 32894 14786
rect 33758 14726 33898 14786
rect 34762 14726 34796 14786
rect 2736 14150 2774 14210
rect 3638 14150 3778 14210
rect 4642 14150 4782 14210
rect 5646 14150 5786 14210
rect 6650 14150 6790 14210
rect 7654 14150 7794 14210
rect 8658 14150 8798 14210
rect 9662 14150 9802 14210
rect 10666 14150 10806 14210
rect 11670 14150 11810 14210
rect 12674 14150 12814 14210
rect 13678 14150 13818 14210
rect 14682 14150 14822 14210
rect 15686 14150 15826 14210
rect 16690 14150 16830 14210
rect 17694 14150 17834 14210
rect 18698 14150 18838 14210
rect 19702 14150 19842 14210
rect 20706 14150 20846 14210
rect 21710 14150 21850 14210
rect 22714 14150 22854 14210
rect 23718 14150 23858 14210
rect 24722 14150 24862 14210
rect 25726 14150 25866 14210
rect 26730 14150 26870 14210
rect 27734 14150 27874 14210
rect 28738 14150 28878 14210
rect 29742 14150 29882 14210
rect 30746 14150 30886 14210
rect 31750 14150 31890 14210
rect 32754 14150 32894 14210
rect 33758 14150 33898 14210
rect 34762 14150 34796 14210
rect 1046 14067 1067 14138
rect 1138 14067 1162 14138
rect 1233 14067 1271 14138
rect 1342 14067 1366 14138
rect 1437 14067 1460 14138
rect 1046 13134 1460 14067
rect 36064 14138 36478 15071
rect 36064 14067 36085 14138
rect 36156 14067 36180 14138
rect 36251 14067 36289 14138
rect 36360 14067 36384 14138
rect 36455 14067 36478 14138
rect 2888 13896 2948 14036
rect 3464 13896 3524 14036
rect 3892 13896 3952 14036
rect 4468 13896 4528 14036
rect 4896 13896 4956 14036
rect 5472 13896 5532 14036
rect 5900 13896 5960 14036
rect 6476 13896 6536 14036
rect 6904 13896 6964 14036
rect 7480 13896 7540 14036
rect 7908 13896 7968 14036
rect 8484 13896 8544 14036
rect 8912 13896 8972 14036
rect 9488 13896 9548 14036
rect 9916 13896 9976 14036
rect 10492 13896 10552 14036
rect 10920 13896 10980 14036
rect 11496 13896 11556 14036
rect 11924 13896 11984 14036
rect 12500 13896 12560 14036
rect 12928 13896 12988 14036
rect 13504 13896 13564 14036
rect 13932 13896 13992 14036
rect 14508 13896 14568 14036
rect 14936 13896 14996 14036
rect 15512 13896 15572 14036
rect 15940 13896 16000 14036
rect 16516 13896 16576 14036
rect 16944 13896 17004 14036
rect 17520 13896 17580 14036
rect 17948 13896 18008 14036
rect 18524 13896 18584 14036
rect 18952 13896 19012 14036
rect 19528 13896 19588 14036
rect 19956 13896 20016 14036
rect 20532 13896 20592 14036
rect 20960 13896 21020 14036
rect 21536 13896 21596 14036
rect 21964 13896 22024 14036
rect 22540 13896 22600 14036
rect 22968 13896 23028 14036
rect 23544 13896 23604 14036
rect 23972 13896 24032 14036
rect 24548 13896 24608 14036
rect 24976 13896 25036 14036
rect 25552 13896 25612 14036
rect 25980 13896 26040 14036
rect 26556 13896 26616 14036
rect 26984 13896 27044 14036
rect 27560 13896 27620 14036
rect 27988 13896 28048 14036
rect 28564 13896 28624 14036
rect 28992 13896 29052 14036
rect 29568 13896 29628 14036
rect 29996 13896 30056 14036
rect 30572 13896 30632 14036
rect 31000 13896 31060 14036
rect 31576 13896 31636 14036
rect 32004 13896 32064 14036
rect 32580 13896 32640 14036
rect 33008 13896 33068 14036
rect 33584 13896 33644 14036
rect 34012 13896 34072 14036
rect 34588 13896 34648 14036
rect 2736 13722 2774 13782
rect 3638 13722 3778 13782
rect 4642 13722 4782 13782
rect 5646 13722 5786 13782
rect 6650 13722 6790 13782
rect 7654 13722 7794 13782
rect 8658 13722 8798 13782
rect 9662 13722 9802 13782
rect 10666 13722 10806 13782
rect 11670 13722 11810 13782
rect 12674 13722 12814 13782
rect 13678 13722 13818 13782
rect 14682 13722 14822 13782
rect 15686 13722 15826 13782
rect 16690 13722 16830 13782
rect 17694 13722 17834 13782
rect 18698 13722 18838 13782
rect 19702 13722 19842 13782
rect 20706 13722 20846 13782
rect 21710 13722 21850 13782
rect 22714 13722 22854 13782
rect 23718 13722 23858 13782
rect 24722 13722 24862 13782
rect 25726 13722 25866 13782
rect 26730 13722 26870 13782
rect 27734 13722 27874 13782
rect 28738 13722 28878 13782
rect 29742 13722 29882 13782
rect 30746 13722 30886 13782
rect 31750 13722 31890 13782
rect 32754 13722 32894 13782
rect 33758 13722 33898 13782
rect 34762 13722 34796 13782
rect 2736 13146 2774 13206
rect 3638 13146 3778 13206
rect 4642 13146 4782 13206
rect 5646 13146 5786 13206
rect 6650 13146 6790 13206
rect 7654 13146 7794 13206
rect 8658 13146 8798 13206
rect 9662 13146 9802 13206
rect 10666 13146 10806 13206
rect 11670 13146 11810 13206
rect 12674 13146 12814 13206
rect 13678 13146 13818 13206
rect 14682 13146 14822 13206
rect 15686 13146 15826 13206
rect 16690 13146 16830 13206
rect 17694 13146 17834 13206
rect 18698 13146 18838 13206
rect 19702 13146 19842 13206
rect 20706 13146 20846 13206
rect 21710 13146 21850 13206
rect 22714 13146 22854 13206
rect 23718 13146 23858 13206
rect 24722 13146 24862 13206
rect 25726 13146 25866 13206
rect 26730 13146 26870 13206
rect 27734 13146 27874 13206
rect 28738 13146 28878 13206
rect 29742 13146 29882 13206
rect 30746 13146 30886 13206
rect 31750 13146 31890 13206
rect 32754 13146 32894 13206
rect 33758 13146 33898 13206
rect 34762 13146 34796 13206
rect 1046 13063 1067 13134
rect 1138 13063 1162 13134
rect 1233 13063 1271 13134
rect 1342 13063 1366 13134
rect 1437 13063 1460 13134
rect 1046 12130 1460 13063
rect 36064 13134 36478 14067
rect 36540 18332 36954 18799
rect 41602 18788 42322 18806
rect 41602 18638 41930 18788
rect 42142 18638 42322 18788
rect 41602 18624 42322 18638
rect 36540 18307 37602 18332
rect 36540 18243 37431 18307
rect 37495 18243 37602 18307
rect 41908 18264 42322 18624
rect 36540 18195 37602 18243
rect 36540 18131 37430 18195
rect 37494 18131 37602 18195
rect 36540 18077 37602 18131
rect 41602 18246 42322 18264
rect 41602 18096 41930 18246
rect 42142 18096 42322 18246
rect 41602 18082 42322 18096
rect 36540 18013 37430 18077
rect 37494 18013 37602 18077
rect 36540 17988 37602 18013
rect 36540 17866 36954 17988
rect 36540 17795 36561 17866
rect 36632 17795 36656 17866
rect 36727 17795 36765 17866
rect 36836 17795 36860 17866
rect 36931 17795 36954 17866
rect 36540 16862 36954 17795
rect 41908 17708 42322 18082
rect 41602 17690 42322 17708
rect 41602 17540 41930 17690
rect 42142 17540 42322 17690
rect 41602 17526 42322 17540
rect 36540 16791 36561 16862
rect 36632 16791 36656 16862
rect 36727 16791 36765 16862
rect 36836 16791 36860 16862
rect 36931 16791 36954 16862
rect 36540 15858 36954 16791
rect 37394 16650 37602 16680
rect 37394 16586 37423 16650
rect 37487 16586 37602 16650
rect 37394 16558 37602 16586
rect 37394 16494 37423 16558
rect 37487 16494 37602 16558
rect 37394 16467 37602 16494
rect 37394 16403 37423 16467
rect 37487 16403 37602 16467
rect 37394 16381 37602 16403
rect 41602 16545 41847 16558
rect 41602 16388 41707 16545
rect 41821 16388 41847 16545
rect 41602 16374 41847 16388
rect 36540 15787 36561 15858
rect 36632 15787 36656 15858
rect 36727 15787 36765 15858
rect 36836 15787 36860 15858
rect 36931 15787 36954 15858
rect 36540 14854 36954 15787
rect 41602 15655 41847 15668
rect 41602 15498 41707 15655
rect 41821 15498 41847 15655
rect 41602 15484 41847 15498
rect 36540 14783 36561 14854
rect 36632 14783 36656 14854
rect 36727 14783 36765 14854
rect 36836 14783 36860 14854
rect 36931 14783 36954 14854
rect 41908 14806 42322 17526
rect 36540 14332 36954 14783
rect 41602 14788 42322 14806
rect 41602 14638 41930 14788
rect 42142 14638 42322 14788
rect 41602 14624 42322 14638
rect 36540 14307 37602 14332
rect 36540 14243 37431 14307
rect 37495 14243 37602 14307
rect 41908 14264 42322 14624
rect 36540 14195 37602 14243
rect 36540 14131 37430 14195
rect 37494 14131 37602 14195
rect 36540 14077 37602 14131
rect 41602 14246 42322 14264
rect 41602 14096 41930 14246
rect 42142 14096 42322 14246
rect 41602 14082 42322 14096
rect 36540 14013 37430 14077
rect 37494 14013 37602 14077
rect 36540 13988 37602 14013
rect 36540 13850 36954 13988
rect 36540 13779 36561 13850
rect 36632 13779 36656 13850
rect 36727 13779 36765 13850
rect 36836 13779 36860 13850
rect 36931 13779 36954 13850
rect 36540 13636 36954 13779
rect 41908 13708 42322 14082
rect 36538 13356 36954 13636
rect 41602 13690 42322 13708
rect 41602 13540 41930 13690
rect 42142 13540 42322 13690
rect 41602 13526 42322 13540
rect 36064 13063 36085 13134
rect 36156 13063 36180 13134
rect 36251 13063 36289 13134
rect 36360 13063 36384 13134
rect 36455 13063 36478 13134
rect 2888 12892 2948 13032
rect 3464 12892 3524 13032
rect 3892 12892 3952 13032
rect 4468 12892 4528 13032
rect 4896 12892 4956 13032
rect 5472 12892 5532 13032
rect 5900 12892 5960 13032
rect 6476 12892 6536 13032
rect 6904 12892 6964 13032
rect 7480 12892 7540 13032
rect 7908 12892 7968 13032
rect 8484 12892 8544 13032
rect 8912 12892 8972 13032
rect 9488 12892 9548 13032
rect 9916 12892 9976 13032
rect 10492 12892 10552 13032
rect 10920 12892 10980 13032
rect 11496 12892 11556 13032
rect 11924 12892 11984 13032
rect 12500 12892 12560 13032
rect 12928 12892 12988 13032
rect 13504 12892 13564 13032
rect 13932 12892 13992 13032
rect 14508 12892 14568 13032
rect 14936 12892 14996 13032
rect 15512 12892 15572 13032
rect 15940 12892 16000 13032
rect 16516 12892 16576 13032
rect 16944 12892 17004 13032
rect 17520 12892 17580 13032
rect 17948 12892 18008 13032
rect 18524 12892 18584 13032
rect 18952 12892 19012 13032
rect 19528 12892 19588 13032
rect 19956 12892 20016 13032
rect 20532 12892 20592 13032
rect 20960 12892 21020 13032
rect 21536 12892 21596 13032
rect 21964 12892 22024 13032
rect 22540 12892 22600 13032
rect 22968 12892 23028 13032
rect 23544 12892 23604 13032
rect 23972 12892 24032 13032
rect 24548 12892 24608 13032
rect 24976 12892 25036 13032
rect 25552 12892 25612 13032
rect 25980 12892 26040 13032
rect 26556 12892 26616 13032
rect 26984 12892 27044 13032
rect 27560 12892 27620 13032
rect 27988 12892 28048 13032
rect 28564 12892 28624 13032
rect 28992 12892 29052 13032
rect 29568 12892 29628 13032
rect 29996 12892 30056 13032
rect 30572 12892 30632 13032
rect 31000 12892 31060 13032
rect 31576 12892 31636 13032
rect 32004 12892 32064 13032
rect 32580 12892 32640 13032
rect 33008 12892 33068 13032
rect 33584 12892 33644 13032
rect 34012 12892 34072 13032
rect 34588 12892 34648 13032
rect 2736 12718 2774 12778
rect 3638 12718 3778 12778
rect 4642 12718 4782 12778
rect 5646 12718 5786 12778
rect 6650 12718 6790 12778
rect 7654 12718 7794 12778
rect 8658 12718 8798 12778
rect 9662 12718 9802 12778
rect 10666 12718 10806 12778
rect 11670 12718 11810 12778
rect 12674 12718 12814 12778
rect 13678 12718 13818 12778
rect 14682 12718 14822 12778
rect 15686 12718 15826 12778
rect 16690 12718 16830 12778
rect 17694 12718 17834 12778
rect 18698 12718 18838 12778
rect 19702 12718 19842 12778
rect 20706 12718 20846 12778
rect 21710 12718 21850 12778
rect 22714 12718 22854 12778
rect 23718 12718 23858 12778
rect 24722 12718 24862 12778
rect 25726 12718 25866 12778
rect 26730 12718 26870 12778
rect 27734 12718 27874 12778
rect 28738 12718 28878 12778
rect 29742 12718 29882 12778
rect 30746 12718 30886 12778
rect 31750 12718 31890 12778
rect 32754 12718 32894 12778
rect 33758 12718 33898 12778
rect 34762 12718 34796 12778
rect 36064 12594 36478 13063
rect 36064 12530 36094 12594
rect 36158 12530 36190 12594
rect 36254 12530 36286 12594
rect 36350 12530 36382 12594
rect 36446 12530 36478 12594
rect 36064 12503 36478 12530
rect 36064 12439 36094 12503
rect 36158 12439 36190 12503
rect 36254 12439 36286 12503
rect 36350 12439 36382 12503
rect 36446 12439 36478 12503
rect 36064 12412 36478 12439
rect 36064 12348 36094 12412
rect 36158 12348 36190 12412
rect 36254 12348 36286 12412
rect 36350 12348 36382 12412
rect 36446 12348 36478 12412
rect 2736 12142 2774 12202
rect 3638 12142 3778 12202
rect 4642 12142 4782 12202
rect 5646 12142 5786 12202
rect 6650 12142 6790 12202
rect 7654 12142 7794 12202
rect 8658 12142 8798 12202
rect 9662 12142 9802 12202
rect 10666 12142 10806 12202
rect 11670 12142 11810 12202
rect 12674 12142 12814 12202
rect 13678 12142 13818 12202
rect 14682 12142 14822 12202
rect 15686 12142 15826 12202
rect 16690 12142 16830 12202
rect 17694 12142 17834 12202
rect 18698 12142 18838 12202
rect 19702 12142 19842 12202
rect 20706 12142 20846 12202
rect 21710 12142 21850 12202
rect 22714 12142 22854 12202
rect 23718 12142 23858 12202
rect 24722 12142 24862 12202
rect 25726 12142 25866 12202
rect 26730 12142 26870 12202
rect 27734 12142 27874 12202
rect 28738 12142 28878 12202
rect 29742 12142 29882 12202
rect 30746 12142 30886 12202
rect 31750 12142 31890 12202
rect 32754 12142 32894 12202
rect 33758 12142 33898 12202
rect 34762 12142 34796 12202
rect 1046 12059 1067 12130
rect 1138 12059 1162 12130
rect 1233 12059 1271 12130
rect 1342 12059 1366 12130
rect 1437 12059 1460 12130
rect 1046 11126 1460 12059
rect 36064 12130 36478 12348
rect 36064 12059 36085 12130
rect 36156 12059 36180 12130
rect 36251 12059 36289 12130
rect 36360 12059 36384 12130
rect 36455 12059 36478 12130
rect 2888 11888 2948 12028
rect 3464 11888 3524 12028
rect 3892 11888 3952 12028
rect 4468 11888 4528 12028
rect 4896 11888 4956 12028
rect 5472 11888 5532 12028
rect 5900 11888 5960 12028
rect 6476 11888 6536 12028
rect 6904 11888 6964 12028
rect 7480 11888 7540 12028
rect 7908 11888 7968 12028
rect 8484 11888 8544 12028
rect 8912 11888 8972 12028
rect 9488 11888 9548 12028
rect 9916 11888 9976 12028
rect 10492 11888 10552 12028
rect 10920 11888 10980 12028
rect 11496 11888 11556 12028
rect 11924 11888 11984 12028
rect 12500 11888 12560 12028
rect 12928 11888 12988 12028
rect 13504 11888 13564 12028
rect 13932 11888 13992 12028
rect 14508 11888 14568 12028
rect 14936 11888 14996 12028
rect 15512 11888 15572 12028
rect 15940 11888 16000 12028
rect 16516 11888 16576 12028
rect 16944 11888 17004 12028
rect 17520 11888 17580 12028
rect 17948 11888 18008 12028
rect 18524 11888 18584 12028
rect 18952 11888 19012 12028
rect 19528 11888 19588 12028
rect 19956 11888 20016 12028
rect 20532 11888 20592 12028
rect 20960 11888 21020 12028
rect 21536 11888 21596 12028
rect 21964 11888 22024 12028
rect 22540 11888 22600 12028
rect 22968 11888 23028 12028
rect 23544 11888 23604 12028
rect 23972 11888 24032 12028
rect 24548 11888 24608 12028
rect 24976 11888 25036 12028
rect 25552 11888 25612 12028
rect 25980 11888 26040 12028
rect 26556 11888 26616 12028
rect 26984 11888 27044 12028
rect 27560 11888 27620 12028
rect 27988 11888 28048 12028
rect 28564 11888 28624 12028
rect 28992 11888 29052 12028
rect 29568 11888 29628 12028
rect 29996 11888 30056 12028
rect 30572 11888 30632 12028
rect 31000 11888 31060 12028
rect 31576 11888 31636 12028
rect 32004 11888 32064 12028
rect 32580 11888 32640 12028
rect 33008 11888 33068 12028
rect 33584 11888 33644 12028
rect 34012 11888 34072 12028
rect 34588 11888 34648 12028
rect 2736 11714 2774 11774
rect 3638 11714 3778 11774
rect 4642 11714 4782 11774
rect 5646 11714 5786 11774
rect 6650 11714 6790 11774
rect 7654 11714 7794 11774
rect 8658 11714 8798 11774
rect 9662 11714 9802 11774
rect 10666 11714 10806 11774
rect 11670 11714 11810 11774
rect 12674 11714 12814 11774
rect 13678 11714 13818 11774
rect 14682 11714 14822 11774
rect 15686 11714 15826 11774
rect 16690 11714 16830 11774
rect 17694 11714 17834 11774
rect 18698 11714 18838 11774
rect 19702 11714 19842 11774
rect 20706 11714 20846 11774
rect 21710 11714 21850 11774
rect 22714 11714 22854 11774
rect 23718 11714 23858 11774
rect 24722 11714 24862 11774
rect 25726 11714 25866 11774
rect 26730 11714 26870 11774
rect 27734 11714 27874 11774
rect 28738 11714 28878 11774
rect 29742 11714 29882 11774
rect 30746 11714 30886 11774
rect 31750 11714 31890 11774
rect 32754 11714 32894 11774
rect 33758 11714 33898 11774
rect 34762 11714 34796 11774
rect 2736 11138 2774 11198
rect 3638 11138 3778 11198
rect 4642 11138 4782 11198
rect 5646 11138 5786 11198
rect 6650 11138 6790 11198
rect 7654 11138 7794 11198
rect 8658 11138 8798 11198
rect 9662 11138 9802 11198
rect 10666 11138 10806 11198
rect 11670 11138 11810 11198
rect 12674 11138 12814 11198
rect 13678 11138 13818 11198
rect 14682 11138 14822 11198
rect 15686 11138 15826 11198
rect 16690 11138 16830 11198
rect 17694 11138 17834 11198
rect 18698 11138 18838 11198
rect 19702 11138 19842 11198
rect 20706 11138 20846 11198
rect 21710 11138 21850 11198
rect 22714 11138 22854 11198
rect 23718 11138 23858 11198
rect 24722 11138 24862 11198
rect 25726 11138 25866 11198
rect 26730 11138 26870 11198
rect 27734 11138 27874 11198
rect 28738 11138 28878 11198
rect 29742 11138 29882 11198
rect 30746 11138 30886 11198
rect 31750 11138 31890 11198
rect 32754 11138 32894 11198
rect 33758 11138 33898 11198
rect 34762 11138 34796 11198
rect 1046 11055 1067 11126
rect 1138 11055 1162 11126
rect 1233 11055 1271 11126
rect 1342 11055 1366 11126
rect 1437 11055 1460 11126
rect 1046 10122 1460 11055
rect 36064 11126 36478 12059
rect 36064 11055 36085 11126
rect 36156 11055 36180 11126
rect 36251 11055 36289 11126
rect 36360 11055 36384 11126
rect 36455 11055 36478 11126
rect 2888 10884 2948 11024
rect 3464 10884 3524 11024
rect 3892 10884 3952 11024
rect 4468 10884 4528 11024
rect 4896 10884 4956 11024
rect 5472 10884 5532 11024
rect 5900 10884 5960 11024
rect 6476 10884 6536 11024
rect 6904 10884 6964 11024
rect 7480 10884 7540 11024
rect 7908 10884 7968 11024
rect 8484 10884 8544 11024
rect 8912 10884 8972 11024
rect 9488 10884 9548 11024
rect 9916 10884 9976 11024
rect 10492 10884 10552 11024
rect 10920 10884 10980 11024
rect 11496 10884 11556 11024
rect 11924 10884 11984 11024
rect 12500 10884 12560 11024
rect 12928 10884 12988 11024
rect 13504 10884 13564 11024
rect 13932 10884 13992 11024
rect 14508 10884 14568 11024
rect 14936 10884 14996 11024
rect 15512 10884 15572 11024
rect 15940 10884 16000 11024
rect 16516 10884 16576 11024
rect 16944 10884 17004 11024
rect 17520 10884 17580 11024
rect 17948 10884 18008 11024
rect 18524 10884 18584 11024
rect 18952 10884 19012 11024
rect 19528 10884 19588 11024
rect 19956 10884 20016 11024
rect 20532 10884 20592 11024
rect 20960 10884 21020 11024
rect 21536 10884 21596 11024
rect 21964 10884 22024 11024
rect 22540 10884 22600 11024
rect 22968 10884 23028 11024
rect 23544 10884 23604 11024
rect 23972 10884 24032 11024
rect 24548 10884 24608 11024
rect 24976 10884 25036 11024
rect 25552 10884 25612 11024
rect 25980 10884 26040 11024
rect 26556 10884 26616 11024
rect 26984 10884 27044 11024
rect 27560 10884 27620 11024
rect 27988 10884 28048 11024
rect 28564 10884 28624 11024
rect 28992 10884 29052 11024
rect 29568 10884 29628 11024
rect 29996 10884 30056 11024
rect 30572 10884 30632 11024
rect 31000 10884 31060 11024
rect 31576 10884 31636 11024
rect 32004 10884 32064 11024
rect 32580 10884 32640 11024
rect 33008 10884 33068 11024
rect 33584 10884 33644 11024
rect 34012 10884 34072 11024
rect 34588 10884 34648 11024
rect 2736 10710 2774 10770
rect 3638 10710 3778 10770
rect 4642 10710 4782 10770
rect 5646 10710 5786 10770
rect 6650 10710 6790 10770
rect 7654 10710 7794 10770
rect 8658 10710 8798 10770
rect 9662 10710 9802 10770
rect 10666 10710 10806 10770
rect 11670 10710 11810 10770
rect 12674 10710 12814 10770
rect 13678 10710 13818 10770
rect 14682 10710 14822 10770
rect 15686 10710 15826 10770
rect 16690 10710 16830 10770
rect 17694 10710 17834 10770
rect 18698 10710 18838 10770
rect 19702 10710 19842 10770
rect 20706 10710 20846 10770
rect 21710 10710 21850 10770
rect 22714 10710 22854 10770
rect 23718 10710 23858 10770
rect 24722 10710 24862 10770
rect 25726 10710 25866 10770
rect 26730 10710 26870 10770
rect 27734 10710 27874 10770
rect 28738 10710 28878 10770
rect 29742 10710 29882 10770
rect 30746 10710 30886 10770
rect 31750 10710 31890 10770
rect 32754 10710 32894 10770
rect 33758 10710 33898 10770
rect 34762 10710 34796 10770
rect 2736 10134 2774 10194
rect 3638 10134 3778 10194
rect 4642 10134 4782 10194
rect 5646 10134 5786 10194
rect 6650 10134 6790 10194
rect 7654 10134 7794 10194
rect 8658 10134 8798 10194
rect 9662 10134 9802 10194
rect 10666 10134 10806 10194
rect 11670 10134 11810 10194
rect 12674 10134 12814 10194
rect 13678 10134 13818 10194
rect 14682 10134 14822 10194
rect 15686 10134 15826 10194
rect 16690 10134 16830 10194
rect 17694 10134 17834 10194
rect 18698 10134 18838 10194
rect 19702 10134 19842 10194
rect 20706 10134 20846 10194
rect 21710 10134 21850 10194
rect 22714 10134 22854 10194
rect 23718 10134 23858 10194
rect 24722 10134 24862 10194
rect 25726 10134 25866 10194
rect 26730 10134 26870 10194
rect 27734 10134 27874 10194
rect 28738 10134 28878 10194
rect 29742 10134 29882 10194
rect 30746 10134 30886 10194
rect 31750 10134 31890 10194
rect 32754 10134 32894 10194
rect 33758 10134 33898 10194
rect 34762 10134 34796 10194
rect 1046 10051 1067 10122
rect 1138 10051 1162 10122
rect 1233 10051 1271 10122
rect 1342 10051 1366 10122
rect 1437 10051 1460 10122
rect 1046 9118 1460 10051
rect 36064 10122 36478 11055
rect 36064 10051 36085 10122
rect 36156 10051 36180 10122
rect 36251 10051 36289 10122
rect 36360 10051 36384 10122
rect 36455 10051 36478 10122
rect 2888 9880 2948 10020
rect 3464 9880 3524 10020
rect 3892 9880 3952 10020
rect 4468 9880 4528 10020
rect 4896 9880 4956 10020
rect 5472 9880 5532 10020
rect 5900 9880 5960 10020
rect 6476 9880 6536 10020
rect 6904 9880 6964 10020
rect 7480 9880 7540 10020
rect 7908 9880 7968 10020
rect 8484 9880 8544 10020
rect 8912 9880 8972 10020
rect 9488 9880 9548 10020
rect 9916 9880 9976 10020
rect 10492 9880 10552 10020
rect 10920 9880 10980 10020
rect 11496 9880 11556 10020
rect 11924 9880 11984 10020
rect 12500 9880 12560 10020
rect 12928 9880 12988 10020
rect 13504 9880 13564 10020
rect 13932 9880 13992 10020
rect 14508 9880 14568 10020
rect 14936 9880 14996 10020
rect 15512 9880 15572 10020
rect 15940 9880 16000 10020
rect 16516 9880 16576 10020
rect 16944 9880 17004 10020
rect 17520 9880 17580 10020
rect 17948 9880 18008 10020
rect 18524 9880 18584 10020
rect 18952 9880 19012 10020
rect 19528 9880 19588 10020
rect 19956 9880 20016 10020
rect 20532 9880 20592 10020
rect 20960 9880 21020 10020
rect 21536 9880 21596 10020
rect 21964 9880 22024 10020
rect 22540 9880 22600 10020
rect 22968 9880 23028 10020
rect 23544 9880 23604 10020
rect 23972 9880 24032 10020
rect 24548 9880 24608 10020
rect 24976 9880 25036 10020
rect 25552 9880 25612 10020
rect 25980 9880 26040 10020
rect 26556 9880 26616 10020
rect 26984 9880 27044 10020
rect 27560 9880 27620 10020
rect 27988 9880 28048 10020
rect 28564 9880 28624 10020
rect 28992 9880 29052 10020
rect 29568 9880 29628 10020
rect 29996 9880 30056 10020
rect 30572 9880 30632 10020
rect 31000 9880 31060 10020
rect 31576 9880 31636 10020
rect 32004 9880 32064 10020
rect 32580 9880 32640 10020
rect 33008 9880 33068 10020
rect 33584 9880 33644 10020
rect 34012 9880 34072 10020
rect 34588 9880 34648 10020
rect 2736 9706 2774 9766
rect 3638 9706 3778 9766
rect 4642 9706 4782 9766
rect 5646 9706 5786 9766
rect 6650 9706 6790 9766
rect 7654 9706 7794 9766
rect 8658 9706 8798 9766
rect 9662 9706 9802 9766
rect 10666 9706 10806 9766
rect 11670 9706 11810 9766
rect 12674 9706 12814 9766
rect 13678 9706 13818 9766
rect 14682 9706 14822 9766
rect 15686 9706 15826 9766
rect 16690 9706 16830 9766
rect 17694 9706 17834 9766
rect 18698 9706 18838 9766
rect 19702 9706 19842 9766
rect 20706 9706 20846 9766
rect 21710 9706 21850 9766
rect 22714 9706 22854 9766
rect 23718 9706 23858 9766
rect 24722 9706 24862 9766
rect 25726 9706 25866 9766
rect 26730 9706 26870 9766
rect 27734 9706 27874 9766
rect 28738 9706 28878 9766
rect 29742 9706 29882 9766
rect 30746 9706 30886 9766
rect 31750 9706 31890 9766
rect 32754 9706 32894 9766
rect 33758 9706 33898 9766
rect 34762 9706 34796 9766
rect 2736 9130 2774 9190
rect 3638 9130 3778 9190
rect 4642 9130 4782 9190
rect 5646 9130 5786 9190
rect 6650 9130 6790 9190
rect 7654 9130 7794 9190
rect 8658 9130 8798 9190
rect 9662 9130 9802 9190
rect 10666 9130 10806 9190
rect 11670 9130 11810 9190
rect 12674 9130 12814 9190
rect 13678 9130 13818 9190
rect 14682 9130 14822 9190
rect 15686 9130 15826 9190
rect 16690 9130 16830 9190
rect 17694 9130 17834 9190
rect 18698 9130 18838 9190
rect 19702 9130 19842 9190
rect 20706 9130 20846 9190
rect 21710 9130 21850 9190
rect 22714 9130 22854 9190
rect 23718 9130 23858 9190
rect 24722 9130 24862 9190
rect 25726 9130 25866 9190
rect 26730 9130 26870 9190
rect 27734 9130 27874 9190
rect 28738 9130 28878 9190
rect 29742 9130 29882 9190
rect 30746 9130 30886 9190
rect 31750 9130 31890 9190
rect 32754 9130 32894 9190
rect 33758 9130 33898 9190
rect 34762 9130 34796 9190
rect 1046 9047 1067 9118
rect 1138 9047 1162 9118
rect 1233 9047 1271 9118
rect 1342 9047 1366 9118
rect 1437 9047 1460 9118
rect 1046 8114 1460 9047
rect 36064 9118 36478 10051
rect 36064 9047 36085 9118
rect 36156 9047 36180 9118
rect 36251 9047 36289 9118
rect 36360 9047 36384 9118
rect 36455 9047 36478 9118
rect 2888 8876 2948 9016
rect 3464 8876 3524 9016
rect 3892 8876 3952 9016
rect 4468 8876 4528 9016
rect 4896 8876 4956 9016
rect 5472 8876 5532 9016
rect 5900 8876 5960 9016
rect 6476 8876 6536 9016
rect 6904 8876 6964 9016
rect 7480 8876 7540 9016
rect 7908 8876 7968 9016
rect 8484 8876 8544 9016
rect 8912 8876 8972 9016
rect 9488 8876 9548 9016
rect 9916 8876 9976 9016
rect 10492 8876 10552 9016
rect 10920 8876 10980 9016
rect 11496 8876 11556 9016
rect 11924 8876 11984 9016
rect 12500 8876 12560 9016
rect 12928 8876 12988 9016
rect 13504 8876 13564 9016
rect 13932 8876 13992 9016
rect 14508 8876 14568 9016
rect 14936 8876 14996 9016
rect 15512 8876 15572 9016
rect 15940 8876 16000 9016
rect 16516 8876 16576 9016
rect 16944 8876 17004 9016
rect 17520 8876 17580 9016
rect 17948 8876 18008 9016
rect 18524 8876 18584 9016
rect 18952 8876 19012 9016
rect 19528 8876 19588 9016
rect 19956 8876 20016 9016
rect 20532 8876 20592 9016
rect 20960 8876 21020 9016
rect 21536 8876 21596 9016
rect 21964 8876 22024 9016
rect 22540 8876 22600 9016
rect 22968 8876 23028 9016
rect 23544 8876 23604 9016
rect 23972 8876 24032 9016
rect 24548 8876 24608 9016
rect 24976 8876 25036 9016
rect 25552 8876 25612 9016
rect 25980 8876 26040 9016
rect 26556 8876 26616 9016
rect 26984 8876 27044 9016
rect 27560 8876 27620 9016
rect 27988 8876 28048 9016
rect 28564 8876 28624 9016
rect 28992 8876 29052 9016
rect 29568 8876 29628 9016
rect 29996 8876 30056 9016
rect 30572 8876 30632 9016
rect 31000 8876 31060 9016
rect 31576 8876 31636 9016
rect 32004 8876 32064 9016
rect 32580 8876 32640 9016
rect 33008 8876 33068 9016
rect 33584 8876 33644 9016
rect 34012 8876 34072 9016
rect 34588 8876 34648 9016
rect 2736 8702 2774 8762
rect 3638 8702 3778 8762
rect 4642 8702 4782 8762
rect 5646 8702 5786 8762
rect 6650 8702 6790 8762
rect 7654 8702 7794 8762
rect 8658 8702 8798 8762
rect 9662 8702 9802 8762
rect 10666 8702 10806 8762
rect 11670 8702 11810 8762
rect 12674 8702 12814 8762
rect 13678 8702 13818 8762
rect 14682 8702 14822 8762
rect 15686 8702 15826 8762
rect 16690 8702 16830 8762
rect 17694 8702 17834 8762
rect 18698 8702 18838 8762
rect 19702 8702 19842 8762
rect 20706 8702 20846 8762
rect 21710 8702 21850 8762
rect 22714 8702 22854 8762
rect 23718 8702 23858 8762
rect 24722 8702 24862 8762
rect 25726 8702 25866 8762
rect 26730 8702 26870 8762
rect 27734 8702 27874 8762
rect 28738 8702 28878 8762
rect 29742 8702 29882 8762
rect 30746 8702 30886 8762
rect 31750 8702 31890 8762
rect 32754 8702 32894 8762
rect 33758 8702 33898 8762
rect 34762 8702 34796 8762
rect 36064 8501 36478 9047
rect 36064 8437 36094 8501
rect 36158 8437 36190 8501
rect 36254 8437 36286 8501
rect 36350 8437 36382 8501
rect 36446 8437 36478 8501
rect 36064 8410 36478 8437
rect 36064 8346 36094 8410
rect 36158 8346 36190 8410
rect 36254 8346 36286 8410
rect 36350 8346 36382 8410
rect 36446 8346 36478 8410
rect 36064 8319 36478 8346
rect 36064 8255 36094 8319
rect 36158 8255 36190 8319
rect 36254 8255 36286 8319
rect 36350 8255 36382 8319
rect 36446 8255 36478 8319
rect 2736 8126 2774 8186
rect 3638 8126 3778 8186
rect 4642 8126 4782 8186
rect 5646 8126 5786 8186
rect 6650 8126 6790 8186
rect 7654 8126 7794 8186
rect 8658 8126 8798 8186
rect 9662 8126 9802 8186
rect 10666 8126 10806 8186
rect 11670 8126 11810 8186
rect 12674 8126 12814 8186
rect 13678 8126 13818 8186
rect 14682 8126 14822 8186
rect 15686 8126 15826 8186
rect 16690 8126 16830 8186
rect 17694 8126 17834 8186
rect 18698 8126 18838 8186
rect 19702 8126 19842 8186
rect 20706 8126 20846 8186
rect 21710 8126 21850 8186
rect 22714 8126 22854 8186
rect 23718 8126 23858 8186
rect 24722 8126 24862 8186
rect 25726 8126 25866 8186
rect 26730 8126 26870 8186
rect 27734 8126 27874 8186
rect 28738 8126 28878 8186
rect 29742 8126 29882 8186
rect 30746 8126 30886 8186
rect 31750 8126 31890 8186
rect 32754 8126 32894 8186
rect 33758 8126 33898 8186
rect 34762 8126 34796 8186
rect 1046 8043 1067 8114
rect 1138 8043 1162 8114
rect 1233 8043 1271 8114
rect 1342 8043 1366 8114
rect 1437 8043 1460 8114
rect 1046 7110 1460 8043
rect 36064 8114 36478 8255
rect 36064 8043 36085 8114
rect 36156 8043 36180 8114
rect 36251 8043 36289 8114
rect 36360 8043 36384 8114
rect 36455 8043 36478 8114
rect 2888 7872 2948 8012
rect 3464 7872 3524 8012
rect 3892 7872 3952 8012
rect 4468 7872 4528 8012
rect 4896 7872 4956 8012
rect 5472 7872 5532 8012
rect 5900 7872 5960 8012
rect 6476 7872 6536 8012
rect 6904 7872 6964 8012
rect 7480 7872 7540 8012
rect 7908 7872 7968 8012
rect 8484 7872 8544 8012
rect 8912 7872 8972 8012
rect 9488 7872 9548 8012
rect 9916 7872 9976 8012
rect 10492 7872 10552 8012
rect 10920 7872 10980 8012
rect 11496 7872 11556 8012
rect 11924 7872 11984 8012
rect 12500 7872 12560 8012
rect 12928 7872 12988 8012
rect 13504 7872 13564 8012
rect 13932 7872 13992 8012
rect 14508 7872 14568 8012
rect 14936 7872 14996 8012
rect 15512 7872 15572 8012
rect 15940 7872 16000 8012
rect 16516 7872 16576 8012
rect 16944 7872 17004 8012
rect 17520 7872 17580 8012
rect 17948 7872 18008 8012
rect 18524 7872 18584 8012
rect 18952 7872 19012 8012
rect 19528 7872 19588 8012
rect 19956 7872 20016 8012
rect 20532 7872 20592 8012
rect 20960 7872 21020 8012
rect 21536 7872 21596 8012
rect 21964 7872 22024 8012
rect 22540 7872 22600 8012
rect 22968 7872 23028 8012
rect 23544 7872 23604 8012
rect 23972 7872 24032 8012
rect 24548 7872 24608 8012
rect 24976 7872 25036 8012
rect 25552 7872 25612 8012
rect 25980 7872 26040 8012
rect 26556 7872 26616 8012
rect 26984 7872 27044 8012
rect 27560 7872 27620 8012
rect 27988 7872 28048 8012
rect 28564 7872 28624 8012
rect 28992 7872 29052 8012
rect 29568 7872 29628 8012
rect 29996 7872 30056 8012
rect 30572 7872 30632 8012
rect 31000 7872 31060 8012
rect 31576 7872 31636 8012
rect 32004 7872 32064 8012
rect 32580 7872 32640 8012
rect 33008 7872 33068 8012
rect 33584 7872 33644 8012
rect 34012 7872 34072 8012
rect 34588 7872 34648 8012
rect 2736 7698 2774 7758
rect 3638 7698 3778 7758
rect 4642 7698 4782 7758
rect 5646 7698 5786 7758
rect 6650 7698 6790 7758
rect 7654 7698 7794 7758
rect 8658 7698 8798 7758
rect 9662 7698 9802 7758
rect 10666 7698 10806 7758
rect 11670 7698 11810 7758
rect 12674 7698 12814 7758
rect 13678 7698 13818 7758
rect 14682 7698 14822 7758
rect 15686 7698 15826 7758
rect 16690 7698 16830 7758
rect 17694 7698 17834 7758
rect 18698 7698 18838 7758
rect 19702 7698 19842 7758
rect 20706 7698 20846 7758
rect 21710 7698 21850 7758
rect 22714 7698 22854 7758
rect 23718 7698 23858 7758
rect 24722 7698 24862 7758
rect 25726 7698 25866 7758
rect 26730 7698 26870 7758
rect 27734 7698 27874 7758
rect 28738 7698 28878 7758
rect 29742 7698 29882 7758
rect 30746 7698 30886 7758
rect 31750 7698 31890 7758
rect 32754 7698 32894 7758
rect 33758 7698 33898 7758
rect 34762 7698 34796 7758
rect 2736 7122 2774 7182
rect 3638 7122 3778 7182
rect 4642 7122 4782 7182
rect 5646 7122 5786 7182
rect 6650 7122 6790 7182
rect 7654 7122 7794 7182
rect 8658 7122 8798 7182
rect 9662 7122 9802 7182
rect 10666 7122 10806 7182
rect 11670 7122 11810 7182
rect 12674 7122 12814 7182
rect 13678 7122 13818 7182
rect 14682 7122 14822 7182
rect 15686 7122 15826 7182
rect 16690 7122 16830 7182
rect 17694 7122 17834 7182
rect 18698 7122 18838 7182
rect 19702 7122 19842 7182
rect 20706 7122 20846 7182
rect 21710 7122 21850 7182
rect 22714 7122 22854 7182
rect 23718 7122 23858 7182
rect 24722 7122 24862 7182
rect 25726 7122 25866 7182
rect 26730 7122 26870 7182
rect 27734 7122 27874 7182
rect 28738 7122 28878 7182
rect 29742 7122 29882 7182
rect 30746 7122 30886 7182
rect 31750 7122 31890 7182
rect 32754 7122 32894 7182
rect 33758 7122 33898 7182
rect 34762 7122 34796 7182
rect 1046 7039 1067 7110
rect 1138 7039 1162 7110
rect 1233 7039 1271 7110
rect 1342 7039 1366 7110
rect 1437 7039 1460 7110
rect 1046 6106 1460 7039
rect 36064 7110 36478 8043
rect 36540 12846 36954 13356
rect 36540 12775 36561 12846
rect 36632 12775 36656 12846
rect 36727 12775 36765 12846
rect 36836 12775 36860 12846
rect 36931 12775 36954 12846
rect 36540 11842 36954 12775
rect 37394 12592 37602 12622
rect 37394 12528 37423 12592
rect 37487 12528 37602 12592
rect 37394 12500 37602 12528
rect 37394 12436 37423 12500
rect 37487 12436 37602 12500
rect 37394 12409 37602 12436
rect 37394 12345 37423 12409
rect 37487 12345 37602 12409
rect 41602 12545 41847 12558
rect 41602 12388 41707 12545
rect 41821 12388 41847 12545
rect 41602 12374 41847 12388
rect 37394 12323 37602 12345
rect 36540 11771 36561 11842
rect 36632 11771 36656 11842
rect 36727 11771 36765 11842
rect 36836 11771 36860 11842
rect 36931 11771 36954 11842
rect 36540 10838 36954 11771
rect 41602 11655 41847 11668
rect 41602 11498 41707 11655
rect 41821 11498 41847 11655
rect 41602 11484 41847 11498
rect 36540 10767 36561 10838
rect 36632 10767 36656 10838
rect 36727 10767 36765 10838
rect 36836 10767 36860 10838
rect 36931 10767 36954 10838
rect 41908 10806 42322 13526
rect 36540 10332 36954 10767
rect 41602 10788 42322 10806
rect 41602 10638 41930 10788
rect 42142 10638 42322 10788
rect 41602 10624 42322 10638
rect 36540 10307 37602 10332
rect 36540 10243 37431 10307
rect 37495 10243 37602 10307
rect 41908 10264 42322 10624
rect 36540 10195 37602 10243
rect 36540 10131 37430 10195
rect 37494 10131 37602 10195
rect 36540 10077 37602 10131
rect 41602 10246 42322 10264
rect 41602 10096 41930 10246
rect 42142 10096 42322 10246
rect 41602 10082 42322 10096
rect 36540 10013 37430 10077
rect 37494 10013 37602 10077
rect 36540 9988 37602 10013
rect 36540 9834 36954 9988
rect 36540 9763 36561 9834
rect 36632 9763 36656 9834
rect 36727 9763 36765 9834
rect 36836 9763 36860 9834
rect 36931 9763 36954 9834
rect 36540 8830 36954 9763
rect 41908 9708 42322 10082
rect 41602 9690 42322 9708
rect 41602 9540 41930 9690
rect 42142 9540 42322 9690
rect 41602 9526 42322 9540
rect 36540 8759 36561 8830
rect 36632 8759 36656 8830
rect 36727 8759 36765 8830
rect 36836 8759 36860 8830
rect 36931 8759 36954 8830
rect 36540 7826 36954 8759
rect 41602 8545 41847 8558
rect 37394 8499 37602 8529
rect 37394 8435 37423 8499
rect 37487 8435 37602 8499
rect 37394 8407 37602 8435
rect 37394 8343 37423 8407
rect 37487 8343 37602 8407
rect 41602 8388 41707 8545
rect 41821 8388 41847 8545
rect 41602 8374 41847 8388
rect 37394 8316 37602 8343
rect 37394 8252 37423 8316
rect 37487 8252 37602 8316
rect 37394 8230 37602 8252
rect 36540 7755 36561 7826
rect 36632 7755 36656 7826
rect 36727 7755 36765 7826
rect 36836 7755 36860 7826
rect 36931 7755 36954 7826
rect 36540 7620 36954 7755
rect 36538 7340 36954 7620
rect 41602 7655 41847 7668
rect 41602 7498 41707 7655
rect 41821 7498 41847 7655
rect 41602 7484 41847 7498
rect 36064 7039 36085 7110
rect 36156 7039 36180 7110
rect 36251 7039 36289 7110
rect 36360 7039 36384 7110
rect 36455 7039 36478 7110
rect 2888 6868 2948 7008
rect 3464 6868 3524 7008
rect 3892 6868 3952 7008
rect 4468 6868 4528 7008
rect 4896 6868 4956 7008
rect 5472 6868 5532 7008
rect 5900 6868 5960 7008
rect 6476 6868 6536 7008
rect 6904 6868 6964 7008
rect 7480 6868 7540 7008
rect 7908 6868 7968 7008
rect 8484 6868 8544 7008
rect 8912 6868 8972 7008
rect 9488 6868 9548 7008
rect 9916 6868 9976 7008
rect 10492 6868 10552 7008
rect 10920 6868 10980 7008
rect 11496 6868 11556 7008
rect 11924 6868 11984 7008
rect 12500 6868 12560 7008
rect 12928 6868 12988 7008
rect 13504 6868 13564 7008
rect 13932 6868 13992 7008
rect 14508 6868 14568 7008
rect 14936 6868 14996 7008
rect 15512 6868 15572 7008
rect 15940 6868 16000 7008
rect 16516 6868 16576 7008
rect 16944 6868 17004 7008
rect 17520 6868 17580 7008
rect 17948 6868 18008 7008
rect 18524 6868 18584 7008
rect 18952 6868 19012 7008
rect 19528 6868 19588 7008
rect 19956 6868 20016 7008
rect 20532 6868 20592 7008
rect 20960 6868 21020 7008
rect 21536 6868 21596 7008
rect 21964 6868 22024 7008
rect 22540 6868 22600 7008
rect 22968 6868 23028 7008
rect 23544 6868 23604 7008
rect 23972 6868 24032 7008
rect 24548 6868 24608 7008
rect 24976 6868 25036 7008
rect 25552 6868 25612 7008
rect 25980 6868 26040 7008
rect 26556 6868 26616 7008
rect 26984 6868 27044 7008
rect 27560 6868 27620 7008
rect 27988 6868 28048 7008
rect 28564 6868 28624 7008
rect 28992 6868 29052 7008
rect 29568 6868 29628 7008
rect 29996 6868 30056 7008
rect 30572 6868 30632 7008
rect 31000 6868 31060 7008
rect 31576 6868 31636 7008
rect 32004 6868 32064 7008
rect 32580 6868 32640 7008
rect 33008 6868 33068 7008
rect 33584 6868 33644 7008
rect 34012 6868 34072 7008
rect 34588 6868 34648 7008
rect 2736 6694 2774 6754
rect 3638 6694 3778 6754
rect 4642 6694 4782 6754
rect 5646 6694 5786 6754
rect 6650 6694 6790 6754
rect 7654 6694 7794 6754
rect 8658 6694 8798 6754
rect 9662 6694 9802 6754
rect 10666 6694 10806 6754
rect 11670 6694 11810 6754
rect 12674 6694 12814 6754
rect 13678 6694 13818 6754
rect 14682 6694 14822 6754
rect 15686 6694 15826 6754
rect 16690 6694 16830 6754
rect 17694 6694 17834 6754
rect 18698 6694 18838 6754
rect 19702 6694 19842 6754
rect 20706 6694 20846 6754
rect 21710 6694 21850 6754
rect 22714 6694 22854 6754
rect 23718 6694 23858 6754
rect 24722 6694 24862 6754
rect 25726 6694 25866 6754
rect 26730 6694 26870 6754
rect 27734 6694 27874 6754
rect 28738 6694 28878 6754
rect 29742 6694 29882 6754
rect 30746 6694 30886 6754
rect 31750 6694 31890 6754
rect 32754 6694 32894 6754
rect 33758 6694 33898 6754
rect 34762 6694 34796 6754
rect 36064 6576 36478 7039
rect 36540 6822 36954 7340
rect 36540 6751 36561 6822
rect 36632 6751 36656 6822
rect 36727 6751 36765 6822
rect 36836 6751 36860 6822
rect 36931 6751 36954 6822
rect 41908 6806 42322 9526
rect 36064 6294 36480 6576
rect 36540 6330 36954 6751
rect 41602 6788 42322 6806
rect 41602 6638 41930 6788
rect 42142 6638 42322 6788
rect 41602 6624 42322 6638
rect 36540 6305 37602 6330
rect 2736 6118 2774 6178
rect 3638 6118 3778 6178
rect 4642 6118 4782 6178
rect 5646 6118 5786 6178
rect 6650 6118 6790 6178
rect 7654 6118 7794 6178
rect 8658 6118 8798 6178
rect 9662 6118 9802 6178
rect 10666 6118 10806 6178
rect 11670 6118 11810 6178
rect 12674 6118 12814 6178
rect 13678 6118 13818 6178
rect 14682 6118 14822 6178
rect 15686 6118 15826 6178
rect 16690 6118 16830 6178
rect 17694 6118 17834 6178
rect 18698 6118 18838 6178
rect 19702 6118 19842 6178
rect 20706 6118 20846 6178
rect 21710 6118 21850 6178
rect 22714 6118 22854 6178
rect 23718 6118 23858 6178
rect 24722 6118 24862 6178
rect 25726 6118 25866 6178
rect 26730 6118 26870 6178
rect 27734 6118 27874 6178
rect 28738 6118 28878 6178
rect 29742 6118 29882 6178
rect 30746 6118 30886 6178
rect 31750 6118 31890 6178
rect 32754 6118 32894 6178
rect 33758 6118 33898 6178
rect 34762 6118 34796 6178
rect 1046 6035 1067 6106
rect 1138 6035 1162 6106
rect 1233 6035 1271 6106
rect 1342 6035 1366 6106
rect 1437 6035 1460 6106
rect 1046 5102 1460 6035
rect 36064 6106 36478 6294
rect 36064 6035 36085 6106
rect 36156 6035 36180 6106
rect 36251 6035 36289 6106
rect 36360 6035 36384 6106
rect 36455 6035 36478 6106
rect 2888 5864 2948 6004
rect 3464 5864 3524 6004
rect 3892 5864 3952 6004
rect 4468 5864 4528 6004
rect 4896 5864 4956 6004
rect 5472 5864 5532 6004
rect 5900 5864 5960 6004
rect 6476 5864 6536 6004
rect 6904 5864 6964 6004
rect 7480 5864 7540 6004
rect 7908 5864 7968 6004
rect 8484 5864 8544 6004
rect 8912 5864 8972 6004
rect 9488 5864 9548 6004
rect 9916 5864 9976 6004
rect 10492 5864 10552 6004
rect 10920 5864 10980 6004
rect 11496 5864 11556 6004
rect 11924 5864 11984 6004
rect 12500 5864 12560 6004
rect 12928 5864 12988 6004
rect 13504 5864 13564 6004
rect 13932 5864 13992 6004
rect 14508 5864 14568 6004
rect 14936 5864 14996 6004
rect 15512 5864 15572 6004
rect 15940 5864 16000 6004
rect 16516 5864 16576 6004
rect 16944 5864 17004 6004
rect 17520 5864 17580 6004
rect 17948 5864 18008 6004
rect 18524 5864 18584 6004
rect 18952 5864 19012 6004
rect 19528 5864 19588 6004
rect 19956 5864 20016 6004
rect 20532 5864 20592 6004
rect 20960 5864 21020 6004
rect 21536 5864 21596 6004
rect 21964 5864 22024 6004
rect 22540 5864 22600 6004
rect 22968 5864 23028 6004
rect 23544 5864 23604 6004
rect 23972 5864 24032 6004
rect 24548 5864 24608 6004
rect 24976 5864 25036 6004
rect 25552 5864 25612 6004
rect 25980 5864 26040 6004
rect 26556 5864 26616 6004
rect 26984 5864 27044 6004
rect 27560 5864 27620 6004
rect 27988 5864 28048 6004
rect 28564 5864 28624 6004
rect 28992 5864 29052 6004
rect 29568 5864 29628 6004
rect 29996 5864 30056 6004
rect 30572 5864 30632 6004
rect 31000 5864 31060 6004
rect 31576 5864 31636 6004
rect 32004 5864 32064 6004
rect 32580 5864 32640 6004
rect 33008 5864 33068 6004
rect 33584 5864 33644 6004
rect 34012 5864 34072 6004
rect 34588 5864 34648 6004
rect 2736 5690 2774 5750
rect 3638 5690 3778 5750
rect 4642 5690 4782 5750
rect 5646 5690 5786 5750
rect 6650 5690 6790 5750
rect 7654 5690 7794 5750
rect 8658 5690 8798 5750
rect 9662 5690 9802 5750
rect 10666 5690 10806 5750
rect 11670 5690 11810 5750
rect 12674 5690 12814 5750
rect 13678 5690 13818 5750
rect 14682 5690 14822 5750
rect 15686 5690 15826 5750
rect 16690 5690 16830 5750
rect 17694 5690 17834 5750
rect 18698 5690 18838 5750
rect 19702 5690 19842 5750
rect 20706 5690 20846 5750
rect 21710 5690 21850 5750
rect 22714 5690 22854 5750
rect 23718 5690 23858 5750
rect 24722 5690 24862 5750
rect 25726 5690 25866 5750
rect 26730 5690 26870 5750
rect 27734 5690 27874 5750
rect 28738 5690 28878 5750
rect 29742 5690 29882 5750
rect 30746 5690 30886 5750
rect 31750 5690 31890 5750
rect 32754 5690 32894 5750
rect 33758 5690 33898 5750
rect 34762 5690 34796 5750
rect 2736 5114 2774 5174
rect 3638 5114 3778 5174
rect 4642 5114 4782 5174
rect 5646 5114 5786 5174
rect 6650 5114 6790 5174
rect 7654 5114 7794 5174
rect 8658 5114 8798 5174
rect 9662 5114 9802 5174
rect 10666 5114 10806 5174
rect 11670 5114 11810 5174
rect 12674 5114 12814 5174
rect 13678 5114 13818 5174
rect 14682 5114 14822 5174
rect 15686 5114 15826 5174
rect 16690 5114 16830 5174
rect 17694 5114 17834 5174
rect 18698 5114 18838 5174
rect 19702 5114 19842 5174
rect 20706 5114 20846 5174
rect 21710 5114 21850 5174
rect 22714 5114 22854 5174
rect 23718 5114 23858 5174
rect 24722 5114 24862 5174
rect 25726 5114 25866 5174
rect 26730 5114 26870 5174
rect 27734 5114 27874 5174
rect 28738 5114 28878 5174
rect 29742 5114 29882 5174
rect 30746 5114 30886 5174
rect 31750 5114 31890 5174
rect 32754 5114 32894 5174
rect 33758 5114 33898 5174
rect 34762 5114 34796 5174
rect 1046 5031 1067 5102
rect 1138 5031 1162 5102
rect 1233 5031 1271 5102
rect 1342 5031 1366 5102
rect 1437 5031 1460 5102
rect 1046 4098 1460 5031
rect 36064 5102 36478 6035
rect 36064 5031 36085 5102
rect 36156 5031 36180 5102
rect 36251 5031 36289 5102
rect 36360 5031 36384 5102
rect 36455 5031 36478 5102
rect 2888 4860 2948 5000
rect 3464 4860 3524 5000
rect 3892 4860 3952 5000
rect 4468 4860 4528 5000
rect 4896 4860 4956 5000
rect 5472 4860 5532 5000
rect 5900 4860 5960 5000
rect 6476 4860 6536 5000
rect 6904 4860 6964 5000
rect 7480 4860 7540 5000
rect 7908 4860 7968 5000
rect 8484 4860 8544 5000
rect 8912 4860 8972 5000
rect 9488 4860 9548 5000
rect 9916 4860 9976 5000
rect 10492 4860 10552 5000
rect 10920 4860 10980 5000
rect 11496 4860 11556 5000
rect 11924 4860 11984 5000
rect 12500 4860 12560 5000
rect 12928 4860 12988 5000
rect 13504 4860 13564 5000
rect 13932 4860 13992 5000
rect 14508 4860 14568 5000
rect 14936 4860 14996 5000
rect 15512 4860 15572 5000
rect 15940 4860 16000 5000
rect 16516 4860 16576 5000
rect 16944 4860 17004 5000
rect 17520 4860 17580 5000
rect 17948 4860 18008 5000
rect 18524 4860 18584 5000
rect 18952 4860 19012 5000
rect 19528 4860 19588 5000
rect 19956 4860 20016 5000
rect 20532 4860 20592 5000
rect 20960 4860 21020 5000
rect 21536 4860 21596 5000
rect 21964 4860 22024 5000
rect 22540 4860 22600 5000
rect 22968 4860 23028 5000
rect 23544 4860 23604 5000
rect 23972 4860 24032 5000
rect 24548 4860 24608 5000
rect 24976 4860 25036 5000
rect 25552 4860 25612 5000
rect 25980 4860 26040 5000
rect 26556 4860 26616 5000
rect 26984 4860 27044 5000
rect 27560 4860 27620 5000
rect 27988 4860 28048 5000
rect 28564 4860 28624 5000
rect 28992 4860 29052 5000
rect 29568 4860 29628 5000
rect 29996 4860 30056 5000
rect 30572 4860 30632 5000
rect 31000 4860 31060 5000
rect 31576 4860 31636 5000
rect 32004 4860 32064 5000
rect 32580 4860 32640 5000
rect 33008 4860 33068 5000
rect 33584 4860 33644 5000
rect 34012 4860 34072 5000
rect 34588 4860 34648 5000
rect 2736 4686 2774 4746
rect 3638 4686 3778 4746
rect 4642 4686 4782 4746
rect 5646 4686 5786 4746
rect 6650 4686 6790 4746
rect 7654 4686 7794 4746
rect 8658 4686 8798 4746
rect 9662 4686 9802 4746
rect 10666 4686 10806 4746
rect 11670 4686 11810 4746
rect 12674 4686 12814 4746
rect 13678 4686 13818 4746
rect 14682 4686 14822 4746
rect 15686 4686 15826 4746
rect 16690 4686 16830 4746
rect 17694 4686 17834 4746
rect 18698 4686 18838 4746
rect 19702 4686 19842 4746
rect 20706 4686 20846 4746
rect 21710 4686 21850 4746
rect 22714 4686 22854 4746
rect 23718 4686 23858 4746
rect 24722 4686 24862 4746
rect 25726 4686 25866 4746
rect 26730 4686 26870 4746
rect 27734 4686 27874 4746
rect 28738 4686 28878 4746
rect 29742 4686 29882 4746
rect 30746 4686 30886 4746
rect 31750 4686 31890 4746
rect 32754 4686 32894 4746
rect 33758 4686 33898 4746
rect 34762 4686 34796 4746
rect 2736 4110 2774 4170
rect 3638 4110 3778 4170
rect 4642 4110 4782 4170
rect 5646 4110 5786 4170
rect 6650 4110 6790 4170
rect 7654 4110 7794 4170
rect 8658 4110 8798 4170
rect 9662 4110 9802 4170
rect 10666 4110 10806 4170
rect 11670 4110 11810 4170
rect 12674 4110 12814 4170
rect 13678 4110 13818 4170
rect 14682 4110 14822 4170
rect 15686 4110 15826 4170
rect 16690 4110 16830 4170
rect 17694 4110 17834 4170
rect 18698 4110 18838 4170
rect 19702 4110 19842 4170
rect 20706 4110 20846 4170
rect 21710 4110 21850 4170
rect 22714 4110 22854 4170
rect 23718 4110 23858 4170
rect 24722 4110 24862 4170
rect 25726 4110 25866 4170
rect 26730 4110 26870 4170
rect 27734 4110 27874 4170
rect 28738 4110 28878 4170
rect 29742 4110 29882 4170
rect 30746 4110 30886 4170
rect 31750 4110 31890 4170
rect 32754 4110 32894 4170
rect 33758 4110 33898 4170
rect 34762 4110 34796 4170
rect 1046 4027 1067 4098
rect 1138 4027 1162 4098
rect 1233 4027 1271 4098
rect 1342 4027 1366 4098
rect 1437 4027 1460 4098
rect 1046 3092 1460 4027
rect 36064 4098 36478 5031
rect 36064 4027 36085 4098
rect 36156 4027 36180 4098
rect 36251 4027 36289 4098
rect 36360 4027 36384 4098
rect 36455 4027 36478 4098
rect 2888 3856 2948 3996
rect 3464 3856 3524 3996
rect 3892 3856 3952 3996
rect 4468 3856 4528 3996
rect 4896 3856 4956 3996
rect 5472 3856 5532 3996
rect 5900 3856 5960 3996
rect 6476 3856 6536 3996
rect 6904 3856 6964 3996
rect 7480 3856 7540 3996
rect 7908 3856 7968 3996
rect 8484 3856 8544 3996
rect 8912 3856 8972 3996
rect 9488 3856 9548 3996
rect 9916 3856 9976 3996
rect 10492 3856 10552 3996
rect 10920 3856 10980 3996
rect 11496 3856 11556 3996
rect 11924 3856 11984 3996
rect 12500 3856 12560 3996
rect 12928 3856 12988 3996
rect 13504 3856 13564 3996
rect 13932 3856 13992 3996
rect 14508 3856 14568 3996
rect 14936 3856 14996 3996
rect 15512 3856 15572 3996
rect 15940 3856 16000 3996
rect 16516 3856 16576 3996
rect 16944 3856 17004 3996
rect 17520 3856 17580 3996
rect 17948 3856 18008 3996
rect 18524 3856 18584 3996
rect 18952 3856 19012 3996
rect 19528 3856 19588 3996
rect 19956 3856 20016 3996
rect 20532 3856 20592 3996
rect 20960 3856 21020 3996
rect 21536 3856 21596 3996
rect 21964 3856 22024 3996
rect 22540 3856 22600 3996
rect 22968 3856 23028 3996
rect 23544 3856 23604 3996
rect 23972 3856 24032 3996
rect 24548 3856 24608 3996
rect 24976 3856 25036 3996
rect 25552 3856 25612 3996
rect 25980 3856 26040 3996
rect 26556 3856 26616 3996
rect 26984 3856 27044 3996
rect 27560 3856 27620 3996
rect 27988 3856 28048 3996
rect 28564 3856 28624 3996
rect 28992 3856 29052 3996
rect 29568 3856 29628 3996
rect 29996 3856 30056 3996
rect 30572 3856 30632 3996
rect 31000 3856 31060 3996
rect 31576 3856 31636 3996
rect 32004 3856 32064 3996
rect 32580 3856 32640 3996
rect 33008 3856 33068 3996
rect 33584 3856 33644 3996
rect 34012 3856 34072 3996
rect 34588 3856 34648 3996
rect 2736 3682 2774 3742
rect 3638 3682 3778 3742
rect 4642 3682 4782 3742
rect 5646 3682 5786 3742
rect 6650 3682 6790 3742
rect 7654 3682 7794 3742
rect 8658 3682 8798 3742
rect 9662 3682 9802 3742
rect 10666 3682 10806 3742
rect 11670 3682 11810 3742
rect 12674 3682 12814 3742
rect 13678 3682 13818 3742
rect 14682 3682 14822 3742
rect 15686 3682 15826 3742
rect 16690 3682 16830 3742
rect 17694 3682 17834 3742
rect 18698 3682 18838 3742
rect 19702 3682 19842 3742
rect 20706 3682 20846 3742
rect 21710 3682 21850 3742
rect 22714 3682 22854 3742
rect 23718 3682 23858 3742
rect 24722 3682 24862 3742
rect 25726 3682 25866 3742
rect 26730 3682 26870 3742
rect 27734 3682 27874 3742
rect 28738 3682 28878 3742
rect 29742 3682 29882 3742
rect 30746 3682 30886 3742
rect 31750 3682 31890 3742
rect 32754 3682 32894 3742
rect 33758 3682 33898 3742
rect 34762 3682 34796 3742
rect 36064 3589 36478 4027
rect 36064 3525 36094 3589
rect 36158 3525 36190 3589
rect 36254 3525 36286 3589
rect 36350 3525 36382 3589
rect 36446 3525 36478 3589
rect 36064 3498 36478 3525
rect 36064 3434 36094 3498
rect 36158 3434 36190 3498
rect 36254 3434 36286 3498
rect 36350 3434 36382 3498
rect 36446 3434 36478 3498
rect 36064 3407 36478 3434
rect 36064 3343 36094 3407
rect 36158 3343 36190 3407
rect 36254 3343 36286 3407
rect 36350 3343 36382 3407
rect 36446 3343 36478 3407
rect 2736 3106 2774 3166
rect 3638 3106 3778 3166
rect 4642 3106 4782 3166
rect 5646 3106 5786 3166
rect 6650 3106 6790 3166
rect 7654 3106 7794 3166
rect 8658 3106 8798 3166
rect 9662 3106 9802 3166
rect 10666 3106 10806 3166
rect 11670 3106 11810 3166
rect 12674 3106 12814 3166
rect 13678 3106 13818 3166
rect 14682 3106 14822 3166
rect 15686 3106 15826 3166
rect 16690 3106 16830 3166
rect 17694 3106 17834 3166
rect 18698 3106 18838 3166
rect 19702 3106 19842 3166
rect 20706 3106 20846 3166
rect 21710 3106 21850 3166
rect 22714 3106 22854 3166
rect 23718 3106 23858 3166
rect 24722 3106 24862 3166
rect 25726 3106 25866 3166
rect 26730 3106 26870 3166
rect 27734 3106 27874 3166
rect 28738 3106 28878 3166
rect 29742 3106 29882 3166
rect 30746 3106 30886 3166
rect 31750 3106 31890 3166
rect 32754 3106 32894 3166
rect 33758 3106 33898 3166
rect 34762 3106 34796 3166
rect 1046 3021 1067 3092
rect 1138 3021 1162 3092
rect 1233 3021 1271 3092
rect 1342 3021 1366 3092
rect 1437 3021 1460 3092
rect 1046 2089 1460 3021
rect 36064 3094 36478 3343
rect 36064 3023 36085 3094
rect 36156 3023 36180 3094
rect 36251 3023 36289 3094
rect 36360 3023 36384 3094
rect 36455 3023 36478 3094
rect 2888 2958 2948 2992
rect 3464 2958 3524 2992
rect 3892 2852 3952 2992
rect 4468 2852 4528 2992
rect 4896 2852 4956 2992
rect 5472 2852 5532 2992
rect 5900 2852 5960 2992
rect 6476 2852 6536 2992
rect 6904 2852 6964 2992
rect 7480 2852 7540 2992
rect 7908 2852 7968 2992
rect 8484 2852 8544 2992
rect 8912 2852 8972 2992
rect 9488 2852 9548 2992
rect 9916 2852 9976 2992
rect 10492 2852 10552 2992
rect 10920 2852 10980 2992
rect 11496 2852 11556 2992
rect 11924 2852 11984 2992
rect 12500 2852 12560 2992
rect 12928 2852 12988 2992
rect 13504 2852 13564 2992
rect 13932 2852 13992 2992
rect 14508 2852 14568 2992
rect 14936 2852 14996 2992
rect 15512 2852 15572 2992
rect 15940 2852 16000 2992
rect 16516 2852 16576 2992
rect 16944 2852 17004 2992
rect 17520 2852 17580 2992
rect 17948 2852 18008 2992
rect 18524 2852 18584 2992
rect 18952 2852 19012 2992
rect 19528 2852 19588 2992
rect 19956 2852 20016 2992
rect 20532 2852 20592 2992
rect 20960 2852 21020 2992
rect 21536 2852 21596 2992
rect 21964 2852 22024 2992
rect 22540 2852 22600 2992
rect 22968 2852 23028 2992
rect 23544 2852 23604 2992
rect 23972 2852 24032 2992
rect 24548 2852 24608 2992
rect 24976 2852 25036 2992
rect 25552 2852 25612 2992
rect 25980 2852 26040 2992
rect 26556 2852 26616 2992
rect 26984 2852 27044 2992
rect 27560 2852 27620 2992
rect 27988 2852 28048 2992
rect 28564 2852 28624 2992
rect 28992 2852 29052 2992
rect 29568 2852 29628 2992
rect 29996 2852 30056 2992
rect 30572 2852 30632 2992
rect 31000 2852 31060 2992
rect 31576 2852 31636 2992
rect 32004 2852 32064 2992
rect 32580 2852 32640 2992
rect 33008 2852 33068 2992
rect 33584 2852 33644 2992
rect 34012 2852 34072 2992
rect 34588 2852 34648 2992
rect 3744 2678 3778 2738
rect 4642 2678 4782 2738
rect 5646 2678 5786 2738
rect 6650 2678 6790 2738
rect 7654 2678 7794 2738
rect 8658 2678 8798 2738
rect 9662 2678 9802 2738
rect 10666 2678 10806 2738
rect 11670 2678 11810 2738
rect 12674 2678 12814 2738
rect 13678 2678 13818 2738
rect 14682 2678 14822 2738
rect 15686 2678 15826 2738
rect 16690 2678 16830 2738
rect 17694 2678 17834 2738
rect 18698 2678 18838 2738
rect 19702 2678 19842 2738
rect 20706 2678 20846 2738
rect 21710 2678 21850 2738
rect 22714 2678 22854 2738
rect 23718 2678 23858 2738
rect 24722 2678 24862 2738
rect 25726 2678 25866 2738
rect 26730 2678 26870 2738
rect 27734 2678 27874 2738
rect 28738 2678 28878 2738
rect 29742 2678 29882 2738
rect 30746 2678 30886 2738
rect 31750 2678 31890 2738
rect 32754 2678 32894 2738
rect 33758 2678 33898 2738
rect 34762 2678 34796 2738
rect 3744 2102 3778 2162
rect 4642 2102 4782 2162
rect 5646 2102 5786 2162
rect 6650 2102 6790 2162
rect 7654 2102 7794 2162
rect 8658 2102 8798 2162
rect 9662 2102 9802 2162
rect 10666 2102 10806 2162
rect 11670 2102 11810 2162
rect 12674 2102 12814 2162
rect 13678 2102 13818 2162
rect 14682 2102 14822 2162
rect 15686 2102 15826 2162
rect 16690 2102 16830 2162
rect 17694 2102 17834 2162
rect 18698 2102 18838 2162
rect 19702 2102 19842 2162
rect 20706 2102 20846 2162
rect 21710 2102 21850 2162
rect 22714 2102 22854 2162
rect 23718 2102 23858 2162
rect 24722 2102 24862 2162
rect 25726 2102 25866 2162
rect 26730 2102 26870 2162
rect 27734 2102 27874 2162
rect 28738 2102 28878 2162
rect 29742 2102 29882 2162
rect 30746 2102 30886 2162
rect 31750 2102 31890 2162
rect 32754 2102 32894 2162
rect 33758 2102 33898 2162
rect 34762 2102 34796 2162
rect 1046 2018 1067 2089
rect 1138 2018 1162 2089
rect 1233 2018 1271 2089
rect 1342 2018 1366 2089
rect 1437 2018 1460 2089
rect 1046 1434 1460 2018
rect 36064 2090 36478 3023
rect 36064 2019 36085 2090
rect 36156 2019 36180 2090
rect 36251 2019 36289 2090
rect 36360 2019 36384 2090
rect 36455 2019 36478 2090
rect 3892 1848 3952 1988
rect 4468 1950 4528 1988
rect 4896 1950 4956 1988
rect 5472 1950 5532 1988
rect 5900 1950 5960 1988
rect 6476 1950 6536 1988
rect 6904 1950 6964 1988
rect 7480 1950 7540 1988
rect 7908 1950 7968 1988
rect 8484 1950 8544 1988
rect 8912 1950 8972 1988
rect 9488 1950 9548 1988
rect 9916 1950 9976 1988
rect 10492 1950 10552 1988
rect 10920 1950 10980 1988
rect 11496 1950 11556 1988
rect 11924 1950 11984 1988
rect 12500 1950 12560 1988
rect 12928 1950 12988 1988
rect 13504 1950 13564 1988
rect 13932 1950 13992 1988
rect 14508 1950 14568 1988
rect 14936 1950 14996 1988
rect 15512 1950 15572 1988
rect 15940 1950 16000 1988
rect 16516 1950 16576 1988
rect 16944 1950 17004 1988
rect 17520 1950 17580 1988
rect 17948 1950 18008 1988
rect 18524 1848 18584 1988
rect 18952 1848 19012 1988
rect 19528 1848 19588 1988
rect 19956 1950 20016 1988
rect 20532 1950 20592 1988
rect 20960 1950 21020 1988
rect 21536 1950 21596 1988
rect 21964 1950 22024 1988
rect 22540 1950 22600 1988
rect 22968 1950 23028 1988
rect 23544 1950 23604 1988
rect 23972 1950 24032 1988
rect 24548 1950 24608 1988
rect 24976 1950 25036 1988
rect 25552 1950 25612 1988
rect 25980 1950 26040 1988
rect 26556 1950 26616 1988
rect 26984 1950 27044 1988
rect 27560 1950 27620 1988
rect 27988 1950 28048 1988
rect 28564 1950 28624 1988
rect 28992 1950 29052 1988
rect 29568 1950 29628 1988
rect 29996 1950 30056 1988
rect 30572 1950 30632 1988
rect 31000 1950 31060 1988
rect 31576 1950 31636 1988
rect 32004 1950 32064 1988
rect 32580 1950 32640 1988
rect 33008 1950 33068 1988
rect 33584 1950 33644 1988
rect 34012 1950 34072 1988
rect 34300 1848 34360 1988
rect 34588 1950 34648 1988
rect 18698 1674 18838 1734
rect 19702 1674 19842 1734
rect 1046 1363 1067 1434
rect 1138 1363 1162 1434
rect 1233 1363 1271 1434
rect 1342 1363 1366 1434
rect 1437 1363 1460 1434
rect 1046 1324 1460 1363
rect 1046 1253 1067 1324
rect 1138 1253 1162 1324
rect 1233 1253 1271 1324
rect 1342 1253 1366 1324
rect 1437 1253 1460 1324
rect 1046 1085 1460 1253
rect 1046 1014 1067 1085
rect 1138 1014 1162 1085
rect 1233 1014 1271 1085
rect 1342 1014 1366 1085
rect 1437 1014 1460 1085
rect 1046 42 1460 1014
rect 36064 1086 36478 2019
rect 36064 1015 36085 1086
rect 36156 1015 36180 1086
rect 36251 1015 36289 1086
rect 36360 1015 36384 1086
rect 36455 1015 36478 1086
rect 34300 0 34360 962
rect 36064 881 36478 1015
rect 36064 817 36094 881
rect 36158 817 36190 881
rect 36254 817 36286 881
rect 36350 817 36382 881
rect 36446 817 36478 881
rect 36064 790 36478 817
rect 36064 726 36094 790
rect 36158 726 36190 790
rect 36254 726 36286 790
rect 36350 726 36382 790
rect 36446 726 36478 790
rect 36064 699 36478 726
rect 36064 635 36094 699
rect 36158 635 36190 699
rect 36254 635 36286 699
rect 36350 635 36382 699
rect 36446 635 36478 699
rect 36064 172 36478 635
rect 36540 6241 37431 6305
rect 37495 6241 37602 6305
rect 41908 6264 42322 6624
rect 36540 6193 37602 6241
rect 36540 6129 37430 6193
rect 37494 6129 37602 6193
rect 36540 6075 37602 6129
rect 41602 6246 42322 6264
rect 41602 6096 41930 6246
rect 42142 6096 42322 6246
rect 41602 6082 42322 6096
rect 36540 6011 37430 6075
rect 37494 6011 37602 6075
rect 36540 5986 37602 6011
rect 36540 5818 36954 5986
rect 36540 5747 36561 5818
rect 36632 5747 36656 5818
rect 36727 5747 36765 5818
rect 36836 5747 36860 5818
rect 36931 5747 36954 5818
rect 36540 4814 36954 5747
rect 41908 5708 42322 6082
rect 41602 5690 42322 5708
rect 41602 5540 41930 5690
rect 42142 5540 42322 5690
rect 41602 5526 42322 5540
rect 36540 4743 36561 4814
rect 36632 4743 36656 4814
rect 36727 4743 36765 4814
rect 36836 4743 36860 4814
rect 36931 4743 36954 4814
rect 36540 3810 36954 4743
rect 41602 4545 41847 4558
rect 41602 4388 41707 4545
rect 41821 4388 41847 4545
rect 41602 4374 41847 4388
rect 36540 3739 36561 3810
rect 36632 3739 36656 3810
rect 36727 3739 36765 3810
rect 36836 3739 36860 3810
rect 36931 3739 36954 3810
rect 36540 2806 36954 3739
rect 41602 3655 41847 3668
rect 37394 3587 37602 3617
rect 37394 3523 37423 3587
rect 37487 3523 37602 3587
rect 37394 3495 37602 3523
rect 37394 3431 37423 3495
rect 37487 3431 37602 3495
rect 41602 3498 41707 3655
rect 41821 3498 41847 3655
rect 41602 3484 41847 3498
rect 37394 3404 37602 3431
rect 37394 3340 37423 3404
rect 37487 3340 37602 3404
rect 37394 3318 37602 3340
rect 41908 2806 42322 5526
rect 36540 2735 36561 2806
rect 36632 2735 36656 2806
rect 36727 2735 36765 2806
rect 36836 2735 36860 2806
rect 36931 2735 36954 2806
rect 36540 2336 36954 2735
rect 41602 2788 42322 2806
rect 41602 2638 41930 2788
rect 42142 2638 42322 2788
rect 41602 2624 42322 2638
rect 36540 2311 37602 2336
rect 36540 2247 37431 2311
rect 37495 2247 37602 2311
rect 41908 2264 42322 2624
rect 36540 2199 37602 2247
rect 36540 2135 37430 2199
rect 37494 2135 37602 2199
rect 36540 2081 37602 2135
rect 41602 2246 42322 2264
rect 41602 2096 41930 2246
rect 42142 2096 42322 2246
rect 41602 2082 42322 2096
rect 36540 2017 37430 2081
rect 37494 2017 37602 2081
rect 36540 1992 37602 2017
rect 36540 1802 36954 1992
rect 36540 1731 36561 1802
rect 36632 1731 36656 1802
rect 36727 1731 36765 1802
rect 36836 1731 36860 1802
rect 36931 1731 36954 1802
rect 36540 526 36954 1731
rect 41908 1708 42322 2082
rect 41602 1690 42322 1708
rect 41602 1540 41930 1690
rect 42142 1540 42322 1690
rect 41602 1526 42322 1540
rect 37394 879 37602 909
rect 37394 815 37423 879
rect 37487 815 37602 879
rect 37394 787 37602 815
rect 37394 723 37423 787
rect 37487 723 37602 787
rect 37394 696 37602 723
rect 37394 632 37423 696
rect 37487 632 37602 696
rect 37394 610 37602 632
rect 36540 455 36561 526
rect 36632 455 36656 526
rect 36727 455 36765 526
rect 36836 455 36860 526
rect 36931 455 36954 526
rect 36540 172 36954 455
rect 41602 544 41847 557
rect 41602 387 41707 544
rect 41821 387 41847 544
rect 41602 373 41847 387
rect 41908 166 42322 1526
rect 42396 23656 42810 24168
rect 42396 23494 42410 23656
rect 42648 23494 42810 23656
rect 42396 23250 42810 23494
rect 42396 22838 42422 23250
rect 42634 22838 42810 23250
rect 42396 21492 42810 22838
rect 42396 21080 42422 21492
rect 42634 21080 42810 21492
rect 42396 20546 42810 21080
rect 42396 20384 42410 20546
rect 42648 20384 42810 20546
rect 42396 19656 42810 20384
rect 42396 19494 42410 19656
rect 42648 19494 42810 19656
rect 42396 19250 42810 19494
rect 42396 18838 42422 19250
rect 42634 18838 42810 19250
rect 42396 17492 42810 18838
rect 42396 17080 42422 17492
rect 42634 17080 42810 17492
rect 42396 16546 42810 17080
rect 42396 16384 42410 16546
rect 42648 16384 42810 16546
rect 42396 15656 42810 16384
rect 42396 15494 42410 15656
rect 42648 15494 42810 15656
rect 42396 15250 42810 15494
rect 42396 14838 42422 15250
rect 42634 14838 42810 15250
rect 42396 13492 42810 14838
rect 42396 13080 42422 13492
rect 42634 13080 42810 13492
rect 42396 12546 42810 13080
rect 42396 12384 42410 12546
rect 42648 12384 42810 12546
rect 42396 11656 42810 12384
rect 42396 11494 42410 11656
rect 42648 11494 42810 11656
rect 42396 11250 42810 11494
rect 42396 10838 42422 11250
rect 42634 10838 42810 11250
rect 42396 9492 42810 10838
rect 42396 9080 42422 9492
rect 42634 9080 42810 9492
rect 42396 8546 42810 9080
rect 42396 8384 42410 8546
rect 42648 8384 42810 8546
rect 42396 7656 42810 8384
rect 42396 7494 42410 7656
rect 42648 7494 42810 7656
rect 42396 7250 42810 7494
rect 42396 6838 42422 7250
rect 42634 6838 42810 7250
rect 42396 5492 42810 6838
rect 42396 5080 42422 5492
rect 42634 5080 42810 5492
rect 42396 4546 42810 5080
rect 42396 4384 42410 4546
rect 42648 4384 42810 4546
rect 42396 3656 42810 4384
rect 42396 3494 42410 3656
rect 42648 3494 42810 3656
rect 42396 3250 42810 3494
rect 42396 2838 42422 3250
rect 42634 2838 42810 3250
rect 42396 1492 42810 2838
rect 42396 1080 42422 1492
rect 42634 1080 42810 1492
rect 42396 546 42810 1080
rect 42396 384 42410 546
rect 42648 384 42810 546
rect 42396 168 42810 384
use adc_array_wafflecap_1  adc_array_wafflecap_1_0
timestamp 1664894364
transform 1 0 19772 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_1  adc_array_wafflecap_1_1
timestamp 1664894364
transform 1 0 3708 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_2  adc_array_wafflecap_2_0
timestamp 1665042887
transform 1 0 17764 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_4  adc_array_wafflecap_4_0
timestamp 1664894853
transform 1 0 18768 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_8  adc_array_wafflecap_8_0
array 0 31 1004 0 14 1004
timestamp 1664895084
transform 1 0 2704 0 1 2922
box 0 0 1004 1004
use adc_array_wafflecap_8  adc_array_wafflecap_8_1
array 0 30 1004 0 0 1004
timestamp 1664895084
transform 1 0 3708 0 1 1918
box 0 0 1004 1004
use adc_array_wafflecap_drv  adc_array_wafflecap_drv_0
array 0 0 1004 0 15 1004
timestamp 1664895328
transform 1 0 1700 0 1 1918
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_0
array 0 1 1004 0 0 1004
timestamp 1664895551
transform 1 0 1700 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_1
array 0 12 1004 0 0 1004
timestamp 1664895551
transform 1 0 4712 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_3
array 0 12 1004 0 0 1004
timestamp 1664895551
transform 1 0 20776 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_4
array 0 33 1004 0 0 1004
timestamp 1664895551
transform 1 0 1700 0 1 17982
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_5
array 0 0 1004 0 15 1004
timestamp 1664895551
transform 1 0 34832 0 1 1918
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_6
timestamp 1664895551
transform 1 0 34832 0 1 914
box 0 0 1004 1004
use adc_array_wafflecap_dummy  adc_array_wafflecap_dummy_7
timestamp 1664895551
transform 1 0 2704 0 1 1918
box 0 0 1004 1004
use adc_array_wafflecap_gate  adc_array_wafflecap_gate_0
timestamp 1665691632
transform 1 0 33828 0 1 914
box 0 0 1004 1004
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0
array 0 0 4000 0 5 4000
timestamp 1663849571
transform 1 0 37602 0 1 166
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 8 4000 0 0 4000
timestamp 1663849571
transform 1 0 1602 0 1 20166
box 0 0 4000 4000
<< labels >>
flabel metal4 s 42396 168 42810 24168 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 s 41908 166 42322 24166 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal2 398 0 534 18986 0 FreeSans 1600 90 0 0 vcm
port 3 nsew signal input
rlabel metal2 290 0 358 76 5 sample
port 4 s signal input
rlabel metal2 182 0 250 76 5 sample_n
port 5 s signal input
flabel metal4 s 36540 172 36954 19902 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 36064 172 36478 19902 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 s 570 42 984 24166 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 1046 42 1460 24166 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal2 s 18286 0 18320 42 5 FreeSans 160 0 0 0 en_bit_n[1]
port 71 s signal input
flabel metal2 s 19290 0 19324 42 5 FreeSans 160 0 0 0 en_bit_n[2]
port 70 s signal input
flabel metal2 s 20294 0 20328 42 5 FreeSans 160 0 0 0 en_bit_n[0]
port 72 s signal input
flabel metal2 s 4230 0 4264 42 5 FreeSans 160 0 0 0 en_C0_n
port 73 s signal input
flabel metal2 s 26650 0 26684 42 5 FreeSans 160 0 0 0 col_n[23]
port 46 s signal input
flabel metal2 s 25646 0 25680 42 5 FreeSans 160 0 0 0 col_n[22]
port 47 s signal input
flabel metal2 s 24642 0 24676 42 5 FreeSans 160 0 0 0 col_n[21]
port 48 s signal input
flabel metal2 s 23638 0 23672 42 5 FreeSans 160 0 0 0 col_n[20]
port 49 s signal input
flabel metal2 s 22634 0 22668 42 5 FreeSans 160 0 0 0 col_n[19]
port 50 s signal input
flabel metal2 s 21630 0 21664 42 5 FreeSans 160 0 0 0 col_n[18]
port 51 s signal input
flabel metal2 s 20626 0 20660 42 5 FreeSans 160 0 0 0 col_n[17]
port 52 s signal input
flabel metal2 s 19622 0 19656 42 5 FreeSans 160 0 0 0 col_n[16]
port 53 s signal input
flabel metal2 s 18618 0 18652 42 5 FreeSans 160 0 0 0 col_n[15]
port 54 s signal input
flabel metal2 s 17614 0 17648 42 5 FreeSans 160 0 0 0 col_n[14]
port 55 s signal input
flabel metal2 s 16610 0 16644 42 5 FreeSans 160 0 0 0 col_n[13]
port 56 s signal input
flabel metal2 s 15606 0 15640 42 5 FreeSans 160 0 0 0 col_n[12]
port 57 s signal input
flabel metal2 s 14602 0 14636 42 5 FreeSans 160 0 0 0 col_n[11]
port 58 s signal input
flabel metal2 s 13598 0 13632 42 5 FreeSans 160 0 0 0 col_n[10]
port 59 s signal input
flabel metal2 s 12594 0 12628 42 5 FreeSans 160 0 0 0 col_n[9]
port 60 s signal input
flabel metal2 s 11590 0 11624 42 5 FreeSans 160 0 0 0 col_n[8]
port 61 s signal input
flabel metal2 s 10586 0 10620 42 5 FreeSans 160 0 0 0 col_n[7]
port 62 s signal input
flabel metal2 s 9582 0 9616 42 5 FreeSans 160 0 0 0 col_n[6]
port 63 s signal input
flabel metal2 s 8578 0 8612 42 5 FreeSans 160 0 0 0 col_n[5]
port 64 s signal input
flabel metal2 s 7574 0 7608 42 5 FreeSans 160 0 0 0 col_n[4]
port 65 s signal input
flabel metal2 s 6570 0 6604 42 5 FreeSans 160 0 0 0 col_n[3]
port 66 s signal input
flabel metal2 s 5566 0 5600 42 5 FreeSans 160 0 0 0 col_n[2]
port 67 s signal input
flabel metal2 s 4562 0 4596 42 5 FreeSans 160 0 0 0 col_n[1]
port 68 s signal input
flabel metal2 s 3558 0 3592 42 5 FreeSans 160 0 0 0 col_n[0]
port 69 s signal input
flabel metal2 s 28470 0 28504 42 5 FreeSans 160 0 0 0 col_n[28]
port 41 s signal input
flabel metal2 s 28266 0 28300 42 5 FreeSans 160 0 0 0 col_n[27]
port 42 s signal input
flabel metal2 s 28062 0 28096 42 5 FreeSans 160 0 0 0 col_n[26]
port 43 s signal input
flabel metal2 s 27858 0 27892 42 5 FreeSans 160 0 0 0 col_n[25]
port 44 s signal input
flabel metal2 s 27654 0 27688 42 5 FreeSans 160 0 0 0 col_n[24]
port 45 s signal input
flabel metal2 s 29082 0 29116 42 5 FreeSans 160 0 0 0 col_n[31]
port 38 s signal input
flabel metal2 s 28878 0 28912 42 5 FreeSans 160 0 0 0 col_n[30]
port 39 s signal input
flabel metal2 s 28674 0 28708 42 5 FreeSans 160 0 0 0 col_n[29]
port 40 s signal input
flabel metal4 s 34300 0 34360 58 5 FreeSans 160 0 0 0 ctop
port 77 s signal output
flabel metal1 s 42622 8 42810 124 0 FreeSans 320 0 0 0 analog_in
port 76 nsew signal input
flabel metal1 s 0 17490 106 17518 7 FreeSans 160 0 0 0 rowon_n[15]
port 22 w signal input
flabel metal1 s 0 16486 106 16514 7 FreeSans 160 0 0 0 rowon_n[14]
port 23 w signal input
flabel metal1 s 0 15482 106 15510 7 FreeSans 160 0 0 0 rowon_n[13]
port 24 w signal input
flabel metal1 s 0 14478 106 14506 7 FreeSans 160 0 0 0 rowon_n[12]
port 25 w signal input
flabel metal1 s 0 13474 106 13502 7 FreeSans 160 0 0 0 rowon_n[11]
port 26 w signal input
flabel metal1 s 0 12470 106 12498 7 FreeSans 160 0 0 0 rowon_n[10]
port 27 w signal input
flabel metal1 s 0 11466 106 11494 7 FreeSans 160 0 0 0 rowon_n[9]
port 28 w signal input
flabel metal1 s 0 10462 106 10490 7 FreeSans 160 0 0 0 rowon_n[8]
port 29 w signal input
flabel metal1 s 0 9458 106 9486 7 FreeSans 160 0 0 0 rowon_n[7]
port 30 w signal input
flabel metal1 s 0 8454 106 8482 7 FreeSans 160 0 0 0 rowon_n[6]
port 31 w signal input
flabel metal1 s 0 7450 106 7478 7 FreeSans 160 0 0 0 rowon_n[5]
port 32 w signal input
flabel metal1 s 0 5442 106 5470 7 FreeSans 160 0 0 0 rowon_n[3]
port 34 w signal input
flabel metal1 s 0 4438 106 4466 7 FreeSans 160 0 0 0 rowon_n[2]
port 35 w signal input
flabel metal1 s 0 3434 106 3462 7 FreeSans 160 0 0 0 rowon_n[1]
port 36 w signal input
flabel metal1 s 0 2430 106 2458 7 FreeSans 160 0 0 0 rowon_n[0]
port 37 w signal input
flabel metal1 s 0 17408 106 17436 7 FreeSans 160 0 0 0 row_n[15]
port 6 w signal input
flabel metal1 s 0 16404 106 16432 7 FreeSans 160 0 0 0 row_n[14]
port 7 w signal input
flabel metal1 s 0 15400 106 15428 7 FreeSans 160 0 0 0 row_n[13]
port 8 w signal input
flabel metal1 s 0 14396 106 14424 7 FreeSans 160 0 0 0 row_n[12]
port 9 w signal input
flabel metal1 s 0 13392 106 13420 7 FreeSans 160 0 0 0 row_n[11]
port 10 w signal input
flabel metal1 s 0 12388 106 12416 7 FreeSans 160 0 0 0 row_n[10]
port 11 w signal input
flabel metal1 s 0 11384 106 11412 7 FreeSans 160 0 0 0 row_n[9]
port 12 w signal input
flabel metal1 s 0 10380 106 10408 7 FreeSans 160 0 0 0 row_n[8]
port 13 w signal input
flabel metal1 s 0 9376 106 9404 7 FreeSans 160 0 0 0 row_n[7]
port 14 w signal input
flabel metal1 s 0 8372 106 8400 7 FreeSans 160 0 0 0 row_n[6]
port 15 w signal input
flabel metal1 s 0 7368 106 7396 7 FreeSans 160 0 0 0 row_n[5]
port 16 w signal input
flabel metal1 s 0 6364 106 6392 7 FreeSans 160 0 0 0 row_n[4]
port 17 w signal input
flabel metal1 s 0 5360 106 5388 7 FreeSans 160 0 0 0 row_n[3]
port 18 w signal input
flabel metal1 s 0 4356 106 4384 7 FreeSans 160 0 0 0 row_n[2]
port 19 w signal input
flabel metal1 s 0 3352 106 3380 7 FreeSans 160 0 0 0 row_n[1]
port 20 w signal input
flabel metal1 s 0 2348 106 2376 7 FreeSans 160 0 0 0 row_n[0]
port 21 w signal input
flabel metal1 s 0 6446 106 6474 7 FreeSans 160 0 0 0 rowon_n[4]
port 33 w signal input
flabel metal2 s 34554 0 34593 42 5 FreeSans 160 90 0 0 sw_n
port 75 s signal input
flabel metal2 s 34180 0 34219 42 5 FreeSans 160 90 0 0 sw
port 74 s signal input
<< properties >>
string FIXED_BBOX 0 0 42810 24168
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
