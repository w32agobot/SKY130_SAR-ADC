magic
tech sky130A
magscale 1 2
timestamp 1673727735
<< nwell >>
rect 0 178 208 576
<< nmos >>
rect 62 22 146 52
<< pmos >>
rect 62 364 146 394
rect 62 272 146 302
<< ndiff >>
rect 62 98 146 110
rect 62 64 74 98
rect 134 64 146 98
rect 62 52 146 64
rect 62 10 146 22
rect 62 -24 74 10
rect 134 -24 146 10
rect 62 -36 146 -24
<< pdiff >>
rect 62 442 146 450
rect 62 408 74 442
rect 134 408 146 442
rect 62 394 146 408
rect 62 350 146 364
rect 62 316 74 350
rect 134 316 146 350
rect 62 302 146 316
rect 62 260 146 272
rect 62 226 74 260
rect 134 226 146 260
rect 62 214 146 226
<< ndiffc >>
rect 74 64 134 98
rect 74 -24 134 10
<< pdiffc >>
rect 74 408 134 442
rect 74 316 134 350
rect 74 226 134 260
<< psubdiff >>
rect 62 -124 86 -90
rect 122 -124 146 -90
rect 62 -130 146 -124
<< nsubdiff >>
rect 62 504 86 540
rect 122 504 146 540
<< psubdiffcont >>
rect 86 -124 122 -90
<< nsubdiffcont >>
rect 86 504 122 540
<< poly >>
rect -29 375 62 394
rect -29 296 -19 375
rect 15 364 62 375
rect 146 364 172 394
rect 15 302 46 364
rect 15 296 62 302
rect -29 272 62 296
rect 146 272 172 302
rect -26 55 40 65
rect -26 21 -10 55
rect 24 52 40 55
rect 24 22 62 52
rect 146 22 172 52
rect 24 21 40 22
rect -26 5 40 21
<< polycont >>
rect -19 296 15 375
rect -10 21 24 55
<< locali >>
rect 62 542 86 576
rect 122 542 146 576
rect 62 540 146 542
rect 62 504 86 540
rect 122 519 146 540
rect 122 504 220 519
rect 62 485 220 504
rect 62 444 146 450
rect 58 442 150 444
rect 58 408 74 442
rect 134 408 150 442
rect 58 406 150 408
rect -19 386 15 391
rect 184 352 220 485
rect 50 350 220 352
rect 50 316 74 350
rect 134 316 220 350
rect 50 314 220 316
rect 58 226 74 260
rect 134 226 150 260
rect 62 98 146 226
rect -10 55 24 76
rect 58 64 74 98
rect 134 64 150 98
rect 62 58 146 64
rect -10 0 24 21
rect 58 -24 74 10
rect 134 -24 150 10
rect 62 -90 146 -24
rect 62 -124 86 -90
rect 122 -124 146 -90
rect 62 -130 146 -124
<< viali >>
rect 86 542 122 576
rect 74 408 134 442
rect -19 375 15 386
rect -19 352 15 375
rect -19 296 15 314
rect -19 280 15 296
rect 74 226 134 260
rect -15 21 -10 55
rect -10 21 19 55
rect 86 -124 122 -90
<< metal1 >>
rect 54 576 152 582
rect 54 542 86 576
rect 122 542 152 576
rect 54 536 152 542
rect 66 442 144 456
rect 66 408 74 442
rect 134 408 144 442
rect -25 386 25 398
rect -25 352 -19 386
rect 15 352 25 386
rect -25 314 25 352
rect -25 280 -19 314
rect 15 280 25 314
rect -25 272 25 280
rect -21 55 25 272
rect 66 260 144 408
rect 66 226 74 260
rect 134 226 144 260
rect 66 214 144 226
rect -21 21 -15 55
rect 19 21 25 55
rect -21 0 25 21
rect 56 -90 152 -84
rect 56 -124 86 -90
rect 122 -124 152 -90
rect 56 -130 152 -124
<< labels >>
flabel metal1 -21 0 25 398 0 FreeSans 160 0 0 0 in
port 4 nsew
flabel metal1 66 214 144 267 0 FreeSans 160 0 0 0 out
port 6 nsew
flabel metal1 54 536 152 582 0 FreeSans 160 0 0 0 VDD
port 7 nsew
flabel metal1 56 -130 152 -84 0 FreeSans 160 0 0 0 VSS
port 9 nsew
<< end >>
