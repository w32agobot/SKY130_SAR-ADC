magic
tech sky130A
timestamp 1662997094
<< nwell >>
rect 0 253 47 440
rect 451 253 502 440
<< locali >>
rect 57 443 74 502
rect 427 443 444 502
rect 57 0 74 64
rect 174 0 191 64
rect 210 0 227 64
rect 284 0 301 64
rect 427 0 444 64
<< metal1 >>
rect 0 399 47 427
rect 451 399 502 427
rect 0 370 47 385
rect 451 370 502 385
rect 0 256 47 270
rect 451 256 502 270
rect 0 215 47 229
rect 451 215 502 229
rect 0 187 47 201
rect 451 187 502 201
rect 0 110 47 124
rect 451 110 502 124
rect 0 68 47 96
rect 451 68 502 96
<< metal4 >>
rect 236 456 266 467
rect 236 0 266 5
use adc_array_circuit_150n_Gate  adc_array_circuit_150n_0 ../adc_array_circuit
timestamp 1662997094
transform 1 0 -70 0 1 -221
box 117 285 521 664
use adc_array_wafflecap_8_Gate_25um2  adc_array_wafflecap_8_Gate_25um2_0 ../adc_array_topologies/adc_array_wafflecap_8_topA
timestamp 1662997094
transform 1 0 0 0 1 0
box 0 0 502 502
<< labels >>
rlabel metal1 0 370 0 385 7 sample_n
port 2 w
rlabel metal1 0 256 0 270 7 colon_n
port 3 w
rlabel metal1 0 215 0 229 7 col_n
port 4 w
rlabel metal1 0 187 0 201 7 sample
port 5 w
rlabel metal1 0 110 0 124 7 vcom
port 6 w
rlabel metal1 0 68 0 96 7 VSS
port 7 w
rlabel locali 427 0 444 0 5 row_n
port 8 s
rlabel locali 174 0 191 0 5 sw_n
port 9 s
rlabel locali 284 0 301 0 5 sw
port 11 s
rlabel metal1 0 399 0 427 7 VDD
port 13 w
rlabel locali 210 0 227 0 5 in
port 10 s
rlabel metal4 236 0 266 0 5 ctop
port 14 s
<< end >>
