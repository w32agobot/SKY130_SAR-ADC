magic
tech sky130A
magscale 1 2
timestamp 1661174986
<< error_s >>
rect 182 -1326 240 -1320
rect 374 -1326 432 -1320
rect 566 -1326 624 -1320
rect 758 -1326 816 -1320
rect 182 -1360 194 -1326
rect 374 -1360 386 -1326
rect 566 -1360 578 -1326
rect 758 -1360 770 -1326
rect 182 -1366 240 -1360
rect 374 -1366 432 -1360
rect 566 -1366 624 -1360
rect 758 -1366 816 -1360
rect 86 -1536 144 -1530
rect 278 -1536 336 -1530
rect 470 -1536 528 -1530
rect 662 -1536 720 -1530
rect 86 -1570 98 -1536
rect 278 -1570 290 -1536
rect 470 -1570 482 -1536
rect 662 -1570 674 -1536
rect 86 -1576 144 -1570
rect 278 -1576 336 -1570
rect 470 -1576 528 -1570
rect 662 -1576 720 -1570
<< nwell >>
rect -50 -292 848 8
<< nmos >>
rect 48 -910 78 -510
rect 144 -910 174 -510
rect 240 -910 270 -510
rect 336 -910 366 -510
rect 432 -910 462 -510
rect 528 -910 558 -510
rect 624 -910 654 -510
rect 720 -910 750 -510
<< pmos >>
rect 48 -192 78 -92
rect 144 -192 174 -92
rect 240 -192 270 -92
rect 336 -192 366 -92
rect 432 -192 462 -92
rect 528 -192 558 -92
rect 624 -192 654 -92
rect 720 -192 750 -92
<< ndiff >>
rect -14 -522 48 -510
rect -14 -898 -2 -522
rect 32 -898 48 -522
rect -14 -910 48 -898
rect 78 -522 144 -510
rect 78 -898 94 -522
rect 128 -898 144 -522
rect 78 -910 144 -898
rect 174 -522 240 -510
rect 174 -898 190 -522
rect 224 -898 240 -522
rect 174 -910 240 -898
rect 270 -522 336 -510
rect 270 -898 286 -522
rect 320 -898 336 -522
rect 270 -910 336 -898
rect 366 -522 432 -510
rect 366 -898 382 -522
rect 416 -898 432 -522
rect 366 -910 432 -898
rect 462 -522 528 -510
rect 462 -898 478 -522
rect 512 -898 528 -522
rect 462 -910 528 -898
rect 558 -522 624 -510
rect 558 -898 574 -522
rect 608 -898 624 -522
rect 558 -910 624 -898
rect 654 -522 720 -510
rect 654 -898 670 -522
rect 704 -898 720 -522
rect 654 -910 720 -898
rect 750 -522 812 -510
rect 750 -898 766 -522
rect 800 -898 812 -522
rect 750 -910 812 -898
<< pdiff >>
rect -14 -104 48 -92
rect -14 -180 -2 -104
rect 32 -180 48 -104
rect -14 -192 48 -180
rect 78 -104 144 -92
rect 78 -180 94 -104
rect 128 -180 144 -104
rect 78 -192 144 -180
rect 174 -104 240 -92
rect 174 -180 190 -104
rect 224 -180 240 -104
rect 174 -192 240 -180
rect 270 -104 336 -92
rect 270 -180 286 -104
rect 320 -180 336 -104
rect 270 -192 336 -180
rect 366 -104 432 -92
rect 366 -180 382 -104
rect 416 -180 432 -104
rect 366 -192 432 -180
rect 462 -104 528 -92
rect 462 -180 478 -104
rect 512 -180 528 -104
rect 462 -192 528 -180
rect 558 -104 624 -92
rect 558 -180 574 -104
rect 608 -180 624 -104
rect 558 -192 624 -180
rect 654 -104 720 -92
rect 654 -180 670 -104
rect 704 -180 720 -104
rect 654 -192 720 -180
rect 750 -104 812 -92
rect 750 -180 766 -104
rect 800 -180 812 -104
rect 750 -192 812 -180
<< ndiffc >>
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
<< pdiffc >>
rect -2 -180 32 -104
rect 94 -180 128 -104
rect 190 -180 224 -104
rect 286 -180 320 -104
rect 382 -180 416 -104
rect 478 -180 512 -104
rect 574 -180 608 -104
rect 670 -180 704 -104
rect 766 -180 800 -104
<< poly >>
rect 48 -92 78 -66
rect 144 -92 174 -66
rect 240 -92 270 -66
rect 336 -92 366 -66
rect 432 -92 462 -66
rect 528 -92 558 -66
rect 624 -92 654 -66
rect 720 -92 750 -66
rect 48 -218 78 -192
rect 144 -218 174 -192
rect 240 -218 270 -192
rect 336 -218 366 -192
rect 432 -218 462 -192
rect 528 -218 558 -192
rect 624 -218 654 -192
rect 720 -218 750 -192
rect 48 -250 750 -218
rect 48 -510 78 -484
rect 144 -510 174 -484
rect 240 -510 270 -484
rect 336 -510 366 -484
rect 432 -510 462 -484
rect 528 -510 558 -484
rect 624 -510 654 -484
rect 720 -510 750 -484
rect 48 -938 78 -910
rect 144 -938 174 -910
rect 240 -938 270 -910
rect 336 -938 366 -910
rect 48 -968 366 -938
rect 432 -938 462 -910
rect 528 -938 558 -910
rect 624 -938 654 -910
rect 720 -938 750 -910
rect 432 -968 750 -938
<< locali >>
rect -2 -54 800 -20
rect -2 -104 32 -54
rect -2 -196 32 -180
rect 94 -104 128 -88
rect 94 -256 128 -180
rect 190 -104 224 -54
rect 190 -196 224 -180
rect 286 -104 320 -88
rect 286 -256 320 -180
rect 382 -104 416 -54
rect 382 -196 416 -180
rect 478 -104 512 -88
rect 94 -290 320 -256
rect 286 -438 320 -290
rect 94 -472 320 -438
rect -2 -522 32 -506
rect -2 -972 32 -898
rect 94 -522 128 -472
rect 94 -938 128 -898
rect 190 -522 224 -506
rect 190 -972 224 -898
rect 286 -522 320 -472
rect 478 -252 512 -180
rect 574 -104 608 -54
rect 574 -196 608 -180
rect 670 -104 704 -88
rect 670 -252 704 -180
rect 766 -104 800 -54
rect 766 -196 800 -180
rect 478 -286 704 -252
rect 478 -438 512 -286
rect 478 -472 704 -438
rect 286 -938 320 -898
rect 382 -522 416 -506
rect 382 -972 416 -898
rect 478 -522 512 -472
rect 478 -938 512 -898
rect 574 -522 608 -506
rect 574 -972 608 -898
rect 670 -522 704 -472
rect 670 -938 704 -898
rect 766 -522 800 -506
rect 766 -972 800 -898
rect -2 -1006 800 -972
<< viali >>
rect -2 -180 32 -104
rect 94 -180 128 -104
rect 190 -180 224 -104
rect 286 -180 320 -104
rect 382 -180 416 -104
rect 478 -180 512 -104
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 574 -180 608 -104
rect 670 -180 704 -104
rect 766 -180 800 -104
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
<< metal1 >>
rect -8 -104 38 -92
rect -8 -180 -2 -104
rect 32 -180 38 -104
rect -8 -192 38 -180
rect 88 -104 134 -92
rect 88 -180 94 -104
rect 128 -180 134 -104
rect 88 -192 134 -180
rect 184 -104 230 -92
rect 184 -180 190 -104
rect 224 -180 230 -104
rect 184 -192 230 -180
rect 280 -104 326 -92
rect 280 -180 286 -104
rect 320 -180 326 -104
rect 280 -192 326 -180
rect 376 -104 422 -92
rect 376 -180 382 -104
rect 416 -180 422 -104
rect 376 -192 422 -180
rect 472 -104 518 -92
rect 472 -180 478 -104
rect 512 -180 518 -104
rect 472 -192 518 -180
rect 568 -104 614 -92
rect 568 -180 574 -104
rect 608 -180 614 -104
rect 568 -192 614 -180
rect 664 -104 710 -92
rect 664 -180 670 -104
rect 704 -180 710 -104
rect 664 -192 710 -180
rect 760 -104 806 -92
rect 760 -180 766 -104
rect 800 -180 806 -104
rect 760 -192 806 -180
rect -8 -522 38 -510
rect -8 -898 -2 -522
rect 32 -898 38 -522
rect -8 -910 38 -898
rect 88 -522 134 -510
rect 88 -898 94 -522
rect 128 -898 134 -522
rect 88 -910 134 -898
rect 184 -522 230 -510
rect 184 -898 190 -522
rect 224 -898 230 -522
rect 184 -910 230 -898
rect 280 -522 326 -510
rect 280 -898 286 -522
rect 320 -898 326 -522
rect 280 -910 326 -898
rect 376 -522 422 -510
rect 376 -898 382 -522
rect 416 -898 422 -522
rect 376 -910 422 -898
rect 472 -522 518 -510
rect 472 -898 478 -522
rect 512 -898 518 -522
rect 472 -910 518 -898
rect 568 -522 614 -510
rect 568 -898 574 -522
rect 608 -898 614 -522
rect 568 -910 614 -898
rect 664 -522 710 -510
rect 664 -898 670 -522
rect 704 -898 710 -522
rect 664 -910 710 -898
rect 760 -522 806 -510
rect 760 -898 766 -522
rect 800 -898 806 -522
rect 760 -910 806 -898
use sky130_fd_pr__nfet_01v8_2A3UGD  sky130_fd_pr__nfet_01v8_2A3UGD_0
timestamp 1661174986
transform 1 0 451 0 1 -1448
box -413 -138 413 138
<< end >>
