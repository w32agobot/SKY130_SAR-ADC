magic
tech sky130A
timestamp 1659615172
<< metal2 >>
rect 16 481 486 486
rect 16 453 21 481
rect 49 453 69 481
rect 97 453 117 481
rect 145 453 165 481
rect 193 453 213 481
rect 241 453 261 481
rect 289 453 309 481
rect 337 453 357 481
rect 385 453 405 481
rect 433 453 453 481
rect 481 453 486 481
rect 16 433 486 453
rect 16 405 21 433
rect 49 405 165 433
rect 193 405 309 433
rect 337 405 453 433
rect 481 405 486 433
rect 16 385 486 405
rect 16 357 21 385
rect 49 357 165 385
rect 193 357 309 385
rect 337 357 453 385
rect 481 357 486 385
rect 16 337 486 357
rect 16 309 21 337
rect 49 309 69 337
rect 97 309 117 337
rect 145 309 165 337
rect 193 309 213 337
rect 241 309 261 337
rect 289 309 309 337
rect 337 309 357 337
rect 385 309 405 337
rect 433 309 453 337
rect 481 309 486 337
rect 16 304 486 309
rect 16 289 198 304
rect 16 261 21 289
rect 49 261 165 289
rect 193 261 198 289
rect 304 289 486 304
rect 16 241 198 261
rect 16 213 21 241
rect 49 213 165 241
rect 193 213 198 241
rect 230 230 272 272
rect 304 261 309 289
rect 337 261 453 289
rect 481 261 486 289
rect 304 241 486 261
rect 16 198 198 213
rect 304 213 309 241
rect 337 213 453 241
rect 481 213 486 241
rect 304 198 486 213
rect 16 193 486 198
rect 16 165 21 193
rect 49 165 69 193
rect 97 165 117 193
rect 145 165 165 193
rect 193 165 213 193
rect 241 165 261 193
rect 289 165 309 193
rect 337 165 357 193
rect 385 165 405 193
rect 433 165 453 193
rect 481 165 486 193
rect 16 145 486 165
rect 16 117 21 145
rect 49 117 165 145
rect 193 117 309 145
rect 337 117 453 145
rect 481 117 486 145
rect 16 97 486 117
rect 16 69 21 97
rect 49 69 165 97
rect 193 69 309 97
rect 337 69 453 97
rect 481 69 486 97
rect 16 49 486 69
rect 16 21 21 49
rect 49 21 69 49
rect 97 21 117 49
rect 145 21 165 49
rect 193 21 213 49
rect 241 21 261 49
rect 289 21 309 49
rect 337 21 357 49
rect 385 21 405 49
rect 433 21 453 49
rect 481 21 486 49
rect 16 16 486 21
<< via2 >>
rect 21 453 49 481
rect 69 453 97 481
rect 117 453 145 481
rect 165 453 193 481
rect 213 453 241 481
rect 261 453 289 481
rect 309 453 337 481
rect 357 453 385 481
rect 405 453 433 481
rect 453 453 481 481
rect 21 405 49 433
rect 165 405 193 433
rect 309 405 337 433
rect 453 405 481 433
rect 21 357 49 385
rect 165 357 193 385
rect 309 357 337 385
rect 453 357 481 385
rect 21 309 49 337
rect 69 309 97 337
rect 117 309 145 337
rect 165 309 193 337
rect 213 309 241 337
rect 261 309 289 337
rect 309 309 337 337
rect 357 309 385 337
rect 405 309 433 337
rect 453 309 481 337
rect 21 261 49 289
rect 165 261 193 289
rect 21 213 49 241
rect 165 213 193 241
rect 309 261 337 289
rect 453 261 481 289
rect 309 213 337 241
rect 453 213 481 241
rect 21 165 49 193
rect 69 165 97 193
rect 117 165 145 193
rect 165 165 193 193
rect 213 165 241 193
rect 261 165 289 193
rect 309 165 337 193
rect 357 165 385 193
rect 405 165 433 193
rect 453 165 481 193
rect 21 117 49 145
rect 165 117 193 145
rect 309 117 337 145
rect 453 117 481 145
rect 21 69 49 97
rect 165 69 193 97
rect 309 69 337 97
rect 453 69 481 97
rect 21 21 49 49
rect 69 21 97 49
rect 117 21 145 49
rect 165 21 193 49
rect 213 21 241 49
rect 261 21 289 49
rect 309 21 337 49
rect 357 21 385 49
rect 405 21 433 49
rect 453 21 481 49
<< metal3 >>
rect 18 481 484 484
rect 18 453 21 481
rect 49 453 69 481
rect 97 453 117 481
rect 145 453 165 481
rect 193 453 213 481
rect 241 453 261 481
rect 289 453 309 481
rect 337 453 357 481
rect 385 453 405 481
rect 433 453 453 481
rect 481 453 484 481
rect 18 450 484 453
rect 18 433 52 450
rect 18 405 21 433
rect 49 405 52 433
rect 162 433 196 450
rect 18 385 52 405
rect 18 357 21 385
rect 49 357 52 385
rect 82 412 132 420
rect 82 378 90 412
rect 124 378 132 412
rect 82 370 132 378
rect 162 405 165 433
rect 193 405 196 433
rect 306 433 340 450
rect 162 385 196 405
rect 18 340 52 357
rect 162 357 165 385
rect 193 357 196 385
rect 226 412 276 420
rect 226 378 234 412
rect 268 378 276 412
rect 226 370 276 378
rect 306 405 309 433
rect 337 405 340 433
rect 450 433 484 450
rect 306 385 340 405
rect 162 340 196 357
rect 306 357 309 385
rect 337 357 340 385
rect 370 412 420 420
rect 370 378 378 412
rect 412 378 420 412
rect 370 370 420 378
rect 450 405 453 433
rect 481 405 484 433
rect 450 385 484 405
rect 306 340 340 357
rect 450 357 453 385
rect 481 357 484 385
rect 450 340 484 357
rect 18 337 484 340
rect 18 309 21 337
rect 49 309 69 337
rect 97 309 117 337
rect 145 309 165 337
rect 193 309 213 337
rect 241 309 261 337
rect 289 309 309 337
rect 337 309 357 337
rect 385 309 405 337
rect 433 309 453 337
rect 481 309 484 337
rect 18 306 484 309
rect 18 289 52 306
rect 18 261 21 289
rect 49 261 52 289
rect 162 289 196 306
rect 18 241 52 261
rect 18 213 21 241
rect 49 213 52 241
rect 82 268 132 276
rect 82 234 90 268
rect 124 234 132 268
rect 82 226 132 234
rect 162 261 165 289
rect 193 261 196 289
rect 162 241 196 261
rect 18 196 52 213
rect 162 213 165 241
rect 193 213 196 241
rect 162 196 196 213
rect 306 289 340 306
rect 306 261 309 289
rect 337 261 340 289
rect 450 289 484 306
rect 306 241 340 261
rect 306 213 309 241
rect 337 213 340 241
rect 370 268 420 276
rect 370 234 378 268
rect 412 234 420 268
rect 370 226 420 234
rect 450 261 453 289
rect 481 261 484 289
rect 450 241 484 261
rect 306 196 340 213
rect 450 213 453 241
rect 481 213 484 241
rect 450 196 484 213
rect 18 193 484 196
rect 18 165 21 193
rect 49 165 69 193
rect 97 165 117 193
rect 145 165 165 193
rect 193 165 213 193
rect 241 165 261 193
rect 289 165 309 193
rect 337 165 357 193
rect 385 165 405 193
rect 433 165 453 193
rect 481 165 484 193
rect 18 162 484 165
rect 18 145 52 162
rect 18 117 21 145
rect 49 117 52 145
rect 162 145 196 162
rect 18 97 52 117
rect 18 69 21 97
rect 49 69 52 97
rect 82 124 132 132
rect 82 90 90 124
rect 124 90 132 124
rect 82 82 132 90
rect 162 117 165 145
rect 193 117 196 145
rect 306 145 340 162
rect 162 97 196 117
rect 18 52 52 69
rect 162 69 165 97
rect 193 69 196 97
rect 226 124 276 132
rect 226 90 234 124
rect 268 90 276 124
rect 226 82 276 90
rect 306 117 309 145
rect 337 117 340 145
rect 450 145 484 162
rect 306 97 340 117
rect 162 52 196 69
rect 306 69 309 97
rect 337 69 340 97
rect 370 124 420 132
rect 370 90 378 124
rect 412 90 420 124
rect 370 82 420 90
rect 450 117 453 145
rect 481 117 484 145
rect 450 97 484 117
rect 306 52 340 69
rect 450 69 453 97
rect 481 69 484 97
rect 450 52 484 69
rect 18 49 484 52
rect 18 21 21 49
rect 49 21 69 49
rect 97 21 117 49
rect 145 21 165 49
rect 193 21 213 49
rect 241 21 261 49
rect 289 21 309 49
rect 337 21 357 49
rect 385 21 405 49
rect 433 21 453 49
rect 481 21 484 49
rect 18 18 484 21
<< via3 >>
rect 90 378 124 412
rect 234 378 268 412
rect 378 378 412 412
rect 90 234 124 268
rect 378 234 412 268
rect 90 90 124 124
rect 234 90 268 124
rect 378 90 412 124
<< metal4 >>
rect 92 420 122 467
rect 236 420 266 467
rect 380 420 410 467
rect 82 412 132 420
rect 82 410 90 412
rect 35 380 90 410
rect 82 378 90 380
rect 124 410 132 412
rect 226 412 276 420
rect 226 410 234 412
rect 124 380 234 410
rect 124 378 132 380
rect 82 370 132 378
rect 226 378 234 380
rect 268 410 276 412
rect 370 412 420 420
rect 370 410 378 412
rect 268 380 378 410
rect 268 378 276 380
rect 226 370 276 378
rect 370 378 378 380
rect 412 410 420 412
rect 412 380 467 410
rect 412 378 420 380
rect 370 370 420 378
rect 92 276 122 370
rect 236 323 266 370
rect 380 276 410 370
rect 82 268 132 276
rect 82 266 90 268
rect 35 236 90 266
rect 82 234 90 236
rect 124 266 132 268
rect 370 268 420 276
rect 370 266 378 268
rect 124 236 179 266
rect 323 236 378 266
rect 124 234 132 236
rect 82 226 132 234
rect 370 234 378 236
rect 412 266 420 268
rect 412 236 467 266
rect 412 234 420 236
rect 370 226 420 234
rect 92 132 122 226
rect 236 132 266 179
rect 380 132 410 226
rect 82 124 132 132
rect 82 122 90 124
rect 35 92 90 122
rect 82 90 90 92
rect 124 122 132 124
rect 226 124 276 132
rect 226 122 234 124
rect 124 92 234 122
rect 124 90 132 92
rect 82 82 132 90
rect 226 90 234 92
rect 268 122 276 124
rect 370 124 420 132
rect 370 122 378 124
rect 268 92 378 122
rect 268 90 276 92
rect 226 82 276 90
rect 370 90 378 92
rect 412 122 420 124
rect 412 92 467 122
rect 412 90 420 92
rect 370 82 420 90
rect 92 35 122 82
rect 236 35 266 82
rect 380 35 410 82
<< comment >>
rect 0 486 16 502
rect 486 486 502 502
rect 288 288 304 304
rect 272 272 288 288
rect 214 214 230 230
rect 198 198 214 214
rect 0 0 16 16
rect 486 0 502 16
<< labels >>
rlabel metal2 272 230 272 230 3 symmetry_metal
<< end >>
