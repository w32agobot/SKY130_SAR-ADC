* SPICE3 file created from extract.ext - technology: sky130A

C0 bot_2 m4_9804_1296# 3.18fF
C1 bot_1 dummy_bot 12.54fF
C2 bot_2 dummy_bot 15.18fF
C3 bot_1 m4_13284_1296# 3.32fF
C4 top_4 bot_4 32.39fF
C5 top_8 bot_8 29.82fF
C6 dummy_bot dummy_top 268.14fF
C7 dummy_bot m2_13252_2292# 2.62fF
C8 bot_1 m2_13252_2292# 2.64fF
C9 bot_4 m4_6324_1296# 2.12fF
C10 bot_4 dummy_bot 15.20fF
C11 bot_8 dummy_bot 12.90fF
C12 bot_1 top_1 30.55fF
C13 m2_13252_2292# dummy_top 4.41fF
C14 bot_2 top_2 31.20fF
C15 dummy_top VSUBS 3.66fF
C16 bot_1 VSUBS 2.40fF
C17 bot_2 VSUBS 2.40fF
C18 bot_4 VSUBS 2.40fF
C19 bot_8 VSUBS 2.07fF
C20 dummy_bot VSUBS 33.73fF
