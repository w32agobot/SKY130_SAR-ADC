** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_vcm_generator.sch
.subckt adc_vcm_generator VDD VSS clk vcm
*.PININFO VDD:B VSS:B clk:I vcm:B
X1 clk VDD VSS phi1_n phi1 phi2 phi2_n adc_vcm_clkgen
x_decap_1 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x_decap_2 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x_decap_3 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
X2 phi2_n VDD phi2 mimtop1 VDD VSS adc_vcm_switch
x_cap1_1 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_2 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_3 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_4 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_5 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_6 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_7 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_8 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_9 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_10 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_11 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_12 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_13 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_14 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_15 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_16 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_17 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_18 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_19 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_20 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_21 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_22 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_23 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_24 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_25 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_26 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_27 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_28 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_29 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_30 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_31 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_32 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_33 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_34 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_35 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_36 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_37 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_38 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_39 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap1_40 mimtop1 mimbot1 vcm VSS VSS adc_noise_decoup_cell1
x_cap2_1 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_2 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_3 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_4 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_5 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_6 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_7 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_8 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_9 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_10 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_11 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_12 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_13 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_14 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_15 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_16 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_17 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_18 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_19 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_20 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_21 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_22 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_23 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_24 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_25 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_26 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_27 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_28 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_29 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_30 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_31 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_32 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_33 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_34 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_35 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_36 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_37 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_38 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_39 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
x_cap2_40 mimtop2 VSS vcm VSS VSS adc_noise_decoup_cell1
X4 phi1_n mimbot1 phi1 VSS VDD VSS adc_vcm_switch
X3 phi2_n mimbot1 phi2 mimtop2 VDD VSS adc_vcm_switch
X6 phi1_n mimtop2 phi1 vcm VDD VSS adc_vcm_switch
X5 phi1_n mimtop1 phi1 vcm VDD VSS adc_vcm_switch
**** begin user architecture code

.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
.ends

* expanding   symbol:  adc_vcm_clkgen.sym # of pins=7
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_vcm_clkgen.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_vcm_clkgen.sch
.subckt adc_vcm_clkgen clk VDD VSS phi1_n phi1 phi2 phi2_n
*.PININFO VDD:B VSS:B phi2_n:O phi2:O phi1:O phi1_n:O clk:I
x23 clk VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x2 net6 VSS VSS VDD VDD phi1 sky130_fd_sc_hd__buf_4
x5 net6 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_1
x11 net11 VSS VSS VDD VDD net6 sky130_fd_sc_hd__inv_1
x12 net7 VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_1
x4 net3 VSS VSS VDD VDD phi1_n sky130_fd_sc_hd__buf_4
x7 net4 VSS VSS VDD VDD phi2_n sky130_fd_sc_hd__buf_4
x8 net7 VSS VSS VDD VDD phi2 sky130_fd_sc_hd__buf_4
x3 net1 VSS VSS VDD VDD net8 sky130_fd_sc_hd__dlymetal6s6s_1
x10 net2 VSS VSS VDD VDD net9 sky130_fd_sc_hd__dlymetal6s6s_1
x6 net8 VSS VSS VDD VDD net10 sky130_fd_sc_hd__dlymetal6s6s_1
x13 net9 VSS VSS VDD VDD net13 sky130_fd_sc_hd__dlymetal6s6s_1
x1 net12 VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
x9 net10 VSS VSS VDD VDD net11 sky130_fd_sc_hd__dlymetal6s6s_1
x14 net13 VSS VSS VDD VDD net12 sky130_fd_sc_hd__dlymetal6s6s_1
x15 clk net4 VSS VSS VDD VDD net1 sky130_fd_sc_hd__nand2_1
x16 net3 net5 VSS VSS VDD VDD net2 sky130_fd_sc_hd__nand2_1
.ends


* expanding   symbol:  adc_noise_decoup_cell1.sym # of pins=5
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_noise_decoup_cell1.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_noise_decoup_cell1.sch
.subckt adc_noise_decoup_cell1 mimcap_top mimcap_bot nmoscap_top nmoscap_bot pwell
*.PININFO nmoscap_top:B mimcap_top:B mimcap_bot:B nmoscap_bot:B pwell:B
XC1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 W=17.2 L=17.2 MF=1 m=1
XM1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 L=16.0 W=16.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_vcm_switch.sym # of pins=6
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_vcm_switch.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_vcm_switch.sch
.subckt adc_vcm_switch sw_n a sw b VDD VSS
*.PININFO VSS:B VDD:B sw_n:I sw:I a:B b:B
XM1 a sw_n b VDD sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 a sw b VSS sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
