magic
tech sky130A
magscale 1 2
timestamp 1661177810
<< error_p >>
rect -2389 -700 -2329 700
rect -2309 -700 -2249 700
rect -70 -700 -10 700
rect 10 -700 70 700
rect 2249 -700 2309 700
rect 2329 -700 2389 700
<< metal3 >>
rect -4628 672 -2329 700
rect -4628 -672 -2413 672
rect -2349 -672 -2329 672
rect -4628 -700 -2329 -672
rect -2309 672 -10 700
rect -2309 -672 -94 672
rect -30 -672 -10 672
rect -2309 -700 -10 -672
rect 10 672 2309 700
rect 10 -672 2225 672
rect 2289 -672 2309 672
rect 10 -700 2309 -672
rect 2329 672 4628 700
rect 2329 -672 4544 672
rect 4608 -672 4628 672
rect 2329 -700 4628 -672
<< via3 >>
rect -2413 -672 -2349 672
rect -94 -672 -30 672
rect 2225 -672 2289 672
rect 4544 -672 4608 672
<< mimcap >>
rect -4528 560 -2528 600
rect -4528 -560 -4488 560
rect -2568 -560 -2528 560
rect -4528 -600 -2528 -560
rect -2209 560 -209 600
rect -2209 -560 -2169 560
rect -249 -560 -209 560
rect -2209 -600 -209 -560
rect 110 560 2110 600
rect 110 -560 150 560
rect 2070 -560 2110 560
rect 110 -600 2110 -560
rect 2429 560 4429 600
rect 2429 -560 2469 560
rect 4389 -560 4429 560
rect 2429 -600 4429 -560
<< mimcapcontact >>
rect -4488 -560 -2568 560
rect -2169 -560 -249 560
rect 150 -560 2070 560
rect 2469 -560 4389 560
<< metal4 >>
rect -2429 672 -2333 688
rect -4489 560 -2567 561
rect -4489 -560 -4488 560
rect -2568 -560 -2567 560
rect -4489 -561 -2567 -560
rect -2429 -672 -2413 672
rect -2349 -672 -2333 672
rect -110 672 -14 688
rect -2170 560 -248 561
rect -2170 -560 -2169 560
rect -249 -560 -248 560
rect -2170 -561 -248 -560
rect -2429 -688 -2333 -672
rect -110 -672 -94 672
rect -30 -672 -14 672
rect 2209 672 2305 688
rect 149 560 2071 561
rect 149 -560 150 560
rect 2070 -560 2071 560
rect 149 -561 2071 -560
rect -110 -688 -14 -672
rect 2209 -672 2225 672
rect 2289 -672 2305 672
rect 4528 672 4624 688
rect 2468 560 4390 561
rect 2468 -560 2469 560
rect 4389 -560 4390 560
rect 2468 -561 4390 -560
rect 2209 -688 2305 -672
rect 4528 -672 4544 672
rect 4608 -672 4624 672
rect 4528 -688 4624 -672
<< properties >>
string FIXED_BBOX 2329 -700 4529 700
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 6 val 126.08 carea 2.00 cperi 0.19 nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
