* SPICE3 file created from extract.ext - technology: sky130A

C0 top_4 dummy_bot 8.18fF
C1 top_2 bot_2 19.51fF
C2 top_1 dummy_top 2.71fF
C3 top_8 dummy_bot 6.72fF
C4 dummy_top bot_1 2.83fF
C5 top_2 shielding 11.17fF
C6 shielding bot_2 24.19fF
C7 top_1 dummy_bot 6.98fF
C8 bot_8 shielding 20.80fF
C9 top_2 dummy_top 2.74fF
C10 dummy_top bot_2 2.46fF
C11 bot_4 shielding 24.18fF
C12 top_1 bot_1 19.13fF
C13 dummy_top shielding 52.57fF
C14 top_4 shielding 11.59fF
C15 top_2 dummy_bot 7.44fF
C16 top_8 shielding 10.53fF
C17 top_4 bot_4 20.23fF
C18 dummy_bot shielding 183.35fF
C19 dummy_top top_4 2.86fF
C20 top_8 bot_8 18.69fF
C21 dummy_bot bot_8 2.08fF
C22 top_1 shielding 10.96fF
C23 dummy_top top_8 2.61fF
C24 shielding bot_1 24.56fF
C25 dummy_top dummy_bot 136.37fF
C26 dummy_top VSUBS 3.62fF
C27 shielding VSUBS 61.66fF
C28 bot_1 VSUBS 2.68fF
C29 bot_2 VSUBS 2.71fF
C30 bot_4 VSUBS 2.71fF
C31 bot_8 VSUBS 2.30fF
C32 dummy_bot VSUBS 27.97fF
