VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_clkgen_with_edgedetect
  CLASS BLOCK ;
  FOREIGN adc_clkgen_with_edgedetect ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 64.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 22.720 2.480 24.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.720 2.480 48.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.720 2.480 72.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.720 2.480 96.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.720 2.480 120.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 142.720 2.480 144.320 60.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.720 2.480 18.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.720 2.480 42.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 2.480 66.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.720 2.480 90.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.720 2.480 114.320 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.720 2.480 138.320 60.080 ;
    END
  END VPWR
  PIN clk_comp_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 15.680 160.000 16.280 ;
    END
  END clk_comp_out
  PIN clk_dig_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END clk_dig_out
  PIN dlycontrol1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END dlycontrol1_in[0]
  PIN dlycontrol1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END dlycontrol1_in[1]
  PIN dlycontrol1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END dlycontrol1_in[2]
  PIN dlycontrol1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END dlycontrol1_in[3]
  PIN dlycontrol1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END dlycontrol1_in[4]
  PIN dlycontrol2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END dlycontrol2_in[0]
  PIN dlycontrol2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END dlycontrol2_in[1]
  PIN dlycontrol2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END dlycontrol2_in[2]
  PIN dlycontrol2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END dlycontrol2_in[3]
  PIN dlycontrol2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END dlycontrol2_in[4]
  PIN dlycontrol3_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END dlycontrol3_in[0]
  PIN dlycontrol3_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END dlycontrol3_in[1]
  PIN dlycontrol3_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END dlycontrol3_in[2]
  PIN dlycontrol3_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END dlycontrol3_in[3]
  PIN dlycontrol3_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END dlycontrol3_in[4]
  PIN dlycontrol4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END dlycontrol4_in[0]
  PIN dlycontrol4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END dlycontrol4_in[1]
  PIN dlycontrol4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END dlycontrol4_in[2]
  PIN dlycontrol4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END dlycontrol4_in[3]
  PIN dlycontrol4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END dlycontrol4_in[4]
  PIN dlycontrol4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END dlycontrol4_in[5]
  PIN ena_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END ena_in
  PIN enable_dlycontrol_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END enable_dlycontrol_in
  PIN ndecision_finish_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 47.640 160.000 48.240 ;
    END
  END ndecision_finish_in
  PIN nsample_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END nsample_n_in
  PIN nsample_n_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END nsample_n_out
  PIN nsample_p_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 60.000 100.190 64.000 ;
    END
  END nsample_p_in
  PIN nsample_p_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 60.000 140.210 64.000 ;
    END
  END nsample_p_out
  PIN sample_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END sample_n_in
  PIN sample_n_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END sample_n_out
  PIN sample_p_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 60.000 20.150 64.000 ;
    END
  END sample_p_in
  PIN sample_p_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 60.000 60.170 64.000 ;
    END
  END sample_p_out
  PIN start_conv_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END start_conv_in
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 154.100 59.925 ;
      LAYER met1 ;
        RECT 5.520 0.380 154.100 62.180 ;
      LAYER met2 ;
        RECT 7.910 59.720 19.590 62.210 ;
        RECT 20.430 59.720 59.610 62.210 ;
        RECT 60.450 59.720 99.630 62.210 ;
        RECT 100.470 59.720 139.650 62.210 ;
        RECT 140.490 59.720 150.780 62.210 ;
        RECT 7.910 4.280 150.780 59.720 ;
        RECT 7.910 0.350 19.590 4.280 ;
        RECT 20.430 0.350 59.610 4.280 ;
        RECT 60.450 0.350 99.630 4.280 ;
        RECT 100.470 0.350 139.650 4.280 ;
        RECT 140.490 0.350 150.780 4.280 ;
      LAYER met3 ;
        RECT 4.000 56.800 156.000 60.005 ;
        RECT 4.400 55.400 156.000 56.800 ;
        RECT 4.000 54.760 156.000 55.400 ;
        RECT 4.400 53.360 156.000 54.760 ;
        RECT 4.000 52.720 156.000 53.360 ;
        RECT 4.400 51.320 156.000 52.720 ;
        RECT 4.000 50.680 156.000 51.320 ;
        RECT 4.400 49.280 156.000 50.680 ;
        RECT 4.000 48.640 156.000 49.280 ;
        RECT 4.400 47.240 155.600 48.640 ;
        RECT 4.000 46.600 156.000 47.240 ;
        RECT 4.400 45.200 156.000 46.600 ;
        RECT 4.000 44.560 156.000 45.200 ;
        RECT 4.400 43.160 156.000 44.560 ;
        RECT 4.000 42.520 156.000 43.160 ;
        RECT 4.400 41.120 156.000 42.520 ;
        RECT 4.000 40.480 156.000 41.120 ;
        RECT 4.400 39.080 156.000 40.480 ;
        RECT 4.000 38.440 156.000 39.080 ;
        RECT 4.400 37.040 156.000 38.440 ;
        RECT 4.000 36.400 156.000 37.040 ;
        RECT 4.400 35.000 156.000 36.400 ;
        RECT 4.000 34.360 156.000 35.000 ;
        RECT 4.400 32.960 156.000 34.360 ;
        RECT 4.000 32.320 156.000 32.960 ;
        RECT 4.400 30.920 156.000 32.320 ;
        RECT 4.000 30.280 156.000 30.920 ;
        RECT 4.400 28.880 156.000 30.280 ;
        RECT 4.000 28.240 156.000 28.880 ;
        RECT 4.400 26.840 156.000 28.240 ;
        RECT 4.000 26.200 156.000 26.840 ;
        RECT 4.400 24.800 156.000 26.200 ;
        RECT 4.000 24.160 156.000 24.800 ;
        RECT 4.400 22.760 156.000 24.160 ;
        RECT 4.000 22.120 156.000 22.760 ;
        RECT 4.400 20.720 156.000 22.120 ;
        RECT 4.000 20.080 156.000 20.720 ;
        RECT 4.400 18.680 156.000 20.080 ;
        RECT 4.000 18.040 156.000 18.680 ;
        RECT 4.400 16.680 156.000 18.040 ;
        RECT 4.400 16.640 155.600 16.680 ;
        RECT 4.000 16.000 155.600 16.640 ;
        RECT 4.400 15.280 155.600 16.000 ;
        RECT 4.400 14.600 156.000 15.280 ;
        RECT 4.000 13.960 156.000 14.600 ;
        RECT 4.400 12.560 156.000 13.960 ;
        RECT 4.000 11.920 156.000 12.560 ;
        RECT 4.400 10.520 156.000 11.920 ;
        RECT 4.000 9.880 156.000 10.520 ;
        RECT 4.400 8.480 156.000 9.880 ;
        RECT 4.000 7.840 156.000 8.480 ;
        RECT 4.400 6.440 156.000 7.840 ;
        RECT 4.000 1.535 156.000 6.440 ;
      LAYER met4 ;
        RECT 34.335 8.335 34.665 14.105 ;
  END
END adc_clkgen_with_edgedetect
END LIBRARY

