** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Gate.sch
.subckt adc_array_wafflecap_8_Gate vcom VDD out VSS row_n col_n colon_n sample_n sample in sw sw_n
*.PININFO vcom:B VDD:B out:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I in:B sw:I sw_n:I
x1 VDD row_n col_n colon_n sample_n vcom sample VSS out in sw_n sw adc_array_circuit_150n_gate
.ends

* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_gate.sym # of pins=12
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_gate.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_gate.sch
.subckt adc_array_circuit_150n_gate  VDD row_n col_n colon_n sample_n vcom sample VSS out in sw_n sw
*.PININFO sw:I sw_n:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B sample:I sample_n:I in:B out:B
XM1 in sw_n out VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 in sw out VSS sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
