VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_top
  CLASS BLOCK ;
  FOREIGN adc_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 432.000 BY 403.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 399.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 434.020 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 397.680 434.020 399.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.420 3.280 434.020 399.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.720 -0.020 18.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.720 -0.020 42.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 -0.020 66.320 177.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 224.845 66.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.720 133.310 90.320 177.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.720 224.845 90.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.720 133.310 114.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.720 133.310 138.320 167.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.720 228.660 138.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 160.720 133.310 162.320 167.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 160.720 228.660 162.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 133.310 186.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 133.310 210.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.720 133.310 234.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.720 133.310 258.320 181.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.720 216.280 258.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 280.720 133.310 282.320 182.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 280.720 215.190 282.320 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.720 195.960 306.320 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.720 195.960 330.320 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 352.720 195.960 354.320 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 376.720 173.300 378.320 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.720 173.300 402.320 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.720 -0.020 426.320 402.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 34.080 89.800 35.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 58.080 89.800 59.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 82.080 89.800 83.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 106.080 89.800 107.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 130.080 89.800 131.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 154.080 437.320 155.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 178.080 437.320 179.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 202.080 437.320 203.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 226.080 437.320 227.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 250.080 437.320 251.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 274.080 89.800 275.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 298.080 89.800 299.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 322.080 89.800 323.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 346.080 89.800 347.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 370.080 437.320 371.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 34.080 437.320 35.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 58.080 437.320 59.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 82.080 437.320 83.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 106.080 437.320 107.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 130.080 437.320 131.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 274.080 437.320 275.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 298.080 437.320 299.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 322.080 437.320 323.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 346.080 437.320 347.680 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 402.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 437.320 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 400.980 437.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 435.720 -0.020 437.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.020 -0.020 21.620 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.020 -0.020 45.620 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.020 -0.020 69.620 177.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.020 224.845 69.620 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.020 133.310 93.620 167.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.020 228.660 93.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.020 133.310 117.620 167.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.020 228.660 117.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.020 133.310 141.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.020 133.310 165.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 133.310 189.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.020 133.310 213.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 236.020 133.310 237.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.020 133.310 261.620 182.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.020 215.190 261.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.020 133.310 285.620 181.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.020 216.280 285.620 267.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.020 195.960 309.620 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.020 195.960 333.620 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 356.020 195.960 357.620 226.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 380.020 173.300 381.620 226.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 37.380 89.800 38.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 61.380 89.800 62.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 85.380 89.800 86.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 109.380 89.800 110.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 133.380 437.320 134.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 157.380 437.320 158.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 181.380 437.320 182.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 205.380 437.320 206.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 229.380 437.320 230.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 253.380 437.320 254.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 277.380 89.800 278.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 301.380 89.800 302.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 325.380 89.800 326.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 349.380 89.800 350.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 373.380 437.320 374.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 37.380 437.320 38.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 61.380 437.320 62.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 85.380 437.320 86.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 109.380 437.320 110.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 277.380 437.320 278.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 301.380 437.320 302.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 325.380 437.320 326.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 259.560 349.380 437.320 350.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 418.260 10.640 419.860 391.920 ;
    END
  END VSS
  PIN clk_vcm
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 179.560 432.000 180.160 ;
    END
  END clk_vcm
  PIN config_1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END config_1_in[0]
  PIN config_1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END config_1_in[10]
  PIN config_1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END config_1_in[11]
  PIN config_1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END config_1_in[12]
  PIN config_1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END config_1_in[13]
  PIN config_1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END config_1_in[14]
  PIN config_1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END config_1_in[15]
  PIN config_1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END config_1_in[1]
  PIN config_1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END config_1_in[2]
  PIN config_1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END config_1_in[3]
  PIN config_1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END config_1_in[4]
  PIN config_1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END config_1_in[5]
  PIN config_1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END config_1_in[6]
  PIN config_1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END config_1_in[7]
  PIN config_1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END config_1_in[8]
  PIN config_1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END config_1_in[9]
  PIN config_2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END config_2_in[0]
  PIN config_2_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END config_2_in[10]
  PIN config_2_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END config_2_in[11]
  PIN config_2_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END config_2_in[12]
  PIN config_2_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END config_2_in[13]
  PIN config_2_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END config_2_in[14]
  PIN config_2_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END config_2_in[15]
  PIN config_2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END config_2_in[1]
  PIN config_2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END config_2_in[2]
  PIN config_2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END config_2_in[3]
  PIN config_2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END config_2_in[4]
  PIN config_2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END config_2_in[5]
  PIN config_2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END config_2_in[6]
  PIN config_2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END config_2_in[7]
  PIN config_2_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END config_2_in[8]
  PIN config_2_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END config_2_in[9]
  PIN conversion_finished_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END conversion_finished_out
  PIN dummypin[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 390.360 432.000 390.960 ;
    END
  END dummypin[0]
  PIN dummypin[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 116.320 432.000 116.920 ;
    END
  END dummypin[10]
  PIN dummypin[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 95.240 432.000 95.840 ;
    END
  END dummypin[11]
  PIN dummypin[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 74.160 432.000 74.760 ;
    END
  END dummypin[12]
  PIN dummypin[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 53.080 432.000 53.680 ;
    END
  END dummypin[13]
  PIN dummypin[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 32.000 432.000 32.600 ;
    END
  END dummypin[14]
  PIN dummypin[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 10.920 432.000 11.520 ;
    END
  END dummypin[15]
  PIN dummypin[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 369.280 432.000 369.880 ;
    END
  END dummypin[1]
  PIN dummypin[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 348.200 432.000 348.800 ;
    END
  END dummypin[2]
  PIN dummypin[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 327.120 432.000 327.720 ;
    END
  END dummypin[3]
  PIN dummypin[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 306.040 432.000 306.640 ;
    END
  END dummypin[4]
  PIN dummypin[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 284.960 432.000 285.560 ;
    END
  END dummypin[5]
  PIN dummypin[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 263.880 432.000 264.480 ;
    END
  END dummypin[6]
  PIN dummypin[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 242.800 432.000 243.400 ;
    END
  END dummypin[7]
  PIN dummypin[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 158.480 432.000 159.080 ;
    END
  END dummypin[8]
  PIN dummypin[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 137.400 432.000 138.000 ;
    END
  END dummypin[9]
  PIN inn_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 200.640 432.000 201.240 ;
    END
  END inn_analog
  PIN inp_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.000 221.720 432.000 222.320 ;
    END
  END inp_analog
  PIN result_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END result_out[0]
  PIN result_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END result_out[10]
  PIN result_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END result_out[11]
  PIN result_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END result_out[12]
  PIN result_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END result_out[13]
  PIN result_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END result_out[14]
  PIN result_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END result_out[15]
  PIN result_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END result_out[1]
  PIN result_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END result_out[2]
  PIN result_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END result_out[3]
  PIN result_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END result_out[4]
  PIN result_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END result_out[5]
  PIN result_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END result_out[6]
  PIN result_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END result_out[7]
  PIN result_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END result_out[8]
  PIN result_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END result_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END rst_n
  PIN start_conversion_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END start_conversion_in
  OBS
      LAYER li1 ;
        RECT 5.520 10.000 426.420 391.765 ;
      LAYER met1 ;
        RECT 3.290 5.820 427.270 391.920 ;
      LAYER met2 ;
        RECT 3.320 5.790 427.250 392.205 ;
      LAYER met3 ;
        RECT 4.400 391.360 428.000 392.185 ;
        RECT 4.400 391.320 427.600 391.360 ;
        RECT 4.000 389.960 427.600 391.320 ;
        RECT 4.000 385.240 428.000 389.960 ;
        RECT 4.400 383.840 428.000 385.240 ;
        RECT 4.000 377.760 428.000 383.840 ;
        RECT 4.400 376.360 428.000 377.760 ;
        RECT 4.000 370.280 428.000 376.360 ;
        RECT 4.400 368.880 427.600 370.280 ;
        RECT 4.000 362.800 428.000 368.880 ;
        RECT 4.400 361.400 428.000 362.800 ;
        RECT 4.000 355.320 428.000 361.400 ;
        RECT 4.400 353.920 428.000 355.320 ;
        RECT 4.000 349.200 428.000 353.920 ;
        RECT 4.000 347.840 427.600 349.200 ;
        RECT 4.400 347.800 427.600 347.840 ;
        RECT 4.400 346.440 428.000 347.800 ;
        RECT 4.000 340.360 428.000 346.440 ;
        RECT 4.400 338.960 428.000 340.360 ;
        RECT 4.000 332.880 428.000 338.960 ;
        RECT 4.400 331.480 428.000 332.880 ;
        RECT 4.000 328.120 428.000 331.480 ;
        RECT 4.000 326.720 427.600 328.120 ;
        RECT 4.000 325.400 428.000 326.720 ;
        RECT 4.400 324.000 428.000 325.400 ;
        RECT 4.000 317.920 428.000 324.000 ;
        RECT 4.400 316.520 428.000 317.920 ;
        RECT 4.000 310.440 428.000 316.520 ;
        RECT 4.400 309.040 428.000 310.440 ;
        RECT 4.000 307.040 428.000 309.040 ;
        RECT 4.000 305.640 427.600 307.040 ;
        RECT 4.000 302.960 428.000 305.640 ;
        RECT 4.400 301.560 428.000 302.960 ;
        RECT 4.000 295.480 428.000 301.560 ;
        RECT 4.400 294.080 428.000 295.480 ;
        RECT 4.000 288.000 428.000 294.080 ;
        RECT 4.400 286.600 428.000 288.000 ;
        RECT 4.000 285.960 428.000 286.600 ;
        RECT 4.000 284.560 427.600 285.960 ;
        RECT 4.000 280.520 428.000 284.560 ;
        RECT 4.400 279.120 428.000 280.520 ;
        RECT 4.000 273.040 428.000 279.120 ;
        RECT 4.400 271.640 428.000 273.040 ;
        RECT 4.000 265.560 428.000 271.640 ;
        RECT 4.400 264.880 428.000 265.560 ;
        RECT 4.400 264.160 427.600 264.880 ;
        RECT 4.000 263.480 427.600 264.160 ;
        RECT 4.000 258.080 428.000 263.480 ;
        RECT 4.400 256.680 428.000 258.080 ;
        RECT 4.000 250.600 428.000 256.680 ;
        RECT 4.400 249.200 428.000 250.600 ;
        RECT 4.000 243.800 428.000 249.200 ;
        RECT 4.000 243.120 427.600 243.800 ;
        RECT 4.400 242.400 427.600 243.120 ;
        RECT 4.400 241.720 428.000 242.400 ;
        RECT 4.000 235.640 428.000 241.720 ;
        RECT 4.400 234.240 428.000 235.640 ;
        RECT 4.000 228.160 428.000 234.240 ;
        RECT 4.400 226.760 428.000 228.160 ;
        RECT 4.000 222.720 428.000 226.760 ;
        RECT 4.000 221.320 427.600 222.720 ;
        RECT 4.000 220.680 428.000 221.320 ;
        RECT 4.400 219.280 428.000 220.680 ;
        RECT 4.000 213.200 428.000 219.280 ;
        RECT 4.400 211.800 428.000 213.200 ;
        RECT 4.000 205.720 428.000 211.800 ;
        RECT 4.400 204.320 428.000 205.720 ;
        RECT 4.000 201.640 428.000 204.320 ;
        RECT 4.000 200.240 427.600 201.640 ;
        RECT 4.000 198.240 428.000 200.240 ;
        RECT 4.400 196.840 428.000 198.240 ;
        RECT 4.000 190.760 428.000 196.840 ;
        RECT 4.400 189.360 428.000 190.760 ;
        RECT 4.000 183.280 428.000 189.360 ;
        RECT 4.400 181.880 428.000 183.280 ;
        RECT 4.000 180.560 428.000 181.880 ;
        RECT 4.000 179.160 427.600 180.560 ;
        RECT 4.000 175.800 428.000 179.160 ;
        RECT 4.400 174.400 428.000 175.800 ;
        RECT 4.000 168.320 428.000 174.400 ;
        RECT 4.400 166.920 428.000 168.320 ;
        RECT 4.000 160.840 428.000 166.920 ;
        RECT 4.400 159.480 428.000 160.840 ;
        RECT 4.400 159.440 427.600 159.480 ;
        RECT 4.000 158.080 427.600 159.440 ;
        RECT 4.000 153.360 428.000 158.080 ;
        RECT 4.400 151.960 428.000 153.360 ;
        RECT 4.000 145.880 428.000 151.960 ;
        RECT 4.400 144.480 428.000 145.880 ;
        RECT 4.000 138.400 428.000 144.480 ;
        RECT 4.400 137.000 427.600 138.400 ;
        RECT 4.000 130.920 428.000 137.000 ;
        RECT 4.400 129.520 428.000 130.920 ;
        RECT 4.000 123.440 428.000 129.520 ;
        RECT 4.400 122.040 428.000 123.440 ;
        RECT 4.000 117.320 428.000 122.040 ;
        RECT 4.000 115.960 427.600 117.320 ;
        RECT 4.400 115.920 427.600 115.960 ;
        RECT 4.400 114.560 428.000 115.920 ;
        RECT 4.000 108.480 428.000 114.560 ;
        RECT 4.400 107.080 428.000 108.480 ;
        RECT 4.000 101.000 428.000 107.080 ;
        RECT 4.400 99.600 428.000 101.000 ;
        RECT 4.000 96.240 428.000 99.600 ;
        RECT 4.000 94.840 427.600 96.240 ;
        RECT 4.000 93.520 428.000 94.840 ;
        RECT 4.400 92.120 428.000 93.520 ;
        RECT 4.000 86.040 428.000 92.120 ;
        RECT 4.400 84.640 428.000 86.040 ;
        RECT 4.000 78.560 428.000 84.640 ;
        RECT 4.400 77.160 428.000 78.560 ;
        RECT 4.000 75.160 428.000 77.160 ;
        RECT 4.000 73.760 427.600 75.160 ;
        RECT 4.000 71.080 428.000 73.760 ;
        RECT 4.400 69.680 428.000 71.080 ;
        RECT 4.000 63.600 428.000 69.680 ;
        RECT 4.400 62.200 428.000 63.600 ;
        RECT 4.000 56.120 428.000 62.200 ;
        RECT 4.400 54.720 428.000 56.120 ;
        RECT 4.000 54.080 428.000 54.720 ;
        RECT 4.000 52.680 427.600 54.080 ;
        RECT 4.000 48.640 428.000 52.680 ;
        RECT 4.400 47.240 428.000 48.640 ;
        RECT 4.000 41.160 428.000 47.240 ;
        RECT 4.400 39.760 428.000 41.160 ;
        RECT 4.000 33.680 428.000 39.760 ;
        RECT 4.400 33.000 428.000 33.680 ;
        RECT 4.400 32.280 427.600 33.000 ;
        RECT 4.000 31.600 427.600 32.280 ;
        RECT 4.000 26.200 428.000 31.600 ;
        RECT 4.400 24.800 428.000 26.200 ;
        RECT 4.000 18.720 428.000 24.800 ;
        RECT 4.400 17.320 428.000 18.720 ;
        RECT 4.000 11.920 428.000 17.320 ;
        RECT 4.000 11.240 427.600 11.920 ;
        RECT 4.400 10.520 427.600 11.240 ;
        RECT 4.400 10.000 428.000 10.520 ;
      LAYER met4 ;
        RECT 9.495 10.000 16.320 390.840 ;
        RECT 18.720 10.000 19.620 390.840 ;
        RECT 22.020 10.000 40.320 390.840 ;
        RECT 42.720 10.000 43.620 390.840 ;
        RECT 46.020 224.445 64.320 390.840 ;
        RECT 66.720 224.445 67.620 390.840 ;
        RECT 70.020 267.930 407.850 390.840 ;
        RECT 70.020 224.445 88.320 267.930 ;
        RECT 90.720 228.260 91.620 267.930 ;
        RECT 94.020 228.260 112.320 267.930 ;
        RECT 90.720 224.445 112.320 228.260 ;
        RECT 46.020 177.515 112.320 224.445 ;
        RECT 46.020 10.000 64.320 177.515 ;
        RECT 66.720 10.000 67.620 177.515 ;
        RECT 70.020 132.910 88.320 177.515 ;
        RECT 90.720 167.580 112.320 177.515 ;
        RECT 90.720 132.910 91.620 167.580 ;
        RECT 94.020 132.910 112.320 167.580 ;
        RECT 114.720 228.260 115.620 267.930 ;
        RECT 118.020 228.260 136.320 267.930 ;
        RECT 138.720 228.260 139.620 267.930 ;
        RECT 114.720 167.580 139.620 228.260 ;
        RECT 114.720 132.910 115.620 167.580 ;
        RECT 118.020 132.910 136.320 167.580 ;
        RECT 138.720 132.910 139.620 167.580 ;
        RECT 142.020 228.260 160.320 267.930 ;
        RECT 162.720 228.260 163.620 267.930 ;
        RECT 142.020 167.580 163.620 228.260 ;
        RECT 142.020 132.910 160.320 167.580 ;
        RECT 162.720 132.910 163.620 167.580 ;
        RECT 166.020 132.910 184.320 267.930 ;
        RECT 186.720 132.910 187.620 267.930 ;
        RECT 190.020 132.910 208.320 267.930 ;
        RECT 210.720 132.910 211.620 267.930 ;
        RECT 214.020 132.910 232.320 267.930 ;
        RECT 234.720 132.910 235.620 267.930 ;
        RECT 238.020 215.880 256.320 267.930 ;
        RECT 258.720 215.880 259.620 267.930 ;
        RECT 238.020 214.790 259.620 215.880 ;
        RECT 262.020 214.790 280.320 267.930 ;
        RECT 282.720 215.880 283.620 267.930 ;
        RECT 286.020 227.100 407.850 267.930 ;
        RECT 286.020 215.880 304.320 227.100 ;
        RECT 282.720 214.790 304.320 215.880 ;
        RECT 238.020 195.560 304.320 214.790 ;
        RECT 306.720 195.560 307.620 227.100 ;
        RECT 310.020 195.560 328.320 227.100 ;
        RECT 330.720 195.560 331.620 227.100 ;
        RECT 334.020 195.560 352.320 227.100 ;
        RECT 354.720 195.560 355.620 227.100 ;
        RECT 358.020 195.560 376.320 227.100 ;
        RECT 238.020 183.140 376.320 195.560 ;
        RECT 238.020 182.100 259.620 183.140 ;
        RECT 238.020 132.910 256.320 182.100 ;
        RECT 258.720 132.910 259.620 182.100 ;
        RECT 262.020 132.910 280.320 183.140 ;
        RECT 282.720 182.100 376.320 183.140 ;
        RECT 282.720 132.910 283.620 182.100 ;
        RECT 286.020 172.900 376.320 182.100 ;
        RECT 378.720 172.900 379.620 227.100 ;
        RECT 382.020 172.900 400.320 227.100 ;
        RECT 402.720 172.900 407.850 227.100 ;
        RECT 286.020 132.910 407.850 172.900 ;
        RECT 70.020 10.000 407.850 132.910 ;
      LAYER met5 ;
        RECT 94.400 256.580 254.960 364.890 ;
        RECT 94.400 232.580 254.960 248.480 ;
        RECT 94.400 208.580 254.960 224.480 ;
        RECT 94.400 184.580 254.960 200.480 ;
        RECT 94.400 160.580 254.960 176.480 ;
        RECT 94.400 136.580 254.960 152.480 ;
        RECT 94.400 35.950 254.960 131.780 ;
        RECT 265.680 69.690 298.440 78.350 ;
        RECT 265.730 288.235 298.460 296.560 ;
  END
END adc_top
END LIBRARY

