VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_array_matrix_12bit
  CLASS BLOCK ;
  FOREIGN adc_array_matrix_12bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 214.050 BY 120.840 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2.850 0.210 4.920 120.830 ;
    END
    PORT
      LAYER met4 ;
        RECT 182.700 0.860 184.770 99.510 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.540 0.830 211.610 120.830 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 5.230 0.210 7.300 120.830 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.320 0.860 182.390 99.510 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.980 0.840 214.050 120.840 ;
    END
  END VSS
  PIN vcm
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.210 0.000 186.820 5.745 ;
    END
  END vcm
  PIN sample
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.450 0.000 1.790 11.340 ;
    END
  END sample
  PIN sample_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.910 0.000 1.250 13.180 ;
    END
  END sample_n
  PIN row_n[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 87.040 9.470 87.180 ;
    END
  END row_n[15]
  PIN row_n[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 82.020 9.470 82.160 ;
    END
  END row_n[14]
  PIN row_n[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 77.000 9.470 77.140 ;
    END
  END row_n[13]
  PIN row_n[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 71.980 9.470 72.120 ;
    END
  END row_n[12]
  PIN row_n[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 66.960 9.470 67.100 ;
    END
  END row_n[11]
  PIN row_n[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 61.940 9.470 62.080 ;
    END
  END row_n[10]
  PIN row_n[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 56.920 9.470 57.060 ;
    END
  END row_n[9]
  PIN row_n[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 51.900 9.470 52.040 ;
    END
  END row_n[8]
  PIN row_n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 46.880 9.470 47.020 ;
    END
  END row_n[7]
  PIN row_n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 41.860 9.470 42.000 ;
    END
  END row_n[6]
  PIN row_n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 36.840 9.470 36.980 ;
    END
  END row_n[5]
  PIN row_n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 31.820 9.470 31.960 ;
    END
  END row_n[4]
  PIN row_n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 26.800 9.470 26.940 ;
    END
  END row_n[3]
  PIN row_n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 21.780 9.470 21.920 ;
    END
  END row_n[2]
  PIN row_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 16.760 9.470 16.900 ;
    END
  END row_n[1]
  PIN row_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 11.740 9.470 11.880 ;
    END
  END row_n[0]
  PIN rowon_n[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 87.450 16.070 87.590 ;
    END
  END rowon_n[15]
  PIN rowon_n[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 82.430 16.070 82.570 ;
    END
  END rowon_n[14]
  PIN rowon_n[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 77.410 16.070 77.550 ;
    END
  END rowon_n[13]
  PIN rowon_n[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 72.390 16.070 72.530 ;
    END
  END rowon_n[12]
  PIN rowon_n[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 67.370 16.070 67.510 ;
    END
  END rowon_n[11]
  PIN rowon_n[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 62.350 16.070 62.490 ;
    END
  END rowon_n[10]
  PIN rowon_n[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 57.330 16.070 57.470 ;
    END
  END rowon_n[9]
  PIN rowon_n[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 52.310 16.070 52.450 ;
    END
  END rowon_n[8]
  PIN rowon_n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 47.290 16.070 47.430 ;
    END
  END rowon_n[7]
  PIN rowon_n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 42.270 16.070 42.410 ;
    END
  END rowon_n[6]
  PIN rowon_n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 37.250 16.070 37.390 ;
    END
  END rowon_n[5]
  PIN rowon_n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 32.230 16.070 32.370 ;
    END
  END rowon_n[4]
  PIN rowon_n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 27.210 16.070 27.350 ;
    END
  END rowon_n[3]
  PIN rowon_n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 22.190 16.070 22.330 ;
    END
  END rowon_n[2]
  PIN rowon_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 17.170 16.070 17.310 ;
    END
  END rowon_n[1]
  PIN rowon_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 12.150 16.070 12.290 ;
    END
  END rowon_n[0]
  PIN col_n[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.410 0.000 145.580 1.445 ;
    END
  END col_n[31]
  PIN col_n[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 0.000 144.560 1.825 ;
    END
  END col_n[30]
  PIN col_n[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.370 0.000 143.540 2.205 ;
    END
  END col_n[29]
  PIN col_n[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.350 0.000 142.520 2.590 ;
    END
  END col_n[28]
  PIN col_n[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.330 0.000 141.500 2.985 ;
    END
  END col_n[27]
  PIN col_n[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.310 0.000 140.480 3.335 ;
    END
  END col_n[26]
  PIN col_n[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.290 0.000 139.460 3.715 ;
    END
  END col_n[25]
  PIN col_n[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.270 0.000 138.440 4.290 ;
    END
  END col_n[24]
  PIN col_n[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.250 0.000 133.420 4.290 ;
    END
  END col_n[23]
  PIN col_n[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.230 0.000 128.400 4.290 ;
    END
  END col_n[22]
  PIN col_n[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.210 0.000 123.380 4.290 ;
    END
  END col_n[21]
  PIN col_n[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.190 0.000 118.360 4.290 ;
    END
  END col_n[20]
  PIN col_n[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.170 0.000 113.340 4.290 ;
    END
  END col_n[19]
  PIN col_n[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.150 0.000 108.320 4.290 ;
    END
  END col_n[18]
  PIN col_n[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.300 4.290 ;
    END
  END col_n[17]
  PIN col_n[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.110 0.000 98.280 4.290 ;
    END
  END col_n[16]
  PIN col_n[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.090 0.000 93.260 4.290 ;
    END
  END col_n[15]
  PIN col_n[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.070 0.000 88.240 4.290 ;
    END
  END col_n[14]
  PIN col_n[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.050 0.000 83.220 4.290 ;
    END
  END col_n[13]
  PIN col_n[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.030 0.000 78.200 4.290 ;
    END
  END col_n[12]
  PIN col_n[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.010 0.000 73.180 4.290 ;
    END
  END col_n[11]
  PIN col_n[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.990 0.000 68.160 4.290 ;
    END
  END col_n[10]
  PIN col_n[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.970 0.000 63.140 4.290 ;
    END
  END col_n[9]
  PIN col_n[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.950 0.000 58.120 4.290 ;
    END
  END col_n[8]
  PIN col_n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.930 0.000 53.100 4.290 ;
    END
  END col_n[7]
  PIN col_n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.910 0.000 48.080 4.290 ;
    END
  END col_n[6]
  PIN col_n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.890 0.000 43.060 4.290 ;
    END
  END col_n[5]
  PIN col_n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.870 0.000 38.040 4.290 ;
    END
  END col_n[4]
  PIN col_n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.850 0.000 33.020 4.290 ;
    END
  END col_n[3]
  PIN col_n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.830 0.000 28.000 4.290 ;
    END
  END col_n[2]
  PIN col_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.810 0.000 22.980 4.290 ;
    END
  END col_n[1]
  PIN col_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.790 0.000 17.960 4.285 ;
    END
  END col_n[0]
  PIN en_bit_n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.450 0.000 96.620 4.295 ;
    END
  END en_bit_n[2]
  PIN en_bit_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.430 0.000 91.600 4.295 ;
    END
  END en_bit_n[1]
  PIN en_bit_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.470 0.000 101.640 4.295 ;
    END
  END en_bit_n[0]
  PIN en_C0_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.150 0.000 21.320 4.295 ;
    END
  END en_C0_n
  PIN sw
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.900 0.000 171.095 7.005 ;
    END
  END sw
  PIN sw_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.770 0.000 172.965 7.010 ;
    END
  END sw_n
  PIN analog_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 170.705 0.040 214.050 0.620 ;
    END
  END analog_in
  PIN ctop
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 171.500 0.000 171.800 10.490 ;
    END
  END ctop
  OBS
      LAYER li1 ;
        RECT 5.230 0.830 213.300 120.830 ;
      LAYER met1 ;
        RECT 0.000 87.870 213.300 120.830 ;
        RECT 16.350 87.170 213.300 87.870 ;
        RECT 9.750 86.760 213.300 87.170 ;
        RECT 0.000 82.850 213.300 86.760 ;
        RECT 16.350 82.150 213.300 82.850 ;
        RECT 9.750 81.740 213.300 82.150 ;
        RECT 0.000 77.830 213.300 81.740 ;
        RECT 16.350 77.130 213.300 77.830 ;
        RECT 9.750 76.720 213.300 77.130 ;
        RECT 0.000 72.810 213.300 76.720 ;
        RECT 16.350 72.110 213.300 72.810 ;
        RECT 9.750 71.700 213.300 72.110 ;
        RECT 0.000 67.790 213.300 71.700 ;
        RECT 16.350 67.090 213.300 67.790 ;
        RECT 9.750 66.680 213.300 67.090 ;
        RECT 0.000 62.770 213.300 66.680 ;
        RECT 16.350 62.070 213.300 62.770 ;
        RECT 9.750 61.660 213.300 62.070 ;
        RECT 0.000 57.750 213.300 61.660 ;
        RECT 16.350 57.050 213.300 57.750 ;
        RECT 9.750 56.640 213.300 57.050 ;
        RECT 0.000 52.730 213.300 56.640 ;
        RECT 16.350 52.030 213.300 52.730 ;
        RECT 9.750 51.620 213.300 52.030 ;
        RECT 0.000 47.710 213.300 51.620 ;
        RECT 16.350 47.010 213.300 47.710 ;
        RECT 9.750 46.600 213.300 47.010 ;
        RECT 0.000 42.690 213.300 46.600 ;
        RECT 16.350 41.990 213.300 42.690 ;
        RECT 9.750 41.580 213.300 41.990 ;
        RECT 0.000 37.670 213.300 41.580 ;
        RECT 16.350 36.970 213.300 37.670 ;
        RECT 9.750 36.560 213.300 36.970 ;
        RECT 0.000 32.650 213.300 36.560 ;
        RECT 16.350 31.950 213.300 32.650 ;
        RECT 9.750 31.540 213.300 31.950 ;
        RECT 0.000 27.630 213.300 31.540 ;
        RECT 16.350 26.930 213.300 27.630 ;
        RECT 9.750 26.520 213.300 26.930 ;
        RECT 0.000 22.610 213.300 26.520 ;
        RECT 16.350 21.910 213.300 22.610 ;
        RECT 9.750 21.500 213.300 21.910 ;
        RECT 0.000 17.590 213.300 21.500 ;
        RECT 16.350 16.890 213.300 17.590 ;
        RECT 9.750 16.480 213.300 16.890 ;
        RECT 0.000 12.570 213.300 16.480 ;
        RECT 16.350 11.870 213.300 12.570 ;
        RECT 9.750 11.460 213.300 11.870 ;
        RECT 0.000 0.900 213.300 11.460 ;
        RECT 0.000 0.040 170.425 0.900 ;
      LAYER met2 ;
        RECT 0.910 13.460 213.300 120.830 ;
        RECT 1.530 11.620 213.300 13.460 ;
        RECT 2.070 7.290 213.300 11.620 ;
        RECT 2.070 7.285 172.490 7.290 ;
        RECT 2.070 4.575 170.620 7.285 ;
        RECT 2.070 4.565 20.870 4.575 ;
        RECT 2.070 0.000 17.510 4.565 ;
        RECT 18.240 0.000 20.870 4.565 ;
        RECT 21.600 4.570 91.150 4.575 ;
        RECT 21.600 0.000 22.530 4.570 ;
        RECT 23.260 0.000 27.550 4.570 ;
        RECT 28.280 0.000 32.570 4.570 ;
        RECT 33.300 0.000 37.590 4.570 ;
        RECT 38.320 0.000 42.610 4.570 ;
        RECT 43.340 0.000 47.630 4.570 ;
        RECT 48.360 0.000 52.650 4.570 ;
        RECT 53.380 0.000 57.670 4.570 ;
        RECT 58.400 0.000 62.690 4.570 ;
        RECT 63.420 0.000 67.710 4.570 ;
        RECT 68.440 0.000 72.730 4.570 ;
        RECT 73.460 0.000 77.750 4.570 ;
        RECT 78.480 0.000 82.770 4.570 ;
        RECT 83.500 0.000 87.790 4.570 ;
        RECT 88.520 0.000 91.150 4.570 ;
        RECT 91.880 4.570 96.170 4.575 ;
        RECT 91.880 0.000 92.810 4.570 ;
        RECT 93.540 0.000 96.170 4.570 ;
        RECT 96.900 4.570 101.190 4.575 ;
        RECT 96.900 0.000 97.830 4.570 ;
        RECT 98.560 0.000 101.190 4.570 ;
        RECT 101.920 4.570 170.620 4.575 ;
        RECT 101.920 0.000 102.850 4.570 ;
        RECT 103.580 0.000 107.870 4.570 ;
        RECT 108.600 0.000 112.890 4.570 ;
        RECT 113.620 0.000 117.910 4.570 ;
        RECT 118.640 0.000 122.930 4.570 ;
        RECT 123.660 0.000 127.950 4.570 ;
        RECT 128.680 0.000 132.970 4.570 ;
        RECT 133.700 0.000 137.990 4.570 ;
        RECT 138.720 3.995 170.620 4.570 ;
        RECT 138.720 0.000 139.010 3.995 ;
        RECT 139.740 3.615 170.620 3.995 ;
        RECT 139.740 0.000 140.030 3.615 ;
        RECT 140.760 3.265 170.620 3.615 ;
        RECT 140.760 0.000 141.050 3.265 ;
        RECT 141.780 2.870 170.620 3.265 ;
        RECT 141.780 0.000 142.070 2.870 ;
        RECT 142.800 2.485 170.620 2.870 ;
        RECT 142.800 0.000 143.090 2.485 ;
        RECT 143.820 2.105 170.620 2.485 ;
        RECT 143.820 0.000 144.110 2.105 ;
        RECT 144.840 1.725 170.620 2.105 ;
        RECT 144.840 0.000 145.130 1.725 ;
        RECT 145.860 0.000 170.620 1.725 ;
        RECT 171.375 0.000 172.490 7.285 ;
        RECT 173.245 6.025 213.300 7.290 ;
        RECT 173.245 0.000 184.930 6.025 ;
        RECT 187.100 0.000 213.300 6.025 ;
      LAYER met3 ;
        RECT 2.850 0.830 213.300 120.830 ;
      LAYER met4 ;
        RECT 8.010 99.910 209.140 120.830 ;
        RECT 8.010 10.890 179.920 99.910 ;
        RECT 8.010 0.830 171.100 10.890 ;
        RECT 172.200 0.830 179.920 10.890 ;
        RECT 185.170 0.830 209.140 99.910 ;
  END
END adc_array_matrix_12bit
END LIBRARY

