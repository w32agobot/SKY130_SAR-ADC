* NGSPICE file created from sky130_mm_sc_hd_dly5ns.ext - technology: sky130A

.subckt sky130_mm_sc_hd_dly5ns_postlayout VPWR in out VGND VPB VNB 
X0 cap_top VGND sky130_fd_pr__cap_mim_m3_1 l=1.93e+06u w=3.695e+06u
X1 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=2.478e+11p ps=2.86e+06u w=420000u l=4e+06u
X2 a_1154_296# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X3 out cap_top a_1154_296# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X4 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=4e+06u
X5 cap_top VGND sky130_fd_pr__cap_mim_m3_1 l=1.93e+06u w=2.38e+06u
X6 out cap_top a_1176_80# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X7 a_1176_80# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1176_80# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 VGND out a_1154_296# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10 a_1154_296# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11 VPWR out a_1176_80# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

