** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_matrix_12bit.sch
.subckt adc_array_matrix_12bit VDD VSS vcm sample sample_n row_n[0] row_n[1] row_n[2] row_n[3]
+ row_n[4] row_n[5] row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12] row_n[13] row_n[14]
+ row_n[15] rowon_n[0] rowon_n[1] rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6] rowon_n[7] rowon_n[8]
+ rowon_n[9] rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13] rowon_n[14] rowon_n[15] col_n[0] col_n[1] col_n[2]
+ col_n[3] col_n[4] col_n[5] col_n[6] col_n[7] col_n[8] col_n[9] col_n[10] col_n[11] col_n[12] col_n[13]
+ col_n[14] col_n[15] col_n[16] col_n[17] col_n[18] col_n[19] col_n[20] col_n[21] col_n[22] col_n[23] col_n[24]
+ col_n[25] col_n[26] col_n[27] col_n[28] col_n[29] col_n[30] col_n[31] en_bit_n[0] en_bit_n[1] en_bit_n[2]
+ en_C0_n sw sw_n analog_in ctop
*.PININFO VDD:B VSS:B vcm:B sample:I sample_n:I row_n[0:15]:I rowon_n[0:15]:I col_n[0:31]:I
*+ en_bit_n[0:2]:I en_C0_n:I sw:I sw_n:I analog_in:I ctop:B
x2 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[1] adc_array_wafflecap_8_8
x3 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[2] adc_array_wafflecap_8_8
x4 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[3] adc_array_wafflecap_8_8
x5 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[4] adc_array_wafflecap_8_8
x6 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[5] adc_array_wafflecap_8_8
x7 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[6] adc_array_wafflecap_8_8
x8 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[7] adc_array_wafflecap_8_8
x9 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[8] adc_array_wafflecap_8_8
x10 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[9] adc_array_wafflecap_8_8
x11 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[10] adc_array_wafflecap_8_8
x12 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[11] adc_array_wafflecap_8_8
x13 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[12] adc_array_wafflecap_8_8
x15 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[14] adc_array_wafflecap_8_8
x16 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[15] adc_array_wafflecap_8_8
x17 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[16] adc_array_wafflecap_8_8
x18 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[17] adc_array_wafflecap_8_8
x19 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[18] adc_array_wafflecap_8_8
x20 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[19] adc_array_wafflecap_8_8
x21 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[20] adc_array_wafflecap_8_8
x22 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[21] adc_array_wafflecap_8_8
x23 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[22] adc_array_wafflecap_8_8
x24 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[23] adc_array_wafflecap_8_8
x25 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[24] adc_array_wafflecap_8_8
x26 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[25] adc_array_wafflecap_8_8
x27 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[26] adc_array_wafflecap_8_8
x28 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[27] adc_array_wafflecap_8_8
x29 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[28] adc_array_wafflecap_8_8
x30 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[29] adc_array_wafflecap_8_8
x31 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[30] adc_array_wafflecap_8_8
x32 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[31] adc_array_wafflecap_8_8
x33 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[0] adc_array_wafflecap_8_8
x34 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[1] adc_array_wafflecap_8_8
x35 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[2] adc_array_wafflecap_8_8
x36 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[3] adc_array_wafflecap_8_8
x37 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[4] adc_array_wafflecap_8_8
x38 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[5] adc_array_wafflecap_8_8
x39 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[6] adc_array_wafflecap_8_8
x40 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[7] adc_array_wafflecap_8_8
x41 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[8] adc_array_wafflecap_8_8
x42 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[9] adc_array_wafflecap_8_8
x43 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[10] adc_array_wafflecap_8_8
x44 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[11] adc_array_wafflecap_8_8
x45 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[12] adc_array_wafflecap_8_8
x46 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[13] adc_array_wafflecap_8_8
x47 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[14] adc_array_wafflecap_8_8
x48 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[15] adc_array_wafflecap_8_8
x49 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[16] adc_array_wafflecap_8_8
x50 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[17] adc_array_wafflecap_8_8
x51 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[18] adc_array_wafflecap_8_8
x52 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[19] adc_array_wafflecap_8_8
x53 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[20] adc_array_wafflecap_8_8
x54 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[21] adc_array_wafflecap_8_8
x55 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[22] adc_array_wafflecap_8_8
x56 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[23] adc_array_wafflecap_8_8
x57 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[24] adc_array_wafflecap_8_8
x58 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[25] adc_array_wafflecap_8_8
x59 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[26] adc_array_wafflecap_8_8
x60 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[27] adc_array_wafflecap_8_8
x61 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[28] adc_array_wafflecap_8_8
x62 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[29] adc_array_wafflecap_8_8
x63 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[30] adc_array_wafflecap_8_8
x64 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS col_n[31] adc_array_wafflecap_8_8
x65 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[0] adc_array_wafflecap_8_8
x66 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[1] adc_array_wafflecap_8_8
x67 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[2] adc_array_wafflecap_8_8
x68 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[3] adc_array_wafflecap_8_8
x69 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[4] adc_array_wafflecap_8_8
x70 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[5] adc_array_wafflecap_8_8
x71 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[6] adc_array_wafflecap_8_8
x72 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[7] adc_array_wafflecap_8_8
x73 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[8] adc_array_wafflecap_8_8
x74 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[9] adc_array_wafflecap_8_8
x75 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[10] adc_array_wafflecap_8_8
x76 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[11] adc_array_wafflecap_8_8
x77 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[12] adc_array_wafflecap_8_8
x78 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[13] adc_array_wafflecap_8_8
x79 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[14] adc_array_wafflecap_8_8
x80 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[15] adc_array_wafflecap_8_8
x81 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[16] adc_array_wafflecap_8_8
x82 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[17] adc_array_wafflecap_8_8
x83 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[18] adc_array_wafflecap_8_8
x84 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[19] adc_array_wafflecap_8_8
x85 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[20] adc_array_wafflecap_8_8
x86 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[21] adc_array_wafflecap_8_8
x87 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[22] adc_array_wafflecap_8_8
x88 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[23] adc_array_wafflecap_8_8
x89 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[24] adc_array_wafflecap_8_8
x90 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[25] adc_array_wafflecap_8_8
x91 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[26] adc_array_wafflecap_8_8
x92 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[27] adc_array_wafflecap_8_8
x93 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[28] adc_array_wafflecap_8_8
x94 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[29] adc_array_wafflecap_8_8
x95 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[30] adc_array_wafflecap_8_8
x96 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS col_n[31] adc_array_wafflecap_8_8
x97 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[0] adc_array_wafflecap_8_8
x98 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[1] adc_array_wafflecap_8_8
x99 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[2] adc_array_wafflecap_8_8
x100 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[3] adc_array_wafflecap_8_8
x101 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[4] adc_array_wafflecap_8_8
x102 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[5] adc_array_wafflecap_8_8
x103 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[6] adc_array_wafflecap_8_8
x104 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[7] adc_array_wafflecap_8_8
x105 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[8] adc_array_wafflecap_8_8
x106 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[9] adc_array_wafflecap_8_8
x107 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[10] adc_array_wafflecap_8_8
x108 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[11] adc_array_wafflecap_8_8
x109 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[12] adc_array_wafflecap_8_8
x110 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[13] adc_array_wafflecap_8_8
x111 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[14] adc_array_wafflecap_8_8
x112 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[15] adc_array_wafflecap_8_8
x113 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[16] adc_array_wafflecap_8_8
x114 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[17] adc_array_wafflecap_8_8
x115 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[18] adc_array_wafflecap_8_8
x116 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[19] adc_array_wafflecap_8_8
x117 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[20] adc_array_wafflecap_8_8
x118 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[21] adc_array_wafflecap_8_8
x119 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[22] adc_array_wafflecap_8_8
x120 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[23] adc_array_wafflecap_8_8
x121 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[24] adc_array_wafflecap_8_8
x122 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[25] adc_array_wafflecap_8_8
x123 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[26] adc_array_wafflecap_8_8
x124 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[27] adc_array_wafflecap_8_8
x125 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[28] adc_array_wafflecap_8_8
x126 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[29] adc_array_wafflecap_8_8
x127 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[30] adc_array_wafflecap_8_8
x128 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS col_n[31] adc_array_wafflecap_8_8
x129 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[0] adc_array_wafflecap_8_8
x130 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[1] adc_array_wafflecap_8_8
x131 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[2] adc_array_wafflecap_8_8
x132 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[3] adc_array_wafflecap_8_8
x133 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[4] adc_array_wafflecap_8_8
x134 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[5] adc_array_wafflecap_8_8
x135 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[6] adc_array_wafflecap_8_8
x136 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[7] adc_array_wafflecap_8_8
x137 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[8] adc_array_wafflecap_8_8
x138 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[9] adc_array_wafflecap_8_8
x139 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[10] adc_array_wafflecap_8_8
x140 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[11] adc_array_wafflecap_8_8
x141 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[12] adc_array_wafflecap_8_8
x142 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[13] adc_array_wafflecap_8_8
x143 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[14] adc_array_wafflecap_8_8
x144 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[15] adc_array_wafflecap_8_8
x145 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[16] adc_array_wafflecap_8_8
x146 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[17] adc_array_wafflecap_8_8
x147 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[18] adc_array_wafflecap_8_8
x148 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[19] adc_array_wafflecap_8_8
x149 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[20] adc_array_wafflecap_8_8
x150 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[21] adc_array_wafflecap_8_8
x151 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[22] adc_array_wafflecap_8_8
x152 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[23] adc_array_wafflecap_8_8
x153 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[24] adc_array_wafflecap_8_8
x154 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[25] adc_array_wafflecap_8_8
x155 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[26] adc_array_wafflecap_8_8
x156 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[27] adc_array_wafflecap_8_8
x157 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[28] adc_array_wafflecap_8_8
x158 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[29] adc_array_wafflecap_8_8
x159 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[30] adc_array_wafflecap_8_8
x160 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS col_n[31] adc_array_wafflecap_8_8
x161 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[0] adc_array_wafflecap_8_8
x162 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[1] adc_array_wafflecap_8_8
x163 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[2] adc_array_wafflecap_8_8
x164 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[3] adc_array_wafflecap_8_8
x165 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[4] adc_array_wafflecap_8_8
x166 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[5] adc_array_wafflecap_8_8
x167 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[6] adc_array_wafflecap_8_8
x168 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[7] adc_array_wafflecap_8_8
x169 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[8] adc_array_wafflecap_8_8
x170 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[9] adc_array_wafflecap_8_8
x171 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[10] adc_array_wafflecap_8_8
x172 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[11] adc_array_wafflecap_8_8
x173 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[12] adc_array_wafflecap_8_8
x174 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[13] adc_array_wafflecap_8_8
x175 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[14] adc_array_wafflecap_8_8
x176 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[15] adc_array_wafflecap_8_8
x177 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[16] adc_array_wafflecap_8_8
x178 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[17] adc_array_wafflecap_8_8
x179 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[18] adc_array_wafflecap_8_8
x180 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[19] adc_array_wafflecap_8_8
x181 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[20] adc_array_wafflecap_8_8
x182 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[21] adc_array_wafflecap_8_8
x183 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[22] adc_array_wafflecap_8_8
x184 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[23] adc_array_wafflecap_8_8
x185 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[24] adc_array_wafflecap_8_8
x186 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[25] adc_array_wafflecap_8_8
x187 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[26] adc_array_wafflecap_8_8
x188 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[27] adc_array_wafflecap_8_8
x189 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[28] adc_array_wafflecap_8_8
x190 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[29] adc_array_wafflecap_8_8
x191 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[30] adc_array_wafflecap_8_8
x192 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS col_n[31] adc_array_wafflecap_8_8
x193 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[0] adc_array_wafflecap_8_8
x194 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[1] adc_array_wafflecap_8_8
x195 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[2] adc_array_wafflecap_8_8
x196 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[3] adc_array_wafflecap_8_8
x197 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[4] adc_array_wafflecap_8_8
x198 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[5] adc_array_wafflecap_8_8
x199 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[6] adc_array_wafflecap_8_8
x200 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[7] adc_array_wafflecap_8_8
x201 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[8] adc_array_wafflecap_8_8
x202 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[9] adc_array_wafflecap_8_8
x203 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[10] adc_array_wafflecap_8_8
x204 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[11] adc_array_wafflecap_8_8
x205 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[12] adc_array_wafflecap_8_8
x206 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[13] adc_array_wafflecap_8_8
x207 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[14] adc_array_wafflecap_8_8
x208 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[15] adc_array_wafflecap_8_8
x209 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[16] adc_array_wafflecap_8_8
x210 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[17] adc_array_wafflecap_8_8
x211 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[18] adc_array_wafflecap_8_8
x212 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[19] adc_array_wafflecap_8_8
x213 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[20] adc_array_wafflecap_8_8
x214 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[21] adc_array_wafflecap_8_8
x215 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[22] adc_array_wafflecap_8_8
x216 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[23] adc_array_wafflecap_8_8
x217 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[24] adc_array_wafflecap_8_8
x218 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[25] adc_array_wafflecap_8_8
x219 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[26] adc_array_wafflecap_8_8
x220 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[27] adc_array_wafflecap_8_8
x221 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[28] adc_array_wafflecap_8_8
x222 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[29] adc_array_wafflecap_8_8
x223 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[30] adc_array_wafflecap_8_8
x224 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS col_n[31] adc_array_wafflecap_8_8
x225 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[0] adc_array_wafflecap_8_8
x226 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[1] adc_array_wafflecap_8_8
x227 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[2] adc_array_wafflecap_8_8
x228 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[3] adc_array_wafflecap_8_8
x229 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[4] adc_array_wafflecap_8_8
x230 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[5] adc_array_wafflecap_8_8
x231 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[6] adc_array_wafflecap_8_8
x232 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[7] adc_array_wafflecap_8_8
x233 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[8] adc_array_wafflecap_8_8
x234 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[9] adc_array_wafflecap_8_8
x235 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[10] adc_array_wafflecap_8_8
x236 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[11] adc_array_wafflecap_8_8
x237 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[12] adc_array_wafflecap_8_8
x238 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[13] adc_array_wafflecap_8_8
x239 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[14] adc_array_wafflecap_8_8
x240 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[15] adc_array_wafflecap_8_8
x241 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[16] adc_array_wafflecap_8_8
x242 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[17] adc_array_wafflecap_8_8
x243 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[18] adc_array_wafflecap_8_8
x244 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[19] adc_array_wafflecap_8_8
x245 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[20] adc_array_wafflecap_8_8
x246 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[21] adc_array_wafflecap_8_8
x247 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[22] adc_array_wafflecap_8_8
x248 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[23] adc_array_wafflecap_8_8
x249 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[24] adc_array_wafflecap_8_8
x250 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[25] adc_array_wafflecap_8_8
x251 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[26] adc_array_wafflecap_8_8
x252 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[27] adc_array_wafflecap_8_8
x253 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[28] adc_array_wafflecap_8_8
x254 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[29] adc_array_wafflecap_8_8
x255 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[30] adc_array_wafflecap_8_8
x256 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS col_n[31] adc_array_wafflecap_8_8
x257 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[0] adc_array_wafflecap_8_8
x258 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[1] adc_array_wafflecap_8_8
x259 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[2] adc_array_wafflecap_8_8
x260 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[3] adc_array_wafflecap_8_8
x261 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[4] adc_array_wafflecap_8_8
x262 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[5] adc_array_wafflecap_8_8
x263 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[6] adc_array_wafflecap_8_8
x264 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[7] adc_array_wafflecap_8_8
x265 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[8] adc_array_wafflecap_8_8
x266 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[9] adc_array_wafflecap_8_8
x267 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[10] adc_array_wafflecap_8_8
x268 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[11] adc_array_wafflecap_8_8
x269 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[12] adc_array_wafflecap_8_8
x270 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[13] adc_array_wafflecap_8_8
x271 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[14] adc_array_wafflecap_8_8
x272 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[15] adc_array_wafflecap_8_8
x273 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[16] adc_array_wafflecap_8_8
x274 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[17] adc_array_wafflecap_8_8
x275 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[18] adc_array_wafflecap_8_8
x276 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[19] adc_array_wafflecap_8_8
x277 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[20] adc_array_wafflecap_8_8
x278 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[21] adc_array_wafflecap_8_8
x279 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[22] adc_array_wafflecap_8_8
x280 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[23] adc_array_wafflecap_8_8
x281 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[24] adc_array_wafflecap_8_8
x282 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[25] adc_array_wafflecap_8_8
x283 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[26] adc_array_wafflecap_8_8
x284 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[27] adc_array_wafflecap_8_8
x285 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[28] adc_array_wafflecap_8_8
x286 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[29] adc_array_wafflecap_8_8
x287 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[30] adc_array_wafflecap_8_8
x288 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS col_n[31] adc_array_wafflecap_8_8
x289 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[0] adc_array_wafflecap_8_8
x290 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[1] adc_array_wafflecap_8_8
x291 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[2] adc_array_wafflecap_8_8
x292 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[3] adc_array_wafflecap_8_8
x293 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[4] adc_array_wafflecap_8_8
x294 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[5] adc_array_wafflecap_8_8
x295 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[6] adc_array_wafflecap_8_8
x296 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[7] adc_array_wafflecap_8_8
x297 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[8] adc_array_wafflecap_8_8
x298 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[9] adc_array_wafflecap_8_8
x299 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[10] adc_array_wafflecap_8_8
x300 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[11] adc_array_wafflecap_8_8
x301 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[12] adc_array_wafflecap_8_8
x302 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[13] adc_array_wafflecap_8_8
x303 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[14] adc_array_wafflecap_8_8
x304 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[15] adc_array_wafflecap_8_8
x305 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[16] adc_array_wafflecap_8_8
x306 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[17] adc_array_wafflecap_8_8
x307 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[18] adc_array_wafflecap_8_8
x308 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[19] adc_array_wafflecap_8_8
x309 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[20] adc_array_wafflecap_8_8
x310 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[21] adc_array_wafflecap_8_8
x311 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[22] adc_array_wafflecap_8_8
x312 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[23] adc_array_wafflecap_8_8
x313 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[24] adc_array_wafflecap_8_8
x314 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[25] adc_array_wafflecap_8_8
x315 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[26] adc_array_wafflecap_8_8
x316 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[27] adc_array_wafflecap_8_8
x317 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[28] adc_array_wafflecap_8_8
x318 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[29] adc_array_wafflecap_8_8
x319 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[30] adc_array_wafflecap_8_8
x320 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS col_n[31] adc_array_wafflecap_8_8
x321 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[0] adc_array_wafflecap_8_8
x322 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[1] adc_array_wafflecap_8_8
x323 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[2] adc_array_wafflecap_8_8
x324 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[3] adc_array_wafflecap_8_8
x325 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[4] adc_array_wafflecap_8_8
x326 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[5] adc_array_wafflecap_8_8
x327 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[6] adc_array_wafflecap_8_8
x328 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[7] adc_array_wafflecap_8_8
x329 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[8] adc_array_wafflecap_8_8
x330 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[9] adc_array_wafflecap_8_8
x331 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[10] adc_array_wafflecap_8_8
x332 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[11] adc_array_wafflecap_8_8
x333 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[12] adc_array_wafflecap_8_8
x334 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[13] adc_array_wafflecap_8_8
x335 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[14] adc_array_wafflecap_8_8
x336 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[15] adc_array_wafflecap_8_8
x337 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[16] adc_array_wafflecap_8_8
x338 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[17] adc_array_wafflecap_8_8
x339 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[18] adc_array_wafflecap_8_8
x340 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[19] adc_array_wafflecap_8_8
x341 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[20] adc_array_wafflecap_8_8
x342 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[21] adc_array_wafflecap_8_8
x343 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[22] adc_array_wafflecap_8_8
x344 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[23] adc_array_wafflecap_8_8
x345 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[24] adc_array_wafflecap_8_8
x346 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[25] adc_array_wafflecap_8_8
x347 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[26] adc_array_wafflecap_8_8
x348 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[27] adc_array_wafflecap_8_8
x349 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[28] adc_array_wafflecap_8_8
x350 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[29] adc_array_wafflecap_8_8
x351 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[30] adc_array_wafflecap_8_8
x352 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS col_n[31] adc_array_wafflecap_8_8
x353 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[0] adc_array_wafflecap_8_8
x354 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[1] adc_array_wafflecap_8_8
x355 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[2] adc_array_wafflecap_8_8
x356 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[3] adc_array_wafflecap_8_8
x357 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[4] adc_array_wafflecap_8_8
x358 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[5] adc_array_wafflecap_8_8
x359 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[6] adc_array_wafflecap_8_8
x360 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[7] adc_array_wafflecap_8_8
x361 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[8] adc_array_wafflecap_8_8
x362 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[9] adc_array_wafflecap_8_8
x363 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[10] adc_array_wafflecap_8_8
x364 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[11] adc_array_wafflecap_8_8
x365 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[12] adc_array_wafflecap_8_8
x366 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[13] adc_array_wafflecap_8_8
x367 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[14] adc_array_wafflecap_8_8
x368 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[15] adc_array_wafflecap_8_8
x369 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[16] adc_array_wafflecap_8_8
x370 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[17] adc_array_wafflecap_8_8
x371 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[18] adc_array_wafflecap_8_8
x372 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[19] adc_array_wafflecap_8_8
x373 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[20] adc_array_wafflecap_8_8
x374 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[21] adc_array_wafflecap_8_8
x375 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[22] adc_array_wafflecap_8_8
x376 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[23] adc_array_wafflecap_8_8
x377 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[24] adc_array_wafflecap_8_8
x378 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[25] adc_array_wafflecap_8_8
x379 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[26] adc_array_wafflecap_8_8
x380 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[27] adc_array_wafflecap_8_8
x381 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[28] adc_array_wafflecap_8_8
x382 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[29] adc_array_wafflecap_8_8
x383 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[30] adc_array_wafflecap_8_8
x384 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS col_n[31] adc_array_wafflecap_8_8
x385 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[0] adc_array_wafflecap_8_8
x386 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[1] adc_array_wafflecap_8_8
x387 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[2] adc_array_wafflecap_8_8
x388 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[3] adc_array_wafflecap_8_8
x389 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[4] adc_array_wafflecap_8_8
x390 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[5] adc_array_wafflecap_8_8
x391 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[6] adc_array_wafflecap_8_8
x392 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[7] adc_array_wafflecap_8_8
x393 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[8] adc_array_wafflecap_8_8
x394 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[9] adc_array_wafflecap_8_8
x395 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[10] adc_array_wafflecap_8_8
x396 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[11] adc_array_wafflecap_8_8
x397 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[12] adc_array_wafflecap_8_8
x398 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[13] adc_array_wafflecap_8_8
x399 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[14] adc_array_wafflecap_8_8
x400 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[15] adc_array_wafflecap_8_8
x401 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[16] adc_array_wafflecap_8_8
x402 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[17] adc_array_wafflecap_8_8
x403 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[18] adc_array_wafflecap_8_8
x404 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[19] adc_array_wafflecap_8_8
x405 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[20] adc_array_wafflecap_8_8
x406 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[21] adc_array_wafflecap_8_8
x407 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[22] adc_array_wafflecap_8_8
x408 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[23] adc_array_wafflecap_8_8
x409 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[24] adc_array_wafflecap_8_8
x410 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[25] adc_array_wafflecap_8_8
x411 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[26] adc_array_wafflecap_8_8
x412 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[27] adc_array_wafflecap_8_8
x413 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[28] adc_array_wafflecap_8_8
x414 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[29] adc_array_wafflecap_8_8
x415 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[30] adc_array_wafflecap_8_8
x416 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS col_n[31] adc_array_wafflecap_8_8
x417 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[0] adc_array_wafflecap_8_8
x418 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[1] adc_array_wafflecap_8_8
x419 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[2] adc_array_wafflecap_8_8
x420 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[3] adc_array_wafflecap_8_8
x421 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[4] adc_array_wafflecap_8_8
x422 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[5] adc_array_wafflecap_8_8
x423 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[6] adc_array_wafflecap_8_8
x424 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[7] adc_array_wafflecap_8_8
x425 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[8] adc_array_wafflecap_8_8
x426 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[9] adc_array_wafflecap_8_8
x427 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[10] adc_array_wafflecap_8_8
x428 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[11] adc_array_wafflecap_8_8
x429 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[12] adc_array_wafflecap_8_8
x430 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[13] adc_array_wafflecap_8_8
x431 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[14] adc_array_wafflecap_8_8
x432 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[15] adc_array_wafflecap_8_8
x433 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[16] adc_array_wafflecap_8_8
x434 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[17] adc_array_wafflecap_8_8
x435 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[18] adc_array_wafflecap_8_8
x436 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[19] adc_array_wafflecap_8_8
x437 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[20] adc_array_wafflecap_8_8
x438 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[21] adc_array_wafflecap_8_8
x439 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[22] adc_array_wafflecap_8_8
x440 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[23] adc_array_wafflecap_8_8
x441 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[24] adc_array_wafflecap_8_8
x442 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[25] adc_array_wafflecap_8_8
x443 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[26] adc_array_wafflecap_8_8
x444 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[27] adc_array_wafflecap_8_8
x445 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[28] adc_array_wafflecap_8_8
x446 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[29] adc_array_wafflecap_8_8
x447 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[30] adc_array_wafflecap_8_8
x448 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS col_n[31] adc_array_wafflecap_8_8
x449 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[0] adc_array_wafflecap_8_8
x450 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[1] adc_array_wafflecap_8_8
x451 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[2] adc_array_wafflecap_8_8
x452 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[3] adc_array_wafflecap_8_8
x453 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[4] adc_array_wafflecap_8_8
x454 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[5] adc_array_wafflecap_8_8
x455 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[6] adc_array_wafflecap_8_8
x456 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[7] adc_array_wafflecap_8_8
x457 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[8] adc_array_wafflecap_8_8
x458 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[9] adc_array_wafflecap_8_8
x459 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[10] adc_array_wafflecap_8_8
x460 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[11] adc_array_wafflecap_8_8
x461 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[12] adc_array_wafflecap_8_8
x462 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[13] adc_array_wafflecap_8_8
x463 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[14] adc_array_wafflecap_8_8
x464 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[15] adc_array_wafflecap_8_8
x465 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[16] adc_array_wafflecap_8_8
x466 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[17] adc_array_wafflecap_8_8
x467 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[18] adc_array_wafflecap_8_8
x468 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[19] adc_array_wafflecap_8_8
x469 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[20] adc_array_wafflecap_8_8
x470 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[21] adc_array_wafflecap_8_8
x471 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[22] adc_array_wafflecap_8_8
x472 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[23] adc_array_wafflecap_8_8
x473 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[24] adc_array_wafflecap_8_8
x474 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[25] adc_array_wafflecap_8_8
x475 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[26] adc_array_wafflecap_8_8
x476 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[27] adc_array_wafflecap_8_8
x477 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[28] adc_array_wafflecap_8_8
x478 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[29] adc_array_wafflecap_8_8
x479 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[30] adc_array_wafflecap_8_8
x480 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS col_n[31] adc_array_wafflecap_8_8
x481 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[0] adc_array_wafflecap_8_8
x482 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[1] adc_array_wafflecap_8_8
x483 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[2] adc_array_wafflecap_8_8
x484 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[3] adc_array_wafflecap_8_8
x485 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[4] adc_array_wafflecap_8_8
x486 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[5] adc_array_wafflecap_8_8
x487 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[6] adc_array_wafflecap_8_8
x488 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[7] adc_array_wafflecap_8_8
x489 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[8] adc_array_wafflecap_8_8
x490 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[9] adc_array_wafflecap_8_8
x491 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[10] adc_array_wafflecap_8_8
x492 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[11] adc_array_wafflecap_8_8
x493 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[12] adc_array_wafflecap_8_8
x494 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[13] adc_array_wafflecap_8_8
x495 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[14] adc_array_wafflecap_8_8
x496 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[15] adc_array_wafflecap_8_8
x497 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[16] adc_array_wafflecap_8_8
x498 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[17] adc_array_wafflecap_8_8
x499 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[18] adc_array_wafflecap_8_8
x500 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[19] adc_array_wafflecap_8_8
x501 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[20] adc_array_wafflecap_8_8
x502 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[21] adc_array_wafflecap_8_8
x503 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[22] adc_array_wafflecap_8_8
x504 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[23] adc_array_wafflecap_8_8
x505 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[24] adc_array_wafflecap_8_8
x506 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[25] adc_array_wafflecap_8_8
x507 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[26] adc_array_wafflecap_8_8
x508 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[27] adc_array_wafflecap_8_8
x509 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[28] adc_array_wafflecap_8_8
x510 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[29] adc_array_wafflecap_8_8
x511 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[30] adc_array_wafflecap_8_8
x512 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS col_n[31] adc_array_wafflecap_8_8
x1025 VDD ctop vcm row_n[0] rowon_n[0] sample_n sample VSS VDD net2 net1 adc_array_wafflecap_8_drv
x1026 VDD ctop vcm row_n[1] rowon_n[1] sample_n sample VSS VDD net4 net3 adc_array_wafflecap_8_drv
x1027 VDD ctop vcm row_n[2] rowon_n[2] sample_n sample VSS VDD net6 net5 adc_array_wafflecap_8_drv
x1028 VDD ctop vcm row_n[3] rowon_n[3] sample_n sample VSS VDD net8 net7 adc_array_wafflecap_8_drv
x1029 VDD ctop vcm row_n[4] rowon_n[4] sample_n sample VSS VDD net10 net9 adc_array_wafflecap_8_drv
x1030 VDD ctop vcm row_n[5] rowon_n[5] sample_n sample VSS VDD net12 net11 adc_array_wafflecap_8_drv
x1031 VDD ctop vcm row_n[6] rowon_n[6] sample_n sample VSS VDD net14 net13 adc_array_wafflecap_8_drv
x1032 VDD ctop vcm row_n[7] rowon_n[7] sample_n sample VSS VDD net16 net15 adc_array_wafflecap_8_drv
x1033 VDD ctop vcm row_n[8] rowon_n[8] sample_n sample VSS VDD net18 net17 adc_array_wafflecap_8_drv
x1034 VDD ctop vcm row_n[9] rowon_n[9] sample_n sample VSS VDD net20 net19 adc_array_wafflecap_8_drv
x1035 VDD ctop vcm row_n[10] rowon_n[10] sample_n sample VSS VDD net22 net21
+ adc_array_wafflecap_8_drv
x1036 VDD ctop vcm row_n[11] rowon_n[11] sample_n sample VSS VDD net24 net23
+ adc_array_wafflecap_8_drv
x1037 VDD ctop vcm row_n[12] rowon_n[12] sample_n sample VSS VDD net26 net25
+ adc_array_wafflecap_8_drv
x1038 VDD ctop vcm row_n[13] rowon_n[13] sample_n sample VSS VDD net28 net27
+ adc_array_wafflecap_8_drv
x1039 VDD ctop vcm row_n[14] rowon_n[14] sample_n sample VSS VDD net30 net29
+ adc_array_wafflecap_8_drv
x1040 VDD ctop vcm row_n[15] rowon_n[15] sample_n sample VSS VDD net32 net31
+ adc_array_wafflecap_8_drv
x1058 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[0] adc_array_wafflecap_8_dummy
x1061 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[3] adc_array_wafflecap_8_dummy
x1062 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[4] adc_array_wafflecap_8_dummy
x1063 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[5] adc_array_wafflecap_8_dummy
x1064 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[6] adc_array_wafflecap_8_dummy
x1065 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[7] adc_array_wafflecap_8_dummy
x1067 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[9] adc_array_wafflecap_8_dummy
x1069 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[11] adc_array_wafflecap_8_dummy
x1071 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[13] adc_array_wafflecap_8_dummy
x1072 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[14] adc_array_wafflecap_8_dummy
x1073 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[8] adc_array_wafflecap_8_dummy
x1075 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[24] adc_array_wafflecap_8_dummy
x1077 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[19] adc_array_wafflecap_8_dummy
x1078 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[20] adc_array_wafflecap_8_dummy
x1079 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[21] adc_array_wafflecap_8_dummy
x1080 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[22] adc_array_wafflecap_8_dummy
x1081 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[23] adc_array_wafflecap_8_dummy
x1083 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[25] adc_array_wafflecap_8_dummy
x1085 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[12] adc_array_wafflecap_8_dummy
x1086 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[28] adc_array_wafflecap_8_dummy
x1087 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[29] adc_array_wafflecap_8_dummy
x1088 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[30] adc_array_wafflecap_8_dummy
x1089 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[27] adc_array_wafflecap_8_dummy
x1090 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS VDD adc_array_wafflecap_8_dummy
x1092 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[0] adc_array_wafflecap_8_dummy
x1093 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[1] adc_array_wafflecap_8_dummy
x1094 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[2] adc_array_wafflecap_8_dummy
x1095 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[3] adc_array_wafflecap_8_dummy
x1096 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[4] adc_array_wafflecap_8_dummy
x1097 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[5] adc_array_wafflecap_8_dummy
x1098 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[6] adc_array_wafflecap_8_dummy
x1099 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[7] adc_array_wafflecap_8_dummy
x1100 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[8] adc_array_wafflecap_8_dummy
x1101 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[9] adc_array_wafflecap_8_dummy
x1102 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[10] adc_array_wafflecap_8_dummy
x1103 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[11] adc_array_wafflecap_8_dummy
x1104 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[12] adc_array_wafflecap_8_dummy
x1105 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[13] adc_array_wafflecap_8_dummy
x1106 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[14] adc_array_wafflecap_8_dummy
x1107 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[15] adc_array_wafflecap_8_dummy
x1108 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[16] adc_array_wafflecap_8_dummy
x1109 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[17] adc_array_wafflecap_8_dummy
x1110 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[18] adc_array_wafflecap_8_dummy
x1111 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[19] adc_array_wafflecap_8_dummy
x1112 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[20] adc_array_wafflecap_8_dummy
x1113 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[21] adc_array_wafflecap_8_dummy
x1114 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[22] adc_array_wafflecap_8_dummy
x1115 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[23] adc_array_wafflecap_8_dummy
x1116 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[24] adc_array_wafflecap_8_dummy
x1117 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[25] adc_array_wafflecap_8_dummy
x1118 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[26] adc_array_wafflecap_8_dummy
x1119 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[27] adc_array_wafflecap_8_dummy
x1120 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[28] adc_array_wafflecap_8_dummy
x1121 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[29] adc_array_wafflecap_8_dummy
x1122 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[30] adc_array_wafflecap_8_dummy
x1123 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS col_n[31] adc_array_wafflecap_8_dummy
x1124 VDD ctop vcm rowon_n[15] rowon_n[15] net35 net36 VSS VDD adc_array_wafflecap_8_dummy
x1125 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS VDD adc_array_wafflecap_8_dummy
x1126 VDD ctop vcm row_n[1] rowon_n[1] net4 net3 VSS VDD adc_array_wafflecap_8_dummy
x1127 VDD ctop vcm row_n[2] rowon_n[2] net6 net5 VSS VDD adc_array_wafflecap_8_dummy
x1128 VDD ctop vcm row_n[3] rowon_n[3] net8 net7 VSS VDD adc_array_wafflecap_8_dummy
x1129 VDD ctop vcm row_n[4] rowon_n[4] net10 net9 VSS VDD adc_array_wafflecap_8_dummy
x1130 VDD ctop vcm row_n[5] rowon_n[5] net12 net11 VSS VDD adc_array_wafflecap_8_dummy
x1131 VDD ctop vcm row_n[6] rowon_n[6] net14 net13 VSS VDD adc_array_wafflecap_8_dummy
x1132 VDD ctop vcm row_n[7] rowon_n[7] net16 net15 VSS VDD adc_array_wafflecap_8_dummy
x1133 VDD ctop vcm row_n[8] rowon_n[8] net18 net17 VSS VDD adc_array_wafflecap_8_dummy
x1134 VDD ctop vcm row_n[9] rowon_n[9] net20 net19 VSS VDD adc_array_wafflecap_8_dummy
x1135 VDD ctop vcm row_n[10] rowon_n[10] net22 net21 VSS VDD adc_array_wafflecap_8_dummy
x1136 VDD ctop vcm row_n[11] rowon_n[11] net24 net23 VSS VDD adc_array_wafflecap_8_dummy
x1137 VDD ctop vcm row_n[12] rowon_n[12] net26 net25 VSS VDD adc_array_wafflecap_8_dummy
x1138 VDD ctop vcm row_n[13] rowon_n[13] net28 net27 VSS VDD adc_array_wafflecap_8_dummy
x1139 VDD ctop vcm row_n[14] rowon_n[14] net30 net29 VSS VDD adc_array_wafflecap_8_dummy
x1140 VDD ctop vcm row_n[15] rowon_n[15] net32 net31 VSS VDD adc_array_wafflecap_8_dummy
x513 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[2] adc_array_wafflecap_8_dummy
x514 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[10] adc_array_wafflecap_8_dummy
x515 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[18] adc_array_wafflecap_8_dummy
x516 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[26] adc_array_wafflecap_8_dummy
x517 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[16] en_bit_n[2] adc_array_wafflecap_8_4
x518 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[15] en_bit_n[1] adc_array_wafflecap_8_2
x519 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[17] en_bit_n[0] adc_array_wafflecap_8_1
x520 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[31] sw analog_in sw_n
+ adc_array_wafflecap_8_gate
x14 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[13] adc_array_wafflecap_8_8
x5211 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5212 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5213 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5214 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5215 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5216 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5217 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5218 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x5219 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x52110 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x52111 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x52112 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x52113 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x52114 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x52115 VDD VSS VDD VSS VSS adc_noise_decoup_cell1
x1 VDD ctop vcm row_n[0] rowon_n[0] net2 net1 VSS col_n[0] adc_array_wafflecap_8_dummy
x521 VDD ctop vcm row_n[0] row_n[0] net33 net34 VSS col_n[1] en_C0_n adc_array_wafflecap_8_1
x522 VDD ctop vcm row_n[0] row_n[0] sample_n sample VSS VDD net33 net34 adc_array_wafflecap_8_drv
x523 VDD ctop vcm rowon_n[15] rowon_n[15] sample_n sample VSS VDD net35 net36
+ adc_array_wafflecap_8_drv
.ends

* expanding   symbol:  adc_array_wafflecap_8_8.sym # of pins=9
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_8.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_8.sch
.subckt adc_array_wafflecap_8_8 VDD ctop vcom col_n colon_n sample_n sample VSS row_n
*.PININFO vcom:B VDD:B ctop:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I
C1 ctop cbot 2.90f
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS adc_array_circuit_8
.ends


* expanding   symbol:  adc_array_wafflecap_8_drv.sym # of pins=11
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_drv.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_drv.sch
.subckt adc_array_wafflecap_8_drv VDD ctop vcom col_n colon_n sample_n_i sample_i VSS row_n
+ sample_n_o sample_o
*.PININFO sample_n_i:I sample_i:I vcom:B VDD:B ctop:B VSS:B sample_n_o:O sample_o:O row_n:I col_n:I
*+ colon_n:I
x1 VDD row_n col_n colon_n sample_n_i vcom sample_i VSS sample_n_o sample_o adc_array_circuit_drv
.ends


* expanding   symbol:  adc_array_wafflecap_8_dummy.sym # of pins=9
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_dummy.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_dummy.sch
.subckt adc_array_wafflecap_8_dummy VDD ctop vcom col_n colon_n sample_n sample VSS row_n
*.PININFO vcom:B VDD:B ctop:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS adc_array_circuit_8
.ends


* expanding   symbol:  adc_array_wafflecap_8_4.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_4.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_4.sch
.subckt adc_array_wafflecap_8_4 VDD ctop vcom col_n colon_n sample_n sample VSS row_n en_n
*.PININFO vcom:B VDD:B ctop:B VSS:B en_n:I row_n:I col_n:I colon_n:I sample_n:I sample:I
C3 ctop cbot 1.46f
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS en_n adc_array_circuit_4
.ends


* expanding   symbol:  adc_array_wafflecap_8_2.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_2.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_2.sch
.subckt adc_array_wafflecap_8_2 VDD ctop vcom col_n colon_n sample_n sample VSS row_n en_n
*.PININFO vcom:B VDD:B ctop:B VSS:B en_n:I row_n:I col_n:I colon_n:I sample_n:I sample:I
C3 ctop cbot 0.72f
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS en_n adc_array_circuit_2
.ends


* expanding   symbol:  adc_array_wafflecap_8_1.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_1.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_1.sch
.subckt adc_array_wafflecap_8_1 VDD ctop vcom col_n colon_n sample_n sample VSS row_n en_n
*.PININFO vcom:B VDD:B ctop:B VSS:B en_n:I row_n:I col_n:I colon_n:I sample_n:I sample:I
C3 ctop cbot 0.36f
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS en_n adc_array_circuit_1
.ends


* expanding   symbol:  adc_array_wafflecap_8_gate.sym # of pins=12
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_gate.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_wafflecap_8_gate.sch
.subckt adc_array_wafflecap_8_gate VDD ctop vcom col_n colon_n sample_n sample VSS row_n sw in sw_n
*.PININFO vcom:B VDD:B ctop:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I in:B sw:I sw_n:I
x1 VDD row_n col_n colon_n sample_n vcom sample VSS ctop in sw_n sw adc_array_circuit_gate
.ends


* expanding   symbol:  adc_noise_decoup_cell1.sym # of pins=5
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_noise_decoup_cell1.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_noise_decoup_cell1.sch
.subckt adc_noise_decoup_cell1 mimcap_top mimcap_bot nmoscap_top nmoscap_bot pwell
*.PININFO nmoscap_top:B mimcap_top:B mimcap_bot:B nmoscap_bot:B pwell:B
XC1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 W=17.2 L=17.2 MF=1
M1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 L=16.0 W=16.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_array_circuit_8.sym # of pins=9
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_8.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_8.sch
.subckt adc_array_circuit_8 VDD row_n Cbot col_n colon_n sample_n vcom sample VSS
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B
M1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M5 vint1 col_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M6 VDD row_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M7 VDD colon_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M8 vint2 colon_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M9 VSS row_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M10 VSS col_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_array_circuit_drv.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_drv.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_drv.sch
.subckt adc_array_circuit_drv VDD row_n col_n colon_n sample_n_i vcom sample_i VSS sample_n_o
+ sample_o
*.PININFO sample_n_i:I sample_i:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B sample_o:O
*+ sample_n_o:O
M6 VDD sample_n_i sample_o VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.6 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M7 VDD sample_i sample_n_o VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.6 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M9 VSS sample_i sample_n_o VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M10 VSS sample_n_i sample_o VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_array_circuit_4.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_4.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_4.sch
.subckt adc_array_circuit_4 VDD row_n Cbot col_n colon_n sample_n vcom sample VSS en_n
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B en_n:I
M1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M5 vint1 en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M6 VDD en_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M7 VDD en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M8 vint2 en_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M9 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M10 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_array_circuit_2.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_2.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_2.sch
.subckt adc_array_circuit_2 VDD row_n Cbot col_n colon_n sample_n vcom sample VSS en_n
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B en_n:I
M1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M5 vint1 en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M6 VDD en_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M7 VDD en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M8 vint2 en_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M9 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M10 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_array_circuit_1.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_1.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_1.sch
.subckt adc_array_circuit_1 VDD row_n Cbot col_n colon_n sample_n vcom sample VSS en_n
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B en_n:I
M1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M5 vint1 en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M6 VDD en_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M7 VDD en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M8 vint2 en_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M9 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M10 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_array_circuit_gate.sym # of pins=12
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_gate.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit_gate.sch
.subckt adc_array_circuit_gate VDD row_n col_n colon_n sample_n vcom sample VSS out in sw_n sw
*.PININFO sw:I sw_n:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B sample:I sample_n:I in:B out:B
X1 sw_n in sw out VDD VSS adc_gate_switch
.ends


* expanding   symbol:  adc_gate_switch.sym # of pins=6
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_gate_switch.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_gate_switch.sch
.subckt adc_gate_switch sw_n a sw b VDD VSS
*.PININFO VSS:B VDD:B sw_n:I sw:I a:B b:B
M1 a sw_n b VDD sky130_fd_pr__pfet_01v8 L=0.22 W=7.6 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M3 a sw b VSS sky130_fd_pr__nfet_01v8 L=0.22 W=7.6 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M2 b sw b VDD sky130_fd_pr__pfet_01v8 L=0.22 W=3.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
M4 b sw_n b VSS sky130_fd_pr__nfet_01v8 L=0.22 W=3.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
