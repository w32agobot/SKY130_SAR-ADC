magic
tech sky130A
magscale 1 2
timestamp 1662560087
<< nwell >>
rect -38 250 1970 582
<< pwell >>
rect 1 -17 1931 214
<< nmos >>
rect 196 98 996 182
rect 1190 80 1220 164
rect 1286 80 1316 164
rect 1490 80 1520 164
rect 1586 80 1616 164
<< pmos >>
rect 1168 296 1198 456
rect 1264 296 1294 456
rect 1584 296 1614 456
rect 1680 296 1710 456
<< pmoslvt >>
rect 196 292 996 460
<< ndiff >>
rect 138 170 196 182
rect 138 110 150 170
rect 184 110 196 170
rect 138 98 196 110
rect 996 170 1054 182
rect 996 110 1008 170
rect 1042 110 1054 170
rect 996 98 1054 110
rect 1130 152 1190 164
rect 1130 92 1140 152
rect 1174 92 1190 152
rect 1130 80 1190 92
rect 1220 152 1286 164
rect 1220 92 1236 152
rect 1270 92 1286 152
rect 1220 80 1286 92
rect 1316 152 1374 164
rect 1316 92 1332 152
rect 1366 92 1374 152
rect 1316 80 1374 92
rect 1428 152 1490 164
rect 1428 92 1440 152
rect 1474 92 1490 152
rect 1428 80 1490 92
rect 1520 152 1586 164
rect 1520 92 1536 152
rect 1570 92 1586 152
rect 1520 80 1586 92
rect 1616 152 1678 164
rect 1616 92 1632 152
rect 1666 92 1678 152
rect 1616 80 1678 92
<< pdiff >>
rect 138 448 196 460
rect 138 304 150 448
rect 184 304 196 448
rect 138 292 196 304
rect 996 448 1054 460
rect 996 304 1008 448
rect 1042 304 1054 448
rect 996 292 1054 304
rect 1108 444 1168 456
rect 1108 308 1118 444
rect 1152 308 1168 444
rect 1108 296 1168 308
rect 1198 444 1264 456
rect 1198 308 1214 444
rect 1248 308 1264 444
rect 1198 296 1264 308
rect 1294 444 1354 456
rect 1294 308 1310 444
rect 1344 308 1354 444
rect 1294 296 1354 308
rect 1522 444 1584 456
rect 1522 308 1534 444
rect 1568 308 1584 444
rect 1522 296 1584 308
rect 1614 444 1680 456
rect 1614 308 1630 444
rect 1664 308 1680 444
rect 1614 296 1680 308
rect 1710 444 1770 456
rect 1710 308 1726 444
rect 1760 308 1770 444
rect 1710 296 1770 308
<< ndiffc >>
rect 150 110 184 170
rect 1008 110 1042 170
rect 1140 92 1174 152
rect 1236 92 1270 152
rect 1332 92 1366 152
rect 1440 92 1474 152
rect 1536 92 1570 152
rect 1632 92 1666 152
<< pdiffc >>
rect 150 304 184 448
rect 1008 304 1042 448
rect 1118 308 1152 444
rect 1214 308 1248 444
rect 1310 308 1344 444
rect 1534 308 1568 444
rect 1630 308 1664 444
rect 1726 308 1760 444
<< poly >>
rect 196 460 996 496
rect 1168 456 1198 490
rect 1264 456 1294 490
rect 1584 456 1614 490
rect 1680 456 1710 490
rect 196 266 996 292
rect 1168 280 1198 296
rect 1264 280 1294 296
rect 196 264 322 266
rect 70 248 322 264
rect 70 214 80 248
rect 114 214 322 248
rect 70 208 322 214
rect 1038 250 1126 258
rect 1168 250 1316 280
rect 1038 248 1220 250
rect 1038 214 1076 248
rect 1110 214 1220 248
rect 70 198 996 208
rect 1038 206 1220 214
rect 1038 202 1126 206
rect 196 182 996 198
rect 1190 164 1220 206
rect 1286 164 1316 250
rect 1376 252 1442 262
rect 1376 218 1392 252
rect 1426 220 1442 252
rect 1584 220 1614 296
rect 1680 220 1710 296
rect 1426 218 1710 220
rect 1376 190 1710 218
rect 1490 164 1520 190
rect 1586 164 1616 190
rect 196 72 996 98
rect 1190 54 1220 80
rect 1286 54 1316 80
rect 1490 54 1520 80
rect 1586 54 1616 80
<< polycont >>
rect 80 214 114 248
rect 1076 214 1110 248
rect 1392 218 1426 252
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 150 448 184 464
rect 150 288 184 304
rect 1008 448 1042 464
rect 17 248 118 264
rect 17 214 80 248
rect 114 214 118 248
rect 17 198 118 214
rect 1008 258 1042 304
rect 1118 444 1152 527
rect 1118 292 1152 308
rect 1214 444 1248 460
rect 1214 292 1248 308
rect 1310 444 1344 460
rect 1310 292 1344 308
rect 1008 248 1126 258
rect 1008 214 1054 248
rect 1110 214 1126 248
rect 1008 202 1126 214
rect 1392 252 1426 268
rect 1460 258 1494 527
rect 1528 444 1568 460
rect 1528 308 1534 444
rect 1528 292 1568 308
rect 1630 444 1664 460
rect 1460 224 1570 258
rect 1392 202 1426 218
rect 150 170 184 186
rect 150 94 184 110
rect 1008 170 1042 202
rect 1008 76 1042 110
rect 1140 152 1174 168
rect 1140 17 1174 92
rect 1236 152 1270 168
rect 1236 76 1270 92
rect 1332 76 1366 92
rect 1440 152 1474 168
rect 1440 76 1474 92
rect 1536 152 1570 224
rect 1630 236 1664 308
rect 1726 444 1766 460
rect 1760 308 1766 444
rect 1726 292 1766 308
rect 1771 254 1817 258
rect 1630 202 1734 236
rect 1536 76 1570 92
rect 1632 152 1666 168
rect 1632 76 1666 92
rect 1700 17 1734 202
rect 1771 220 1777 254
rect 1811 220 1817 254
rect 1771 196 1817 220
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 150 304 184 448
rect 1008 304 1042 434
rect 1214 308 1248 444
rect 1310 308 1344 364
rect 1054 214 1076 248
rect 1076 214 1110 248
rect 1392 218 1426 252
rect 1534 328 1568 444
rect 150 110 184 170
rect 1236 92 1270 152
rect 1332 152 1366 178
rect 1332 144 1366 152
rect 1440 92 1474 132
rect 1726 328 1760 444
rect 1632 92 1666 132
rect 1777 220 1811 254
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 144 448 190 496
rect 144 304 150 448
rect 184 304 190 448
rect 144 292 190 304
rect 1002 434 1048 456
rect 1002 304 1008 434
rect 1042 304 1048 434
rect 1002 258 1048 304
rect 1208 444 1766 456
rect 1208 308 1214 444
rect 1248 422 1534 444
rect 1248 308 1254 422
rect 1208 296 1254 308
rect 1304 364 1350 394
rect 1304 308 1310 364
rect 1344 308 1350 364
rect 1528 328 1534 422
rect 1568 422 1726 444
rect 1568 328 1574 422
rect 1528 316 1574 328
rect 1720 328 1726 422
rect 1760 328 1766 444
rect 1720 316 1766 328
rect 1002 248 1126 258
rect 1002 214 1054 248
rect 1110 214 1126 248
rect 1304 248 1350 308
rect 1386 252 1432 264
rect 1386 248 1392 252
rect 1304 220 1392 248
rect 1002 202 1126 214
rect 1326 218 1392 220
rect 1426 248 1432 252
rect 1765 254 1823 260
rect 1765 248 1777 254
rect 1426 220 1777 248
rect 1811 220 1823 254
rect 1426 218 1432 220
rect 1326 206 1432 218
rect 1765 214 1823 220
rect 144 170 190 182
rect 144 110 150 170
rect 184 110 190 170
rect 1326 178 1372 206
rect 1230 152 1276 164
rect 144 48 190 110
rect 1004 48 1108 136
rect 1230 92 1236 152
rect 1270 104 1276 152
rect 1326 144 1332 178
rect 1366 144 1372 178
rect 1326 132 1372 144
rect 1434 132 1480 144
rect 1434 104 1440 132
rect 1270 92 1440 104
rect 1474 104 1480 132
rect 1626 132 1672 144
rect 1626 104 1632 132
rect 1474 92 1632 104
rect 1666 92 1672 132
rect 1230 76 1672 92
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali 1008 172 1042 172 1 cap_top
flabel metal1 s 0 -48 1932 48 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 0 496 1932 592 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 30 221 64 255 7 FreeSans 160 0 0 0 in
port 1 nsew signal input
flabel metal1 s 1777 220 1811 254 0 FreeSans 160 0 0 0 out
port 2 nsew signal output
flabel nwell s 213 527 247 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 213 527 247 561 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel pwell s 213 -17 247 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 213 -17 247 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
string LEFsource USER
string LEFsymmetry X Y R90
<< end >>
