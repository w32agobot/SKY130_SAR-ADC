* SPICE3 file created from adc_array_fingercap_8(8)x386aF_topB_22um2.ext - technology: sky130A

C0 VSS cbot 3.09fF
C1 ctop cbot 2.75fF
C2 VSS ctop 1.03fF
C3 ctop VSUBS 1.00fF
C4 cbot VSUBS 0.43fF
C5 VSS VSUBS 1.80fF
