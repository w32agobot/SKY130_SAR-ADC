* NGSPICE file created from adc_vcm_generator.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
C0 VPWR VGND 0.03fF
C1 VPB Y 0.02fF
C2 VPB VPWR 0.06fF
C3 A VGND 0.04fF
C4 Y VPWR 0.13fF
C5 A VPB 0.07fF
C6 A Y 0.05fF
C7 VPB VGND 0.01fF
C8 A VPWR 0.05fF
C9 Y VGND 0.10fF
C10 VGND VNB 0.24fF
C11 Y VNB 0.08fF
C12 VPWR VNB 0.21fF
C13 A VNB 0.12fF
C14 VPB VNB 0.34fF
.ends

.subckt pfet_01v8_w500_l500_nf2 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26# VSUBS
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
C0 a_29_n26# w_n224_n36# 0.06fF
C1 a_n129_n26# a_n29_0# 0.00fF
C2 a_n129_n26# a_n187_0# 0.00fF
C3 a_29_n26# a_129_0# 0.00fF
C4 w_n224_n36# a_129_0# 0.00fF
C5 a_29_n26# a_n129_n26# 0.01fF
C6 a_n29_0# a_n187_0# 0.02fF
C7 a_n129_n26# w_n224_n36# 0.06fF
C8 a_29_n26# a_n29_0# 0.00fF
C9 w_n224_n36# a_n29_0# 0.00fF
C10 w_n224_n36# a_n187_0# 0.00fF
C11 a_n29_0# a_129_0# 0.02fF
C12 a_129_0# VSUBS 0.04fF
C13 a_n29_0# VSUBS 0.02fF
C14 a_n187_0# VSUBS 0.04fF
C15 a_29_n26# VSUBS 0.08fF
C16 a_n129_n26# VSUBS 0.08fF
C17 w_n224_n36# VSUBS 0.23fF
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 VGND a_27_47# 0.21fF
C1 A X 0.00fF
C2 VPWR a_27_47# 0.26fF
C3 VGND VPWR 0.07fF
C4 a_27_47# A 0.20fF
C5 VPB X 0.02fF
C6 VGND A 0.02fF
C7 VPWR A 0.02fF
C8 VPB a_27_47# 0.20fF
C9 VPB VGND 0.01fF
C10 VPB VPWR 0.08fF
C11 a_27_47# X 0.29fF
C12 VGND X 0.23fF
C13 VPB A 0.06fF
C14 VPWR X 0.31fF
C15 VGND VNB 0.31fF
C16 X VNB -0.24fF
C17 VPWR VNB 0.24fF
C18 A VNB 0.11fF
C19 VPB VNB 0.60fF
C20 a_27_47# VNB 0.29fF
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VPWR X a_240_47# VNB VPB a_629_47#
+ a_523_47# a_346_47# a_63_47#
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=5.82e+11p ps=5.85e+06u w=650000u l=150000u
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.445e+11p pd=7.95e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
C0 A a_346_47# 0.00fF
C1 VGND X 0.09fF
C2 A VGND 0.02fF
C3 a_63_47# X 0.00fF
C4 A a_63_47# 0.27fF
C5 a_346_47# VGND 0.13fF
C6 a_346_47# a_63_47# 0.00fF
C7 a_240_47# a_629_47# 0.00fF
C8 a_63_47# VGND 0.16fF
C9 VPWR a_240_47# 0.10fF
C10 a_240_47# a_523_47# 0.02fF
C11 VPB a_240_47# 0.15fF
C12 a_240_47# X 0.00fF
C13 A a_240_47# 0.02fF
C14 VPWR a_629_47# 0.15fF
C15 a_346_47# a_240_47# 0.31fF
C16 a_629_47# a_523_47# 0.32fF
C17 a_240_47# VGND 0.10fF
C18 a_240_47# a_63_47# 0.17fF
C19 VPB a_629_47# 0.07fF
C20 VPWR a_523_47# 0.09fF
C21 a_629_47# X 0.14fF
C22 A a_629_47# 0.00fF
C23 VPB VPWR 0.12fF
C24 a_346_47# a_629_47# 0.00fF
C25 VPB a_523_47# 0.15fF
C26 VGND a_629_47# 0.14fF
C27 a_63_47# a_629_47# 0.00fF
C28 VPWR X 0.10fF
C29 A VPWR 0.02fF
C30 X a_523_47# 0.01fF
C31 A a_523_47# 0.00fF
C32 a_346_47# VPWR 0.14fF
C33 VPWR VGND 0.09fF
C34 a_346_47# a_523_47# 0.16fF
C35 VPWR a_63_47# 0.16fF
C36 VPB X 0.03fF
C37 VGND a_523_47# 0.09fF
C38 A VPB 0.12fF
C39 a_63_47# a_523_47# 0.00fF
C40 A X 0.00fF
C41 VPB a_346_47# 0.07fF
C42 VPB VGND 0.01fF
C43 VPB a_63_47# 0.07fF
C44 a_346_47# X 0.00fF
C45 VGND VNB 0.46fF
C46 X VNB 0.04fF
C47 VPWR VNB 0.34fF
C48 A VNB 0.18fF
C49 VPB VNB 0.96fF
C50 a_629_47# VNB 0.03fF
C51 a_523_47# VNB 0.07fF
C52 a_346_47# VNB -0.00fF
C53 a_240_47# VNB 0.07fF
C54 a_63_47# VNB 0.05fF
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 nmoscap_top nmoscap_bot pwell sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
C0 nmoscap_bot mimcap_top 0.32fF
C1 nmoscap_top nmoscap_bot 303.08fF
C2 mimcap_bot nmoscap_bot 34.51fF
C3 nmoscap_top mimcap_top 2.71fF
C4 mimcap_bot mimcap_top 33.65fF
C5 mimcap_bot nmoscap_top 30.43fF
C6 mimcap_top pwell 1.83fF
C7 mimcap_bot pwell 0.60fF
C8 nmoscap_top pwell -17.39fF
C9 nmoscap_bot pwell 31.87fF
.ends

.subckt nfet_01v8_w500_l500_nf2 a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76# a_129_n50#
+ VSUBS
X0 a_129_n50# a_29_n76# a_n29_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_n50# a_n129_n76# a_n187_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
C0 a_n129_n76# a_n29_n50# 0.00fF
C1 a_29_n76# a_n129_n76# 0.01fF
C2 a_n187_n50# a_n129_n76# 0.00fF
C3 a_29_n76# a_n29_n50# 0.00fF
C4 a_n29_n50# a_129_n50# 0.02fF
C5 a_n187_n50# a_n29_n50# 0.02fF
C6 a_29_n76# a_129_n50# 0.00fF
C7 a_129_n50# VSUBS 0.04fF
C8 a_n29_n50# VSUBS 0.02fF
C9 a_n187_n50# VSUBS 0.04fF
C10 a_29_n76# VSUBS 0.14fF
C11 a_n129_n76# VSUBS 0.14fF
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VPWR A 0.06fF
C1 VPB VPWR 0.05fF
C2 Y A 0.12fF
C3 Y VPB 0.01fF
C4 VGND A 0.01fF
C5 VPB VGND 0.01fF
C6 Y VPWR 0.22fF
C7 VGND VPWR 0.03fF
C8 VPWR a_113_47# 0.00fF
C9 Y VGND 0.16fF
C10 Y a_113_47# 0.01fF
C11 VGND a_113_47# 0.00fF
C12 B A 0.05fF
C13 VPB B 0.05fF
C14 B VPWR 0.06fF
C15 VPB A 0.05fF
C16 Y B 0.05fF
C17 B VGND 0.07fF
C18 VGND VNB 0.21fF
C19 Y VNB -0.07fF
C20 VPWR VNB 0.22fF
C21 A VNB 0.12fF
C22 B VNB 0.12fF
C23 VPB VNB 0.34fF
.ends

.subckt adc_vcm_generator VDD VSS clk vcm
Xsky130_fd_sc_hd__inv_1_4 clk VSS VDD sky130_fd_sc_hd__inv_1_4/Y VSS VDD sky130_fd_sc_hd__inv_1
Xpfet_01v8_w500_l500_nf2_0 mimtop2 vcm phi1_n VDD vcm phi1_n VSS pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_1 mimtop1 vcm phi1_n VDD vcm phi1_n VSS pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_0 sky130_fd_sc_hd__inv_1_2/A VSS VDD phi1 VSS VDD sky130_fd_sc_hd__buf_4_0/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_2 mimtop2 mimbot1 phi2_n VDD mimbot1 phi2_n VSS pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_1 sky130_fd_sc_hd__inv_1_2/Y VSS VDD phi1_n VSS VDD sky130_fd_sc_hd__buf_4_1/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_3 VDD mimtop1 phi2_n VDD mimtop1 phi2_n VSS pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_4 mimbot1 VSS phi1_n VDD VSS phi1_n VSS pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_2 sky130_fd_sc_hd__inv_1_3/A VSS VDD phi2 VSS VDD sky130_fd_sc_hd__buf_4_2/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_3 sky130_fd_sc_hd__inv_1_3/Y VSS VDD phi2_n VSS VDD sky130_fd_sc_hd__buf_4_3/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 sky130_fd_sc_hd__nand2_1_0/Y VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_3/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VSS VDD sky130_fd_sc_hd__inv_1_0/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VSS VDD sky130_fd_sc_hd__inv_1_1/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xnfet_01v8_w500_l500_nf2_0 phi1 mimtop2 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_1 phi1 mimtop1 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_0 clk sky130_fd_sc_hd__inv_1_3/Y VSS VDD sky130_fd_sc_hd__nand2_1_0/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_2 phi2 mimtop2 mimbot1 phi2 mimbot1 VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_3 phi2 VDD mimtop1 phi2 mimtop1 VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_4/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_4 phi1 mimbot1 VSS phi1 VSS VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A VSS VDD sky130_fd_sc_hd__inv_1_2/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/A VSS VDD sky130_fd_sc_hd__inv_1_3/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VSS VDD sky130_fd_sc_hd__inv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/A VSS VDD sky130_fd_sc_hd__inv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
C0 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C1 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C3 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C4 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C5 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C6 vcm sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.03fF
C7 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C8 sky130_fd_sc_hd__inv_1_3/Y vcm 0.59fF
C9 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 0.00fF
C10 phi1 mimtop1 0.24fF
C11 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# vcm 0.00fF
C12 mimbot1 mimtop1 11.31fF
C13 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C14 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C15 sky130_fd_sc_hd__inv_1_3/A VDD 0.32fF
C16 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C17 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.00fF
C18 VDD sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.01fF
C19 clk sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C20 sky130_fd_sc_hd__inv_1_3/Y clk 0.01fF
C21 sky130_fd_sc_hd__inv_1_3/Y VDD 1.70fF
C22 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C23 sky130_fd_sc_hd__nand2_1_1/a_113_47# mimbot1 0.00fF
C24 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__inv_1_3/Y 0.08fF
C25 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C26 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_3/A 0.00fF
C27 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# -0.00fF
C28 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C29 mimtop1 sky130_fd_sc_hd__nand2_1_0/Y 0.04fF
C30 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C31 phi1 sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C32 mimbot1 sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C33 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_2/A 0.00fF
C34 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.02fF
C35 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C36 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C37 mimtop1 phi1_n 0.17fF
C38 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C39 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# VDD 0.12fF
C40 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_3/A 0.00fF
C41 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__buf_4_2/a_27_47# 0.26fF
C42 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C43 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C44 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C45 mimtop1 phi2_n 0.09fF
C46 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# vcm 0.00fF
C47 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C48 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.01fF
C49 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C50 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_1/Y 0.01fF
C51 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A -0.00fF
C52 phi1_n sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C53 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C54 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# mimbot1 0.00fF
C55 phi2_n sky130_fd_sc_hd__nand2_1_1/Y 0.01fF
C56 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C57 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C58 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# VDD 0.02fF
C59 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C60 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# clk 0.00fF
C61 phi1 vcm 0.24fF
C62 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C63 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C64 mimbot1 vcm 8.24fF
C65 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C66 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# -0.00fF
C67 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__inv_1_2/Y 0.03fF
C68 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# vcm 0.01fF
C69 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C70 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__inv_1_2/Y 0.07fF
C71 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C72 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# vcm 0.03fF
C73 sky130_fd_sc_hd__nand2_1_0/Y vcm 0.27fF
C74 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C75 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.06fF
C76 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# mimtop1 0.00fF
C77 sky130_fd_sc_hd__dlymetal6s6s_1_3/A phi2 0.00fF
C78 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C79 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C80 phi1_n vcm 0.32fF
C81 phi1 VDD 0.41fF
C82 phi1 clk 0.00fF
C83 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# phi1 0.00fF
C84 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.01fF
C85 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.05fF
C86 mimbot1 VDD 3.15fF
C87 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C88 mimbot1 clk 0.01fF
C89 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 0.00fF
C90 vcm phi2_n 0.05fF
C91 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C92 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C93 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C94 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00fF
C95 phi1 sky130_fd_sc_hd__inv_1_2/A 0.00fF
C96 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# -0.00fF
C97 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# VDD 0.05fF
C98 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C99 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# clk 0.00fF
C100 mimbot1 sky130_fd_sc_hd__inv_1_2/A 0.01fF
C101 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.01fF
C102 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C103 phi1 sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C104 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__inv_1_2/Y 0.07fF
C105 mimbot1 sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C106 sky130_fd_sc_hd__dlymetal6s6s_1_4/A phi1_n 0.00fF
C107 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C108 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# VDD 0.05fF
C109 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# clk 0.00fF
C110 sky130_fd_sc_hd__nand2_1_0/Y clk 0.05fF
C111 sky130_fd_sc_hd__nand2_1_0/Y VDD 0.16fF
C112 sky130_fd_sc_hd__inv_1_0/A phi1 0.00fF
C113 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C114 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C115 sky130_fd_sc_hd__dlymetal6s6s_1_4/A phi2_n 0.00fF
C116 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.01fF
C117 sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C118 VDD phi1_n 1.72fF
C119 phi1_n clk 0.00fF
C120 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# phi1_n 0.01fF
C121 VDD phi2_n 1.35fF
C122 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# phi2_n 0.00fF
C123 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C124 sky130_fd_sc_hd__inv_1_2/A phi1_n 0.00fF
C125 mimtop2 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C126 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 0.00fF
C127 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C128 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C129 sky130_fd_sc_hd__inv_1_0/A phi1_n 0.00fF
C130 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C131 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 0.01fF
C132 sky130_fd_sc_hd__buf_4_2/a_27_47# phi2_n 0.00fF
C133 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.02fF
C134 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C135 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C136 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C137 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C138 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# vcm 0.00fF
C139 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A 0.22fF
C140 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.07fF
C141 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C142 phi2 mimtop1 0.04fF
C143 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C144 sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C145 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C146 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C147 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C148 sky130_fd_sc_hd__buf_4_0/a_27_47# vcm 0.00fF
C149 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__inv_1_3/Y 0.03fF
C150 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# VDD 0.03fF
C151 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C152 phi2 sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C153 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# clk 0.00fF
C154 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C155 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C156 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00fF
C157 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C158 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C159 phi1 sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C160 mimbot1 sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C161 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C162 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C163 sky130_fd_sc_hd__buf_4_0/a_27_47# VDD 0.16fF
C164 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C165 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C166 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00fF
C167 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C168 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C169 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C170 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# vcm 0.00fF
C171 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C172 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C173 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.06fF
C174 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# vcm 0.09fF
C175 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C176 sky130_fd_sc_hd__inv_1_4/Y phi1_n 0.00fF
C177 VDD sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.03fF
C178 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C179 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__inv_1_0/A 0.00fF
C180 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C181 phi2 vcm 0.04fF
C182 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C183 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C184 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C185 mimbot1 sky130_fd_sc_hd__inv_1_3/A 0.00fF
C186 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.01fF
C187 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# VDD 0.04fF
C188 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# vcm 0.00fF
C189 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C190 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# clk 0.00fF
C191 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C192 phi1 sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C193 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.01fF
C194 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C195 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__inv_1_2/Y 0.03fF
C196 mimbot1 sky130_fd_sc_hd__inv_1_3/Y 0.28fF
C197 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# clk 0.00fF
C198 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C199 VDD sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.06fF
C200 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C201 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A -0.00fF
C202 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A -0.00fF
C203 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C204 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C205 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C206 phi2 VDD 0.61fF
C207 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C208 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.01fF
C209 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.01fF
C210 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# phi2 0.00fF
C211 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C212 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C213 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C214 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nand2_1_0/Y 0.28fF
C215 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C216 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C217 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.00fF
C218 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.01fF
C219 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C220 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# VDD 0.08fF
C221 sky130_fd_sc_hd__inv_1_3/Y phi1_n 0.02fF
C222 sky130_fd_sc_hd__inv_1_3/A phi2_n 0.00fF
C223 phi2 sky130_fd_sc_hd__buf_4_2/a_27_47# 0.03fF
C224 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C225 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C226 mimtop1 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C227 sky130_fd_sc_hd__inv_1_3/Y phi2_n 0.01fF
C228 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C229 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C230 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.01fF
C231 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C232 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# VDD 0.04fF
C233 mimtop1 sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C234 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C235 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C236 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C237 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C238 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C239 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C240 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C241 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 0.03fF
C242 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# phi1_n 0.00fF
C243 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C244 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# mimtop1 0.00fF
C245 mimbot1 phi1 0.10fF
C246 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_2/Y 0.31fF
C247 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# phi2_n 0.00fF
C248 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C249 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C250 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C251 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C252 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C253 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__inv_1_3/Y 0.06fF
C254 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C255 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C256 mimtop2 mimtop1 0.02fF
C257 phi1 sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C258 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C259 sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C260 vcm sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C261 mimbot1 sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C262 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C263 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C264 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C265 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C266 phi1 phi1_n 0.91fF
C267 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C268 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.00fF
C269 mimbot1 phi1_n 0.19fF
C270 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C271 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C272 mimbot1 phi2_n 0.20fF
C273 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.02fF
C274 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# phi1_n 0.00fF
C275 mimtop2 sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C276 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C277 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# phi2_n 0.01fF
C278 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C279 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# phi1_n 0.00fF
C280 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C281 sky130_fd_sc_hd__nand2_1_0/Y phi1_n 0.01fF
C282 vcm sky130_fd_sc_hd__inv_1_2/Y 0.52fF
C283 VDD sky130_fd_sc_hd__buf_4_3/a_27_47# 0.21fF
C284 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.00fF
C285 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C286 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C287 sky130_fd_sc_hd__nand2_1_0/Y phi2_n 0.00fF
C288 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# phi2_n 0.00fF
C289 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C290 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# mimtop1 0.00fF
C291 phi1_n phi2_n 0.00fF
C292 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C293 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C294 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C295 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# vcm 0.00fF
C296 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C297 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# 0.00fF
C298 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__inv_1_2/Y 0.09fF
C299 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.07fF
C300 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# vcm 0.00fF
C301 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.08fF
C302 VDD sky130_fd_sc_hd__inv_1_2/Y 0.62fF
C303 clk sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C304 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C305 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C306 phi2 sky130_fd_sc_hd__inv_1_3/A 0.00fF
C307 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C308 mimtop2 vcm 4.08fF
C309 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.03fF
C310 sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.03fF
C311 phi2 sky130_fd_sc_hd__inv_1_3/Y 0.43fF
C312 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_2/Y 0.21fF
C313 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# phi1 0.00fF
C314 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# VDD 0.05fF
C315 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# clk 0.00fF
C316 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.02fF
C317 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.00fF
C318 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.01fF
C319 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/Y 0.03fF
C320 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# VDD 0.01fF
C321 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C322 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# phi2 0.00fF
C323 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# clk 0.00fF
C324 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C325 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C326 sky130_fd_sc_hd__buf_4_0/a_27_47# phi1 0.02fF
C327 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C328 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C329 mimtop2 VDD 2.02fF
C330 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.09fF
C331 sky130_fd_sc_hd__buf_4_0/a_27_47# mimbot1 0.01fF
C332 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 0.06fF
C333 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C334 sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C335 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# phi1_n 0.00fF
C336 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C337 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C338 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C339 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# vcm 0.00fF
C340 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# phi2_n 0.00fF
C341 mimtop2 sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C342 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C343 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C344 sky130_fd_sc_hd__buf_4_0/a_27_47# phi1_n 0.00fF
C345 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C346 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C347 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.01fF
C348 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C349 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.04fF
C350 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C351 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C352 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# VDD 0.09fF
C353 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# clk 0.00fF
C354 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.01fF
C355 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.01fF
C356 phi1 phi2 0.00fF
C357 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C358 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C359 mimbot1 phi2 0.13fF
C360 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C361 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.04fF
C362 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C363 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C364 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# phi1_n 0.00fF
C365 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C366 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C367 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C368 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C369 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.06fF
C370 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.01fF
C371 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# vcm 0.05fF
C372 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# phi1_n 0.01fF
C373 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# phi2_n 0.00fF
C374 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C375 phi2 sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C376 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C377 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# phi2_n 0.00fF
C378 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C379 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C380 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C381 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C382 phi2 phi2_n 0.75fF
C383 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__buf_4_3/a_27_47# 0.07fF
C384 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# phi1_n 0.00fF
C385 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 0.00fF
C386 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# VDD 0.02fF
C387 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# clk 0.00fF
C388 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# phi2_n 0.00fF
C389 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.01fF
C390 vcm sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.09fF
C391 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C392 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C393 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C394 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C395 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_2/Y 0.29fF
C396 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C397 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# -0.00fF
C398 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__inv_1_2/Y 0.05fF
C399 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C400 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C401 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A -0.00fF
C402 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C403 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C404 VDD sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.11fF
C405 clk sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C406 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__inv_1_3/Y 0.07fF
C407 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C408 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C409 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C410 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.01fF
C411 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C412 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# phi2 0.00fF
C413 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.02fF
C414 mimtop2 sky130_fd_sc_hd__inv_1_3/Y 0.23fF
C415 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C416 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C417 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C418 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C419 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C420 sky130_fd_sc_hd__buf_4_0/a_27_47# phi2 0.00fF
C421 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C422 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C423 phi1 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C424 mimbot1 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.01fF
C425 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C426 vcm sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C427 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C428 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# VDD 0.03fF
C429 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00fF
C430 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C431 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C432 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.01fF
C433 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C434 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C435 phi1_n sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C436 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C437 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C438 phi1 sky130_fd_sc_hd__inv_1_2/Y 0.38fF
C439 mimbot1 sky130_fd_sc_hd__inv_1_2/Y 0.34fF
C440 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C441 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C442 phi2_n sky130_fd_sc_hd__buf_4_3/a_27_47# 0.03fF
C443 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# vcm 0.00fF
C444 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C445 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C446 VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.08fF
C447 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__inv_1_2/Y 0.06fF
C448 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C449 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# phi1 0.00fF
C450 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__inv_1_2/Y 0.08fF
C451 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C452 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.02fF
C453 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C454 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.01fF
C455 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.02fF
C456 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C457 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C458 phi1_n sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C459 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C460 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C461 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C462 phi2_n sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C463 mimtop2 phi1 0.09fF
C464 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C465 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C466 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# VDD 0.10fF
C467 mimtop2 mimbot1 1.57fF
C468 VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.04fF
C469 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/A -0.00fF
C470 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C471 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C472 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# phi1_n 0.00fF
C473 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C474 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.06fF
C475 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C476 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# phi1_n 0.01fF
C477 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# phi2_n 0.01fF
C478 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C479 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C480 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.01fF
C481 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.02fF
C482 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.08fF
C483 mimtop2 sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C484 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# phi2_n 0.00fF
C485 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C486 mimtop2 phi1_n 0.14fF
C487 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C488 mimtop2 phi2_n 0.10fF
C489 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C490 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# phi1 0.00fF
C491 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C492 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C493 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.01fF
C494 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C495 mimtop1 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C496 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C497 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C498 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C499 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.01fF
C500 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C501 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C502 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C503 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C504 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C505 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# mimtop1 0.00fF
C506 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C507 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# phi1_n 0.00fF
C508 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C509 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.24fF
C510 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# phi2_n 0.00fF
C511 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C512 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C513 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C514 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C515 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__nand2_1_1/Y 0.01fF
C516 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C517 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00fF
C518 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C519 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C520 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C521 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# vcm 0.00fF
C522 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C523 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C524 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C525 phi2 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.19fF
C526 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# vcm 0.00fF
C527 sky130_fd_sc_hd__buf_4_0/a_27_47# mimtop2 0.00fF
C528 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C529 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C530 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.01fF
C531 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C532 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C533 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__nand2_1_0/Y 0.01fF
C534 sky130_fd_sc_hd__buf_4_1/a_27_47# vcm 0.00fF
C535 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C536 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C537 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.09fF
C538 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# phi1_n 0.01fF
C539 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.04fF
C540 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# VDD 0.06fF
C541 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.02fF
C542 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C543 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# vcm 0.05fF
C544 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# phi2_n 0.00fF
C545 phi2 sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C546 VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.11fF
C547 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# clk 0.00fF
C548 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C549 mimtop1 sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C550 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.01fF
C551 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C552 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C553 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C554 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C555 sky130_fd_sc_hd__inv_1_1/A VDD 0.38fF
C556 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__inv_1_2/Y 0.06fF
C557 vcm sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C558 sky130_fd_sc_hd__buf_4_1/a_27_47# VDD 0.20fF
C559 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C560 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# phi2 0.00fF
C561 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C562 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C563 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A -0.00fF
C564 sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C565 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_2/A 0.00fF
C566 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.02fF
C567 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00fF
C568 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C569 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C570 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C571 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# VDD 0.04fF
C572 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C573 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C574 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# VDD 0.04fF
C575 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# clk 0.00fF
C576 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C577 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.01fF
C578 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_0/A 0.01fF
C579 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C580 mimtop2 phi2 0.12fF
C581 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C582 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C583 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C584 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C585 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C586 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.01fF
C587 VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.05fF
C588 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.01fF
C589 sky130_fd_sc_hd__dlymetal6s6s_1_2/A clk 0.00fF
C590 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.01fF
C591 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C592 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C593 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C594 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# mimbot1 0.00fF
C595 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C596 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C597 vcm sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C598 sky130_fd_sc_hd__nand2_1_0/a_113_47# vcm 0.00fF
C599 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.08fF
C600 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C601 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C602 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# phi2 0.00fF
C603 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C604 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A -0.00fF
C605 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C606 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# VDD 0.04fF
C607 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C608 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C609 VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.11fF
C610 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C611 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C612 sky130_fd_sc_hd__nand2_1_0/a_113_47# VDD -0.00fF
C613 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C614 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C615 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C616 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.01fF
C617 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C618 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.01fF
C619 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C620 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C621 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C622 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C623 sky130_fd_sc_hd__dlymetal6s6s_1_3/A vcm 0.00fF
C624 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C625 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00fF
C626 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# vcm 0.00fF
C627 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C628 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C629 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.06fF
C630 sky130_fd_sc_hd__nand2_1_1/a_113_47# mimtop1 0.00fF
C631 mimtop2 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00fF
C632 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# VDD 0.05fF
C633 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C634 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VDD 0.08fF
C635 mimtop1 sky130_fd_sc_hd__nand2_1_1/Y 0.03fF
C636 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.00fF
C637 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_3/A 0.05fF
C638 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__inv_1_2/Y 0.08fF
C639 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C640 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.01fF
C641 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.01fF
C642 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C643 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_3/Y 0.04fF
C644 VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.04fF
C645 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C646 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C647 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C648 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C649 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C650 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C651 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C652 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__inv_1_0/A 0.00fF
C653 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C654 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C655 mimtop2 sky130_fd_sc_hd__inv_1_2/Y 0.21fF
C656 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C657 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C658 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C659 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.01fF
C660 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.01fF
C661 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C662 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C663 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C664 sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# -0.00fF
C665 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.11fF
C666 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.01fF
C667 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.05fF
C668 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C669 mimtop1 vcm 5.68fF
C670 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.06fF
C671 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# vcm 0.00fF
C672 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C673 sky130_fd_sc_hd__nand2_1_1/a_113_47# vcm 0.00fF
C674 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.01fF
C675 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C676 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__inv_1_2/Y 0.05fF
C677 vcm sky130_fd_sc_hd__nand2_1_1/Y 0.26fF
C678 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00fF
C679 mimtop1 VDD 2.23fF
C680 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C681 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C682 mimtop1 clk 0.18fF
C683 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# mimtop1 0.00fF
C684 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.01fF
C685 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C686 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C687 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C688 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C689 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.03fF
C690 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C691 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C692 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# VDD 0.08fF
C693 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.00fF
C694 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C695 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C696 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.05fF
C697 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C698 sky130_fd_sc_hd__nand2_1_1/a_113_47# VDD 0.00fF
C699 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C700 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C701 phi1 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.18fF
C702 VDD sky130_fd_sc_hd__nand2_1_1/Y 0.19fF
C703 mimbot1 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.03fF
C704 sky130_fd_sc_hd__nand2_1_1/Y clk 0.01fF
C705 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C706 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__buf_4_2/a_27_47# 0.00fF
C707 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00fF
C708 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 0.00fF
C709 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.01fF
C710 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# phi1 0.00fF
C711 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__inv_1_0/A 0.00fF
C712 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# phi1_n 0.00fF
C713 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C714 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# mimbot1 0.00fF
C715 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00fF
C716 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# phi2_n 0.00fF
C717 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C718 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C719 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.06fF
C720 sky130_fd_sc_hd__buf_4_1/a_27_47# phi1_n 0.04fF
C721 sky130_fd_sc_hd__inv_1_1/A phi2_n 0.00fF
C722 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# VDD 0.04fF
C723 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C724 sky130_fd_sc_hd__buf_4_1/a_27_47# phi2_n 0.00fF
C725 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00fF
C726 sky130_fd_sc_hd__dlymetal6s6s_1_4/A vcm 0.00fF
C727 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C728 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C729 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# phi1_n 0.00fF
C730 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C731 VDD vcm 49.83fF
C732 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# phi2_n 0.01fF
C733 vcm clk 0.01fF
C734 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# vcm 0.01fF
C735 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C736 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C737 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C738 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.01fF
C739 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__inv_1_3/Y 0.03fF
C740 sky130_fd_sc_hd__dlymetal6s6s_1_2/A phi2_n 0.00fF
C741 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.01fF
C742 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.01fF
C743 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VDD 0.15fF
C744 sky130_fd_sc_hd__dlymetal6s6s_1_4/A clk 0.00fF
C745 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C746 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.11fF
C747 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.07fF
C748 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C749 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C750 VDD clk 0.30fF
C751 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C752 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# VDD 0.02fF
C753 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# clk 0.00fF
C754 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C755 mimtop1 sky130_fd_sc_hd__inv_1_4/Y 0.04fF
C756 mimbot1 sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C757 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C758 sky130_fd_sc_hd__inv_1_2/A VDD 0.31fF
C759 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C760 sky130_fd_sc_hd__buf_4_2/a_27_47# VDD 0.16fF
C761 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__buf_4_1/a_27_47# 0.01fF
C762 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00fF
C763 sky130_fd_sc_hd__inv_1_0/A VDD 0.37fF
C764 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C765 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C766 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__nand2_1_1/Y 0.02fF
C767 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C768 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/A 0.04fF
C769 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# -0.00fF
C770 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C771 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C772 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C773 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00fF
C774 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00fF
C775 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.00fF
C776 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C777 mimtop1 sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C778 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00fF
C779 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# sky130_fd_sc_hd__inv_1_2/Y 0.03fF
C780 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.01fF
C781 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00fF
C782 sky130_fd_sc_hd__dlymetal6s6s_1_3/A phi1 0.00fF
C783 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00fF
C784 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.00fF
C785 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C786 sky130_fd_sc_hd__inv_1_4/Y vcm 0.01fF
C787 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00fF
C788 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00fF
C789 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C790 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C791 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C792 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00fF
C793 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C794 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00fF
C795 sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00fF
C796 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__nand2_1_0/Y 0.00fF
C797 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00fF
C798 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C799 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00fF
C800 sky130_fd_sc_hd__inv_1_1/A phi2 0.00fF
C801 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00fF
C802 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C803 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C804 phi2 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.00fF
C805 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C806 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00fF
C807 mimtop2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00fF
C808 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.08fF
C809 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C810 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__nand2_1_0/a_113_47# 0.00fF
C811 sky130_fd_sc_hd__inv_1_4/Y VDD 0.15fF
C812 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_3/A 0.01fF
C813 sky130_fd_sc_hd__inv_1_4/Y clk 0.06fF
C814 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00fF
C815 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# phi2 0.00fF
C816 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00fF
C817 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A -0.00fF
C818 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00fF
C819 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C820 phi1 VSS 1.16fF
C821 sky130_fd_sc_hd__nand2_1_1/Y VSS 0.01fF
C822 sky130_fd_sc_hd__inv_1_2/Y VSS -0.27fF
C823 sky130_fd_sc_hd__inv_1_4/Y VSS 0.16fF
C824 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.02fF
C825 phi2 VSS 0.68fF
C826 sky130_fd_sc_hd__nand2_1_0/Y VSS 0.24fF
C827 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS 0.00fF
C828 mimtop1 VSS 0.27fF
C829 mimbot1 VSS -63.65fF
C830 mimtop2 VSS 13.83fF
C831 vcm VSS -781.24fF
C832 VDD VSS -1297.83fF
C833 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VSS 0.07fF
C834 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# VSS 0.05fF
C835 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# VSS 0.07fF
C836 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# VSS -0.01fF
C837 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# VSS 0.06fF
C838 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# VSS 0.05fF
C839 sky130_fd_sc_hd__inv_1_1/A VSS 0.32fF
C840 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# VSS 0.06fF
C841 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# VSS 0.08fF
C842 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# VSS 0.03fF
C843 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# VSS 0.10fF
C844 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# VSS 0.10fF
C845 sky130_fd_sc_hd__inv_1_0/A VSS 0.31fF
C846 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# VSS 0.06fF
C847 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# VSS 0.09fF
C848 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# VSS 0.03fF
C849 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# VSS 0.11fF
C850 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# VSS 0.11fF
C851 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VSS 0.07fF
C852 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# VSS 0.07fF
C853 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# VSS 0.08fF
C854 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# VSS 0.01fF
C855 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# VSS 0.09fF
C856 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# VSS 0.08fF
C857 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VSS 0.01fF
C858 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# VSS 0.02fF
C859 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# VSS 0.05fF
C860 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# VSS -0.01fF
C861 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# VSS 0.06fF
C862 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# VSS 0.04fF
C863 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VSS 0.06fF
C864 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# VSS 0.07fF
C865 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# VSS 0.10fF
C866 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# VSS 0.04fF
C867 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# VSS 0.10fF
C868 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# VSS 0.14fF
C869 sky130_fd_sc_hd__inv_1_3/Y VSS -1.49fF
C870 sky130_fd_sc_hd__buf_4_3/a_27_47# VSS 0.38fF
C871 sky130_fd_sc_hd__inv_1_3/A VSS 0.05fF
C872 sky130_fd_sc_hd__buf_4_2/a_27_47# VSS 0.30fF
C873 phi1_n VSS -0.59fF
C874 phi2_n VSS -0.56fF
C875 sky130_fd_sc_hd__buf_4_1/a_27_47# VSS 0.38fF
C876 sky130_fd_sc_hd__inv_1_2/A VSS 0.06fF
C877 sky130_fd_sc_hd__buf_4_0/a_27_47# VSS 0.29fF
C878 clk VSS 0.53fF
.ends

