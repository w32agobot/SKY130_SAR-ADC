VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO delay_macrocell
  CLASS BLOCK ;
  FOREIGN delay_macrocell ;
  ORIGIN 0.190 0.240 ;
  SIZE 9.500 BY 3.210 ;
  PIN in
    ANTENNAGATEAREA 4.880000 ;
    PORT
      LAYER li1 ;
        RECT -0.160 1.030 0.240 1.300 ;
    END
  END in
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 9.120 2.810 ;
        RECT 0.050 1.520 0.220 2.360 ;
        RECT 5.380 1.520 5.550 2.630 ;
        RECT 7.380 1.350 7.550 2.630 ;
        RECT 7.380 1.180 8.060 1.350 ;
        RECT 7.890 0.380 8.060 1.180 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.050 1.600 0.220 2.280 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.120 2.970 ;
        RECT 0.020 1.540 0.250 2.480 ;
    END
  END VPWR
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190 1.220 9.310 2.910 ;
    END
  END VPB
  PIN out
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.402600 ;
    PORT
      LAYER li1 ;
        RECT 6.340 1.520 6.510 2.360 ;
        RECT 7.040 1.010 7.210 1.340 ;
        RECT 6.340 0.380 6.510 0.890 ;
      LAYER mcon ;
        RECT 6.340 1.600 6.510 1.880 ;
        RECT 7.040 1.090 7.210 1.260 ;
        RECT 6.340 0.720 6.510 0.890 ;
      LAYER met1 ;
        RECT 6.310 1.240 6.540 2.030 ;
        RECT 6.980 1.240 7.270 1.290 ;
        RECT 6.310 1.100 9.120 1.240 ;
        RECT 6.310 0.660 6.540 1.100 ;
        RECT 6.980 1.060 7.270 1.100 ;
    END
  END out
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 8.230 1.350 8.400 2.360 ;
        RECT 8.230 1.180 8.880 1.350 ;
        RECT 0.050 0.380 0.220 0.840 ;
        RECT 5.380 0.090 5.550 0.840 ;
        RECT 8.710 0.090 8.880 1.180 ;
        RECT 0.000 -0.090 9.120 0.090 ;
      LAYER mcon ;
        RECT 0.050 0.460 0.220 0.760 ;
        RECT 0.140 -0.090 0.320 0.090 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT 0.020 0.240 0.250 0.820 ;
        RECT 0.000 -0.240 9.120 0.240 ;
      LAYER via ;
        RECT 1.920 -0.090 2.180 0.180 ;
        RECT 7.050 -0.050 7.330 0.220 ;
      LAYER met2 ;
        RECT 1.790 -0.090 2.380 0.360 ;
        RECT 6.880 -0.090 7.470 0.360 ;
      LAYER via2 ;
        RECT 1.920 -0.060 2.200 0.220 ;
        RECT 7.020 -0.050 7.360 0.270 ;
      LAYER met3 ;
        RECT 1.790 -0.090 2.380 0.360 ;
        RECT 6.880 -0.090 7.470 0.360 ;
      LAYER via3 ;
        RECT 1.920 -0.060 2.240 0.260 ;
        RECT 7.020 -0.050 7.360 0.270 ;
      LAYER met4 ;
        RECT 1.830 0.360 2.270 1.330 ;
        RECT 6.930 0.360 7.380 1.260 ;
        RECT 1.790 -0.090 2.380 0.360 ;
        RECT 6.880 -0.090 7.470 0.360 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.005 0.110 8.790 0.240 ;
        RECT 0.005 0.105 8.880 0.110 ;
        RECT 0.140 -0.090 0.320 0.105 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 4.340 1.290 4.510 2.360 ;
        RECT 4.900 1.520 5.070 2.360 ;
        RECT 5.860 1.520 6.030 2.360 ;
        RECT 6.820 1.520 6.990 2.360 ;
        RECT 7.720 1.520 7.920 2.360 ;
        RECT 8.710 1.520 8.880 2.360 ;
        RECT 4.340 1.010 4.940 1.290 ;
        RECT 4.340 0.380 4.510 1.010 ;
        RECT 4.900 0.380 5.070 0.840 ;
        RECT 5.860 0.380 6.030 0.840 ;
        RECT 6.820 0.380 6.990 0.840 ;
        RECT 7.410 0.380 7.580 0.840 ;
        RECT 8.370 0.380 8.540 0.840 ;
      LAYER mcon ;
        RECT 4.340 1.600 4.510 2.280 ;
        RECT 4.900 1.600 5.070 2.280 ;
        RECT 5.860 1.600 6.030 2.280 ;
        RECT 6.820 1.600 6.990 2.280 ;
        RECT 7.750 1.700 7.920 2.280 ;
        RECT 8.710 1.700 8.880 2.280 ;
        RECT 4.580 1.060 4.860 1.230 ;
        RECT 4.340 0.460 4.510 0.760 ;
        RECT 4.900 0.460 5.070 0.760 ;
        RECT 5.860 0.460 6.030 0.760 ;
        RECT 6.820 0.460 6.990 0.760 ;
        RECT 7.410 0.460 7.580 0.660 ;
        RECT 8.370 0.460 8.540 0.660 ;
      LAYER met1 ;
        RECT 4.310 1.290 4.540 2.340 ;
        RECT 4.870 2.000 5.100 2.340 ;
        RECT 5.830 2.170 8.910 2.340 ;
        RECT 5.830 2.000 6.060 2.170 ;
        RECT 4.870 1.810 6.060 2.000 ;
        RECT 4.870 1.540 5.100 1.810 ;
        RECT 5.830 1.540 6.060 1.810 ;
        RECT 6.790 1.540 7.020 2.170 ;
        RECT 7.720 1.640 7.950 2.170 ;
        RECT 8.680 1.640 8.910 2.170 ;
        RECT 4.310 1.010 4.940 1.290 ;
        RECT 4.310 0.400 4.540 1.010 ;
        RECT 4.870 0.690 5.100 0.820 ;
        RECT 5.830 0.690 6.060 0.820 ;
        RECT 4.870 0.520 6.060 0.690 ;
        RECT 6.790 0.540 7.020 0.820 ;
        RECT 7.380 0.540 7.610 0.720 ;
        RECT 8.340 0.540 8.570 0.720 ;
        RECT 6.790 0.520 8.570 0.540 ;
        RECT 4.870 0.400 5.100 0.520 ;
        RECT 5.830 0.400 8.570 0.520 ;
        RECT 5.830 0.380 7.480 0.400 ;
      LAYER via ;
        RECT 4.580 1.020 4.860 1.280 ;
      LAYER met2 ;
        RECT 4.490 1.010 4.940 1.290 ;
      LAYER via2 ;
        RECT 4.580 1.010 4.860 1.290 ;
      LAYER met3 ;
        RECT 0.270 0.680 8.940 2.480 ;
  END
END delay_macrocell
END LIBRARY

