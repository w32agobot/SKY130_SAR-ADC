* NGSPICE file created from adc_top.ext - technology: sky130A

.subckt adc_top_postlayout result_out[0] result_out[1] result_out[2] result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8] result_out[9]
+ result_out[10] result_out[11] result_out[12] result_out[13] result_out[14] result_out[15] VDD VSS conversion_finished_out rst_n start_conversion_in clk_vcm
+ inp_analog inn_analog
+ config_1_in[0] config_1_in[1] config_1_in[2] config_1_in[3] config_1_in[4] config_1_in[5] config_1_in[6] config_1_in[7] config_1_in[8] config_1_in[9]
+ config_1_in[10] config_1_in[11] config_1_in[12] config_1_in[13] config_1_in[14] config_1_in[15] 
+ config_2_in[0] config_2_in[1] config_2_in[2] config_2_in[3] config_2_in[4] config_2_in[5] config_2_in[6] config_2_in[7] config_2_in[8] config_2_in[9] 
+ config_2_in[10] config_2_in[11] config_2_in[12] config_2_in[13] config_2_in[14] config_2_in[15] 
+ dummypin[0] dummypin[10] dummypin[11] dummypin[12] dummypin[13] dummypin[14] dummypin[15] dummypin[1] dummypin[2] dummypin[3] dummypin[4] dummypin[5] 
+ dummypin[6] dummypin[7] dummypin[8] dummypin[9]  
R_D0 VSS a_11067_67279# 1e15 m=1
R_D1 VSS a_2012_33927# 1e15 m=1
R_D10 VSS a_6835_46823# 1e15 m=1
R_D100 VSS a_5915_35943# 1e15 m=1
R_D101 VSS a_12907_27023# 1e15 m=1
R_D102 VSS a_21187_29415# 1e15 m=1
R_D103 VSS a_12641_37684# 1e15 m=1
R_D104 VSS a_4191_33449# 1e15 m=1
R_D105 VSS a_12341_3311# 1e15 m=1
R_D106 VSS a_27535_30503# 1e15 m=1
R_D107 VSS a_1761_41935# 1e15 m=1
R_D108 VSS a_4891_47388# 1e15 m=1
R_D109 VSS a_12473_36341# 1e15 m=1
R_D11 VSS a_27535_30503# 1e15 m=1
R_D110 VSS a_3339_32463# 1e15 m=1
R_D111 VSS a_27535_30503# 1e15 m=1
R_D112 VSS a_11067_13095# 1e15 m=1
R_D113 VSS a_2099_59861# 1e15 m=1
R_D114 VSS a_5831_39189# 1e15 m=1
R_D115 VSS a_8491_57487# 1e15 m=1
R_Dsky130_fd_pr__diode_pw2nd_05v5116 VSS a_3668_56311# 1e15 m=1
R_D117 VSS a_15607_46805# 1e15 m=1
R_D118 VSS config_2_in[9] 1e15 m=1
R_D119 VSS a_2339_38129# 1e15 m=1
R_D12 VSS a_12621_36091# 1e15 m=1
R_D120 VSS a_10515_63143# 1e15 m=1
R_D121 VSS a_7571_29199# 1e15 m=1
R_D122 VSS a_1761_43567# 1e15 m=1
R_D123 VSS a_7479_54439# 1e15 m=1
R_D124 VSS a_4891_47388# 1e15 m=1
R_D125 VSS a_7841_12167# 1e15 m=1
R_D126 VSS a_8491_27023# 1e15 m=1
R_D127 VSS a_6835_46823# 1e15 m=1
R_D128 VSS config_1_in[11] 1e15 m=1
R_D129 VSS a_2004_42453# 1e15 m=1
R_D13 VSS a_1761_22895# 1e15 m=1
R_D130 VSS a_10055_58791# 1e15 m=1
R_D131 VSS a_3987_19623# 1e15 m=1
R_D132 VSS a_2419_48783# 1e15 m=1
R_D133 VSS a_11067_63143# 1e15 m=1
R_D134 VSS a_2143_15271# 1e15 m=1
R_D135 VSS a_4758_45369# 1e15 m=1
R_D136 VSS a_4443_46607# 1e15 m=1
R_D137 VSS a_7295_44647# 1e15 m=1
R_D138 VSS a_34482_29941# 1e15 m=1
R_D139 VSS a_1768_13103# 1e15 m=1
R_D14 VSS a_2840_66103# 1e15 m=1
R_D140 VSS config_2_in[5] 1e15 m=1
R_D141 VSS a_11067_67279# 1e15 m=1
R_D142 VSS a_12357_37999# 1e15 m=1
R_D143 VSS a_6095_44807# 1e15 m=1
R_D144 VSS a_2606_41079# 1e15 m=1
R_D145 VSS a_12516_7093# 1e15 m=1
R_D146 VSS a_8583_33551# 1e15 m=1
R_D147 VSS a_1761_37039# 1e15 m=1
R_D148 VSS a_7862_34025# 1e15 m=1
R_D149 VSS a_2775_46025# 1e15 m=1
R_D15 VSS config_2_in[8] 1e15 m=1
R_D150 VSS a_6559_59879# 1e15 m=1
R_D151 VSS a_5363_30503# 1e15 m=1
R_D152 VSS a_3339_43023# 1e15 m=1
R_D153 VSS a_1586_21959# 1e15 m=1
R_D154 VSS a_21371_50959# 1e15 m=1
R_D155 VSS a_3339_43023# 1e15 m=1
R_D156 VSS a_3987_19623# 1e15 m=1
R_D157 VSS a_12447_29199# 1e15 m=1
R_D158 VSS a_4482_57863# 1e15 m=1
R_D159 VSS a_27535_30503# 1e15 m=1
R_D16 VSS a_8531_70543# 1e15 m=1
R_D160 VSS a_15607_46805# 1e15 m=1
R_D161 VSS a_8123_56399# 1e15 m=1
R_D162 VSS a_12263_4391# 1e15 m=1
R_D163 VSS a_18979_30287# 1e15 m=1
R_D164 VSS a_11067_66191# 1e15 m=1
R_D165 VSS a_12907_27023# 1e15 m=1
R_D166 VSS a_2012_33927# 1e15 m=1
R_D167 VSS a_6831_63303# 1e15 m=1
R_D168 VSS a_2787_30503# 1e15 m=1
R_D169 VSS a_43267_31055# 1e15 m=1
R_D17 VSS a_1586_51335# 1e15 m=1
R_D170 VSS a_29927_29199# 1e15 m=1
R_D171 VSS a_11251_59879# 1e15 m=1
R_D172 VSS a_19807_28111# 1e15 m=1
R_D173 VSS config_2_in[14] 1e15 m=1
R_D174 VSS a_1586_51335# 1e15 m=1
R_D175 VSS a_5831_39189# 1e15 m=1
R_D176 VSS a_23395_32463# 1e15 m=1
R_D177 VSS a_15607_46805# 1e15 m=1
R_D178 VSS a_29927_29199# 1e15 m=1
R_D179 VSS a_12355_65103# 1e15 m=1
R_D18 VSS a_6559_59879# 1e15 m=1
R_D180 VSS a_12357_37999# 1e15 m=1
R_D181 VSS a_10515_63143# 1e15 m=1
R_D182 VSS a_6831_63303# 1e15 m=1
R_D183 VSS a_7479_54439# 1e15 m=1
R_D184 VSS a_1586_51335# 1e15 m=1
R_D185 VSS a_12357_37999# 1e15 m=1
R_D186 VSS a_6095_44807# 1e15 m=1
R_D187 VSS a_11067_13095# 1e15 m=1
R_D188 VSS a_1761_39215# 1e15 m=1
R_D189 VSS a_12641_37684# 1e15 m=1
R_D19 VSS a_4351_67279# 1e15 m=1
R_D190 VSS a_2235_30503# 1e15 m=1
R_D191 VSS a_23395_32463# 1e15 m=1
R_D192 VSS a_2606_41079# 1e15 m=1
R_D193 VSS a_2411_26133# 1e15 m=1
R_D194 VSS a_11067_13095# 1e15 m=1
R_D195 VSS a_5363_30503# 1e15 m=1
R_D196 VSS a_8583_33551# 1e15 m=1
R_D197 VSS a_4191_33449# 1e15 m=1
R_D198 VSS a_4891_47388# 1e15 m=1
R_D199 VSS a_12473_41781# 1e15 m=1
R_D2 VSS a_5363_30503# 1e15 m=1
R_D20 VSS a_2012_33927# 1e15 m=1
R_D200 VSS config_2_in[6] 1e15 m=1
R_D201 VSS a_2012_33927# 1e15 m=1
R_D202 VSS a_2411_26133# 1e15 m=1
R_D203 VSS a_18151_52263# 1e15 m=1
R_D204 VSS a_2143_15271# 1e15 m=1
R_D205 VSS a_4674_40277# 1e15 m=1
R_D206 VSS a_2606_41079# 1e15 m=1
R_D207 VSS a_21187_29415# 1e15 m=1
R_D208 VSS a_28547_51175# 1e15 m=1
R_D209 VSS a_22843_29415# 1e15 m=1
R_D21 VSS a_2787_32679# 1e15 m=1
R_D210 VSS a_4351_67279# 1e15 m=1
R_D211 VSS a_4443_46607# 1e15 m=1
R_D212 VSS a_1761_49007# 1e15 m=1
R_D213 VSS a_26523_29199# 1e15 m=1
R_D214 VSS a_16863_29415# 1e15 m=1
R_D215 VSS a_19967_41781# 1e15 m=1
R_D216 VSS a_12663_40871# 1e15 m=1
R_D217 VSS a_11067_46823# 1e15 m=1
R_D218 VSS a_3339_43023# 1e15 m=1
R_D219 VSS a_1586_51335# 1e15 m=1
R_D22 VSS a_5682_69367# 1e15 m=1
R_D220 VSS a_2840_66103# 1e15 m=1
R_D221 VSS a_12357_37999# 1e15 m=1
R_D222 VSS a_10055_58791# 1e15 m=1
R_D223 VSS a_15607_46805# 1e15 m=1
R_D224 VSS a_1689_10396# 1e15 m=1
R_D225 VSS a_6559_59663# 1e15 m=1
R_D226 VSS a_1586_18695# 1e15 m=1
R_D227 VSS a_29927_29199# 1e15 m=1
R_D228 VSS a_3987_19623# 1e15 m=1
R_D229 VSS a_20635_29415# 1e15 m=1
R_D23 VSS a_4339_64521# 1e15 m=1
R_D230 VSS a_1761_46287# 1e15 m=1
R_D231 VSS a_6559_59879# 1e15 m=1
R_D232 VSS a_2840_66103# 1e15 m=1
R_D233 VSS a_4674_40277# 1e15 m=1
R_D234 VSS a_7571_29199# 1e15 m=1
R_D235 VSS a_12447_29199# 1e15 m=1
R_D236 VSS a_19807_28111# 1e15 m=1
R_D237 VSS config_1_in[5] 1e15 m=1
R_D238 VSS a_11067_46823# 1e15 m=1
R_D239 VSS a_12907_27023# 1e15 m=1
R_D24 VSS a_4482_57863# 1e15 m=1
R_D240 VSS a_7939_30503# 1e15 m=1
R_D241 VSS a_6835_46823# 1e15 m=1
R_D242 VSS a_11067_13095# 1e15 m=1
R_D243 VSS a_2143_15271# 1e15 m=1
R_D244 VSS a_12381_43957# 1e15 m=1
R_D245 VSS a_25971_52263# 1e15 m=1
R_D246 VSS a_14831_50095# 1e15 m=1
R_D247 VSS a_20267_30503# 1e15 m=1
R_D248 VSS a_20359_29199# 1e15 m=1
R_D249 VSS a_3987_19623# 1e15 m=1
R_D25 VSS a_11067_13095# 1e15 m=1
R_D250 VSS a_12869_2741# 1e15 m=1
R_D251 VSS a_2787_30503# 1e15 m=1
R_D252 VSS a_2872_44111# 1e15 m=1
R_D253 VSS a_8491_41383# 1e15 m=1
R_D254 VSS a_4674_40277# 1e15 m=1
R_D255 VSS a_5682_69367# 1e15 m=1
R_D256 VSS a_12663_40871# 1e15 m=1
R_D257 VSS a_4891_47388# 1e15 m=1
R_D258 VSS a_4482_57863# 1e15 m=1
R_D259 VSS a_29927_29199# 1e15 m=1
R_D26 VSS a_24959_30503# 1e15 m=1
R_D260 VSS a_3339_32463# 1e15 m=1
R_D261 VSS a_2840_66103# 1e15 m=1
R_D262 VSS a_12907_27023# 1e15 m=1
R_D263 VSS a_6095_44807# 1e15 m=1
R_D264 VSS a_3339_43023# 1e15 m=1
R_D265 VSS a_20635_29415# 1e15 m=1
R_D266 VSS a_1770_14441# 1e15 m=1
R_D267 VSS a_22291_29415# 1e15 m=1
R_D268 VSS a_8491_41383# 1e15 m=1
R_D269 VSS a_12516_7093# 1e15 m=1
R_D27 VSS a_1768_13103# 1e15 m=1
R_D270 VSS a_13097_36367# 1e15 m=1
R_D271 VSS a_1761_52815# 1e15 m=1
R_D272 VSS a_1586_21959# 1e15 m=1
R_D273 VSS a_4674_40277# 1e15 m=1
R_D274 VSS a_3987_19623# 1e15 m=1
R_D275 VSS a_2606_41079# 1e15 m=1
R_D276 VSS config_1_in[10] 1e15 m=1
R_D277 VSS a_7479_54439# 1e15 m=1
R_D278 VSS a_3339_30503# 1e15 m=1
R_D279 VSS a_6095_44807# 1e15 m=1
R_D28 VSS a_4215_51157# 1e15 m=1
R_D280 VSS a_4758_45369# 1e15 m=1
R_D281 VSS a_18611_52047# 1e15 m=1
R_D282 VSS a_2419_48783# 1e15 m=1
R_D283 VSS a_4891_47388# 1e15 m=1
R_D284 VSS a_2235_30503# 1e15 m=1
R_D285 VSS a_8583_33551# 1e15 m=1
R_D286 VSS a_5682_69367# 1e15 m=1
R_D287 VSS a_6831_63303# 1e15 m=1
R_D288 VSS a_11619_56615# 1e15 m=1
R_D289 VSS a_2959_47113# 1e15 m=1
R_D29 VSS a_4191_33449# 1e15 m=1
R_D290 VSS a_4215_51157# 1e15 m=1
R_D291 VSS a_13067_38517# 1e15 m=1
R_D292 VSS a_12899_2767# 1e15 m=1
R_D293 VSS a_4811_34855# 1e15 m=1
R_D294 VSS a_2339_38129# 1e15 m=1
R_D295 VSS a_20359_29199# 1e15 m=1
R_D296 VSS a_4891_47388# 1e15 m=1
R_D297 VSS a_2959_47113# 1e15 m=1
R_D298 VSS a_3987_19623# 1e15 m=1
R_D299 VSS a_29927_29199# 1e15 m=1
R_D3 VSS a_12663_35431# 1e15 m=1
R_D30 VSS a_4351_67279# 1e15 m=1
R_D300 VSS a_4119_70741# 1e15 m=1
R_D301 VSS a_2411_26133# 1e15 m=1
R_D302 VSS a_6831_63303# 1e15 m=1
R_D303 VSS a_4215_51157# 1e15 m=1
R_D304 VSS a_2411_26133# 1e15 m=1
R_D305 VSS a_5915_35943# 1e15 m=1
R_D306 VSS a_1689_10396# 1e15 m=1
R_D307 VSS a_4443_46607# 1e15 m=1
R_D308 VSS a_4215_51157# 1e15 m=1
R_D309 VSS a_16863_29415# 1e15 m=1
R_D31 VSS a_4119_70741# 1e15 m=1
R_D310 VSS a_4674_40277# 1e15 m=1
R_D311 VSS rst_n 1e15 m=1
R_D312 VSS a_3339_32463# 1e15 m=1
R_D313 VSS a_1586_21959# 1e15 m=1
R_D314 VSS a_3339_43023# 1e15 m=1
R_D315 VSS a_1586_18695# 1e15 m=1
R_D316 VSS a_18979_30287# 1e15 m=1
R_D317 VSS a_2419_48783# 1e15 m=1
R_D318 VSS config_1_in[1] 1e15 m=1
R_D319 VSS a_2872_44111# 1e15 m=1
R_D32 VSS a_4191_33449# 1e15 m=1
R_D320 VSS a_2143_15271# 1e15 m=1
R_D321 VSS a_12725_44527# 1e15 m=1
R_D322 VSS a_26523_29199# 1e15 m=1
R_D323 VSS a_1761_50639# 1e15 m=1
R_D324 VSS a_1950_59887# 1e15 m=1
R_D325 VSS a_7571_26151# 1e15 m=1
R_D326 VSS a_22843_29415# 1e15 m=1
R_D327 VSS config_2_in[1] 1e15 m=1
R_D328 VSS a_4811_34855# 1e15 m=1
R_D329 VSS a_5363_30503# 1e15 m=1
R_D33 VSS a_13123_38231# 1e15 m=1
R_D330 VSS a_10975_66407# 1e15 m=1
R_D331 VSS a_4351_67279# 1e15 m=1
R_D332 VSS a_10055_58791# 1e15 m=1
R_D333 VSS a_2872_44111# 1e15 m=1
R_D334 VSS a_3987_19623# 1e15 m=1
R_D335 VSS a_7479_54439# 1e15 m=1
R_D336 VSS a_2959_47113# 1e15 m=1
R_D337 VSS a_2004_42453# 1e15 m=1
R_D338 VSS a_11067_46823# 1e15 m=1
R_D339 VSS a_11067_21583# 1e15 m=1
R_D34 VSS a_4811_34855# 1e15 m=1
R_D340 VSS a_18703_29199# 1e15 m=1
R_D341 VSS a_11067_46823# 1e15 m=1
R_D342 VSS a_4215_51157# 1e15 m=1
R_D343 VSS a_3247_20495# 1e15 m=1
R_D344 VSS a_1950_59887# 1e15 m=1
R_D345 VSS a_19807_28111# 1e15 m=1
R_D346 VSS a_4339_64521# 1e15 m=1
R_D347 VSS a_11067_67279# 1e15 m=1
R_D348 VSS a_4351_67279# 1e15 m=1
R_D349 VSS a_38115_52263# 1e15 m=1
R_D35 VSS a_4119_70741# 1e15 m=1
R_D350 VSS a_20359_29199# 1e15 m=1
R_D351 VSS a_2606_41079# 1e15 m=1
R_D352 VSS a_11067_66191# 1e15 m=1
R_D353 VSS a_14287_51175# 1e15 m=1
R_D354 VSS a_4674_40277# 1e15 m=1
R_D355 VSS a_4339_64521# 1e15 m=1
R_D356 VSS a_1770_14441# 1e15 m=1
R_D357 VSS a_7939_30503# 1e15 m=1
R_D358 VSS a_3247_20495# 1e15 m=1
R_D359 VSS a_10687_52553# 1e15 m=1
R_D36 VSS a_4443_46607# 1e15 m=1
R_D360 VSS a_2411_26133# 1e15 m=1
R_D361 VSS a_4482_57863# 1e15 m=1
R_D362 VSS a_6831_63303# 1e15 m=1
R_D363 VSS a_4891_47388# 1e15 m=1
R_D364 VSS a_1768_16367# 1e15 m=1
R_D365 VSS a_2959_47113# 1e15 m=1
R_D366 VSS a_3339_30503# 1e15 m=1
R_D367 VSS a_2840_66103# 1e15 m=1
R_D368 VSS a_12869_2741# 1e15 m=1
R_D369 VSS a_2099_59861# 1e15 m=1
R_D37 VSS a_8295_47388# 1e15 m=1
R_D370 VSS a_5682_69367# 1e15 m=1
R_D371 VSS a_4811_34855# 1e15 m=1
R_D372 VSS a_13643_28327# 1e15 m=1
R_D373 VSS a_4215_51157# 1e15 m=1
R_D374 VSS a_7939_30503# 1e15 m=1
R_D375 VSS a_3339_30503# 1e15 m=1
R_D376 VSS a_6835_46823# 1e15 m=1
R_D377 VSS a_6559_22671# 1e15 m=1
R_D378 VSS a_6835_46823# 1e15 m=1
R_D379 VSS a_8531_70543# 1e15 m=1
R_D38 VSS a_7571_29199# 1e15 m=1
R_D380 VSS a_1761_50639# 1e15 m=1
R_D381 VSS a_2840_66103# 1e15 m=1
R_D382 VSS a_2021_17973# 1e15 m=1
R_D383 VSS a_2787_32679# 1e15 m=1
R_D384 VSS a_6559_59879# 1e15 m=1
R_D385 VSS a_20635_29415# 1e15 m=1
R_D386 VSS a_10515_23975# 1e15 m=1
R_D387 VSS a_2787_32679# 1e15 m=1
R_D388 VSS a_1586_18695# 1e15 m=1
R_D389 VSS a_1950_59887# 1e15 m=1
R_D39 VSS a_11067_47695# 1e15 m=1
R_D390 VSS a_18979_30287# 1e15 m=1
R_D391 VSS a_12907_27023# 1e15 m=1
R_D392 VSS a_5915_35943# 1e15 m=1
R_D393 VSS a_2419_48783# 1e15 m=1
R_D394 VSS a_4443_46607# 1e15 m=1
R_D395 VSS config_2_in[13] 1e15 m=1
R_D396 VSS a_19807_28111# 1e15 m=1
R_D397 VSS a_4758_45369# 1e15 m=1
R_D398 VSS a_20359_29199# 1e15 m=1
R_D399 VSS a_5831_39189# 1e15 m=1
R_D4 VSS a_1586_18695# 1e15 m=1
R_D40 VSS a_25787_28327# 1e15 m=1
R_D400 VSS a_3247_20495# 1e15 m=1
R_D401 VSS a_3339_43023# 1e15 m=1
R_D402 VSS a_5363_30503# 1e15 m=1
R_D403 VSS a_3339_43023# 1e15 m=1
R_D404 VSS a_4339_64521# 1e15 m=1
R_D405 VSS a_12907_27023# 1e15 m=1
R_D406 VSS a_11619_56615# 1e15 m=1
R_D407 VSS a_4191_33449# 1e15 m=1
R_D408 VSS a_7295_44647# 1e15 m=1
R_D409 VSS a_13669_35253# 1e15 m=1
R_D41 VSS a_3668_56311# 1e15 m=1
R_D410 VSS a_29927_29199# 1e15 m=1
R_D411 VSS config_1_in[3] 1e15 m=1
R_D412 VSS a_27535_30503# 1e15 m=1
R_D413 VSS a_6831_63303# 1e15 m=1
R_D414 VSS a_7862_34025# 1e15 m=1
R_D415 VSS a_8295_47388# 1e15 m=1
R_D416 VSS a_10515_63143# 1e15 m=1
R_D417 VSS a_12357_37999# 1e15 m=1
R_D418 VSS a_27535_30503# 1e15 m=1
R_D419 VSS a_11067_46823# 1e15 m=1
R_D42 VSS a_1761_31055# 1e15 m=1
R_D420 VSS a_5682_69367# 1e15 m=1
R_D421 VSS a_6831_63303# 1e15 m=1
R_D422 VSS a_19807_28111# 1e15 m=1
R_D423 VSS config_2_in[3] 1e15 m=1
R_D424 VSS a_2606_41079# 1e15 m=1
R_D425 VSS a_5915_35943# 1e15 m=1
R_D426 VSS a_13669_37429# 1e15 m=1
R_D427 VSS a_19807_28111# 1e15 m=1
R_D428 VSS a_11067_63143# 1e15 m=1
R_D429 VSS a_10515_63143# 1e15 m=1
R_D43 VSS a_20635_29415# 1e15 m=1
R_D430 VSS a_20359_29199# 1e15 m=1
R_D431 VSS config_1_in[0] 1e15 m=1
R_D432 VSS inp_analog 1e15 m=1
R_D433 VSS a_7571_29199# 1e15 m=1
R_D434 VSS a_7295_44647# 1e15 m=1
R_D435 VSS a_14831_50095# 1e15 m=1
R_D436 VSS a_7841_12167# 1e15 m=1
R_D437 VSS config_2_in[12] 1e15 m=1
R_D438 VSS a_5831_39189# 1e15 m=1
R_D439 VSS a_22015_28111# 1e15 m=1
R_D44 VSS a_1950_59887# 1e15 m=1
R_D440 VSS a_19807_28111# 1e15 m=1
R_D441 VSS a_4811_34855# 1e15 m=1
R_D442 VSS a_4351_67279# 1e15 m=1
R_D443 VSS a_4191_33449# 1e15 m=1
R_D444 VSS a_13716_43047# 1e15 m=1
R_D445 VSS a_17599_52263# 1e15 m=1
R_D446 VSS a_26523_28111# 1e15 m=1
R_D447 VSS a_2012_33927# 1e15 m=1
R_D448 VSS a_12516_7093# 1e15 m=1
R_D449 VSS a_3247_20495# 1e15 m=1
R_D45 VSS a_10680_52245# 1e15 m=1
R_D450 VSS a_12473_36341# 1e15 m=1
R_D451 VSS a_1761_32143# 1e15 m=1
R_D452 VSS a_2339_38129# 1e15 m=1
R_D453 VSS a_2143_15271# 1e15 m=1
R_D454 VSS config_1_in[4] 1e15 m=1
R_D455 VSS a_3339_43023# 1e15 m=1
R_D456 VSS a_12725_44527# 1e15 m=1
R_D457 VSS config_2_in[11] 1e15 m=1
R_D458 VSS a_1586_51335# 1e15 m=1
R_D459 VSS a_5915_35943# 1e15 m=1
R_D46 VSS a_26523_28111# 1e15 m=1
R_D460 VSS a_12725_44527# 1e15 m=1
R_D461 VSS a_7571_29199# 1e15 m=1
R_D462 VSS a_4443_46607# 1e15 m=1
R_D463 VSS a_1586_18695# 1e15 m=1
R_D464 VSS a_2606_41079# 1e15 m=1
R_D465 VSS a_20359_29199# 1e15 m=1
R_D466 VSS config_1_in[12] 1e15 m=1
R_D467 VSS a_6467_55527# 1e15 m=1
R_D468 VSS a_2787_30503# 1e15 m=1
R_D469 VSS a_12869_2741# 1e15 m=1
R_D47 VSS a_2235_30503# 1e15 m=1
R_D470 VSS a_2143_15271# 1e15 m=1
R_D471 VSS a_5831_39189# 1e15 m=1
R_D472 VSS a_12907_27023# 1e15 m=1
R_D473 VSS a_4339_64521# 1e15 m=1
R_D474 VSS a_12899_3855# 1e15 m=1
R_D475 VSS a_2339_38129# 1e15 m=1
R_D476 VSS a_10515_63143# 1e15 m=1
R_D477 VSS a_1950_59887# 1e15 m=1
R_D478 VSS a_18979_30287# 1e15 m=1
R_D479 VSS a_6559_22671# 1e15 m=1
R_D48 VSS a_8123_56399# 1e15 m=1
R_D480 VSS config_2_in[0] 1e15 m=1
R_D481 VSS a_2004_42453# 1e15 m=1
R_D482 VSS a_11067_21583# 1e15 m=1
R_D483 VSS a_6559_59879# 1e15 m=1
R_D484 VSS a_2235_30503# 1e15 m=1
R_D485 VSS a_8491_41383# 1e15 m=1
R_D486 VSS a_1689_10396# 1e15 m=1
R_D487 VSS a_7571_26151# 1e15 m=1
R_D488 VSS a_1586_18695# 1e15 m=1
R_D489 VSS a_12381_35836# 1e15 m=1
R_D49 VSS a_20267_30503# 1e15 m=1
R_D490 VSS a_2012_33927# 1e15 m=1
R_D491 VSS config_2_in[4] 1e15 m=1
R_D492 VSS a_11067_46823# 1e15 m=1
R_D493 VSS a_19807_28111# 1e15 m=1
R_D494 VSS a_2004_42453# 1e15 m=1
R_D495 VSS a_3339_43023# 1e15 m=1
R_D496 VSS a_13669_35253# 1e15 m=1
R_D497 VSS a_13716_43047# 1e15 m=1
R_D498 VSS a_5682_69367# 1e15 m=1
R_D499 VSS a_2787_32679# 1e15 m=1
R_D5 VSS a_23395_32463# 1e15 m=1
R_D50 VSS a_18979_30287# 1e15 m=1
R_D500 VSS a_4811_34855# 1e15 m=1
R_D501 VSS a_14831_50095# 1e15 m=1
R_D502 VSS a_4215_51157# 1e15 m=1
R_D503 VSS a_11067_46823# 1e15 m=1
R_D504 VSS a_2787_30503# 1e15 m=1
R_D505 VSS a_3668_56311# 1e15 m=1
R_D506 VSS config_2_in[15] 1e15 m=1
R_D507 VSS a_18703_29199# 1e15 m=1
R_D508 VSS a_13183_52047# 1e15 m=1
R_D509 VSS a_4119_70741# 1e15 m=1
R_D51 VSS config_1_in[15] 1e15 m=1
R_D510 VSS a_11067_47695# 1e15 m=1
R_D511 VSS a_4119_70741# 1e15 m=1
R_D512 VSS a_16863_29415# 1e15 m=1
R_D513 VSS a_2021_22325# 1e15 m=1
R_D514 VSS a_13005_35823# 1e15 m=1
R_D515 VSS a_10055_58791# 1e15 m=1
R_D516 VSS a_1761_52815# 1e15 m=1
R_D517 VSS a_22015_28111# 1e15 m=1
R_D518 VSS a_1803_19087# 1e15 m=1
R_D519 VSS a_10680_52245# 1e15 m=1
R_D52 VSS a_13643_28327# 1e15 m=1
R_D520 VSS a_6467_55527# 1e15 m=1
R_D521 VSS a_10975_66407# 1e15 m=1
R_D522 VSS a_18703_29199# 1e15 m=1
R_D523 VSS a_1689_10396# 1e15 m=1
R_D524 VSS a_2872_44111# 1e15 m=1
R_D525 VSS a_13909_39747# 1e15 m=1
R_D526 VSS a_2012_33927# 1e15 m=1
R_D527 VSS a_1768_16367# 1e15 m=1
R_D528 VSS a_22291_29415# 1e15 m=1
R_D529 VSS a_15607_46805# 1e15 m=1
R_D53 VSS a_25419_50959# 1e15 m=1
R_D530 VSS a_26523_29199# 1e15 m=1
R_D531 VSS a_2004_42453# 1e15 m=1
R_D532 VSS a_12381_35836# 1e15 m=1
R_D533 VSS a_11619_56615# 1e15 m=1
R_D534 VSS a_14831_50095# 1e15 m=1
R_D535 VSS a_34251_52263# 1e15 m=1
R_D536 VSS a_3339_43023# 1e15 m=1
R_D537 VSS a_2775_46025# 1e15 m=1
R_D538 VSS a_5363_30503# 1e15 m=1
R_D539 VSS a_3339_30503# 1e15 m=1
R_D54 VSS a_6559_59663# 1e15 m=1
R_D540 VSS a_11067_67279# 1e15 m=1
R_D541 VSS a_2099_59861# 1e15 m=1
R_D542 VSS a_10975_66407# 1e15 m=1
R_D543 VSS a_2787_32679# 1e15 m=1
R_D544 VSS a_6467_55527# 1e15 m=1
R_D545 VSS a_8531_70543# 1e15 m=1
R_D546 VSS a_3339_43023# 1e15 m=1
R_D547 VSS a_4674_40277# 1e15 m=1
R_D548 VSS a_41872_29423# 1e15 m=1
R_D549 VSS a_8583_33551# 1e15 m=1
R_D55 VSS a_12473_41781# 1e15 m=1
R_D550 VSS a_20635_29415# 1e15 m=1
R_D551 VSS a_2235_30503# 1e15 m=1
R_D552 VSS a_7862_34025# 1e15 m=1
R_D553 VSS a_4215_51157# 1e15 m=1
R_D554 VSS a_41427_52263# 1e15 m=1
R_D555 VSS a_26523_28111# 1e15 m=1
R_D556 VSS a_1689_10396# 1e15 m=1
R_D557 VSS a_2191_68565# 1e15 m=1
R_D558 VSS a_7841_12167# 1e15 m=1
R_D559 VSS config_1_in[7] 1e15 m=1
R_D56 VSS a_10515_22671# 1e15 m=1
R_D560 VSS a_11067_23759# 1e15 m=1
R_D561 VSS a_4119_70741# 1e15 m=1
R_D562 VSS a_27535_30503# 1e15 m=1
R_D563 VSS a_10515_63143# 1e15 m=1
R_D564 VSS clk_vcm 1e15 m=1
R_D565 VSS a_3339_32463# 1e15 m=1
R_D566 VSS a_4811_34855# 1e15 m=1
R_D567 VSS a_20635_29415# 1e15 m=1
R_D568 VSS a_20359_29199# 1e15 m=1
R_D569 VSS a_13643_28327# 1e15 m=1
R_D57 VSS a_11067_13095# 1e15 m=1
R_D570 VSS config_1_in[14] 1e15 m=1
R_D571 VSS a_2959_47113# 1e15 m=1
R_D572 VSS a_4811_34855# 1e15 m=1
R_D573 VSS a_1586_21959# 1e15 m=1
R_D574 VSS a_12473_42869# 1e15 m=1
R_D575 VSS a_15607_46805# 1e15 m=1
R_D576 VSS a_10515_23975# 1e15 m=1
R_D577 VSS a_20635_29415# 1e15 m=1
R_D578 VSS a_7571_29199# 1e15 m=1
R_D579 VSS a_1761_47919# 1e15 m=1
R_D58 VSS a_2787_30503# 1e15 m=1
R_D580 VSS a_10687_52553# 1e15 m=1
R_D581 VSS a_10515_22671# 1e15 m=1
R_D582 VSS a_7939_30503# 1e15 m=1
R_D583 VSS a_7571_26151# 1e15 m=1
R_D584 VSS a_38557_32143# 1e15 m=1
R_D585 VSS a_7841_12167# 1e15 m=1
R_D586 VSS a_41427_52263# 1e15 m=1
R_D587 VSS a_8583_33551# 1e15 m=1
R_D588 VSS a_1689_10396# 1e15 m=1
R_D589 VSS a_2099_59861# 1e15 m=1
R_D59 VSS a_10515_63143# 1e15 m=1
R_D590 VSS a_12641_37684# 1e15 m=1
R_D591 VSS a_3247_20495# 1e15 m=1
R_D592 VSS a_20267_30503# 1e15 m=1
R_D593 VSS a_4482_57863# 1e15 m=1
R_D594 VSS a_1586_51335# 1e15 m=1
R_D595 VSS a_2411_26133# 1e15 m=1
R_D596 VSS a_12725_44527# 1e15 m=1
R_D597 VSS a_12355_65103# 1e15 m=1
R_D598 VSS a_12447_29199# 1e15 m=1
R_D599 VSS a_5915_35943# 1e15 m=1
R_D6 VSS a_4443_46607# 1e15 m=1
R_D60 VSS a_2840_66103# 1e15 m=1
R_D600 VSS a_6559_22671# 1e15 m=1
R_D601 VSS a_1586_18695# 1e15 m=1
R_D602 VSS a_6831_63303# 1e15 m=1
R_D603 VSS a_20359_29199# 1e15 m=1
R_D604 VSS a_4443_46607# 1e15 m=1
R_D605 VSS a_2012_33927# 1e15 m=1
R_D606 VSS a_2235_30503# 1e15 m=1
R_D607 VSS a_12907_56399# 1e15 m=1
R_D608 VSS a_14831_50095# 1e15 m=1
R_D609 VSS a_12663_35431# 1e15 m=1
R_D61 VSS a_4758_45369# 1e15 m=1
R_D610 VSS a_1803_20719# 1e15 m=1
R_D611 VSS a_16863_29415# 1e15 m=1
R_D612 VSS a_10055_58791# 1e15 m=1
R_D613 VSS a_4482_57863# 1e15 m=1
R_D614 VSS a_5363_30503# 1e15 m=1
R_D615 VSS a_11067_67279# 1e15 m=1
R_D616 VSS a_2339_38129# 1e15 m=1
R_D617 VSS a_12907_27023# 1e15 m=1
R_D618 VSS a_11619_3303# 1e15 m=1
R_D619 VSS a_12473_37429# 1e15 m=1
R_D62 VSS a_11067_13095# 1e15 m=1
R_D620 VSS a_12447_29199# 1e15 m=1
R_D621 VSS a_22291_29415# 1e15 m=1
R_D622 VSS a_2775_46025# 1e15 m=1
R_D623 VSS a_2021_17973# 1e15 m=1
R_D624 VSS a_2959_47113# 1e15 m=1
R_D625 VSS a_4339_64521# 1e15 m=1
R_D626 VSS a_6831_63303# 1e15 m=1
R_D627 VSS a_3339_30503# 1e15 m=1
R_D628 VSS a_9503_26151# 1e15 m=1
R_D629 VSS a_2235_30503# 1e15 m=1
R_D63 VSS a_7571_29199# 1e15 m=1
R_D630 VSS a_2191_68565# 1e15 m=1
R_D631 VSS a_14831_50095# 1e15 m=1
R_D632 VSS a_2959_47113# 1e15 m=1
R_D633 VSS a_18979_30287# 1e15 m=1
R_D634 VSS a_12907_27023# 1e15 m=1
R_D635 VSS a_7862_34025# 1e15 m=1
R_D636 VSS a_5682_69367# 1e15 m=1
R_D637 VSS a_1761_52815# 1e15 m=1
R_D638 VSS a_15607_46805# 1e15 m=1
R_D639 VSS a_5915_30287# 1e15 m=1
R_D64 VSS a_11067_67279# 1e15 m=1
R_D640 VSS a_2012_33927# 1e15 m=1
R_D641 VSS a_2419_48783# 1e15 m=1
R_D642 VSS a_3247_20495# 1e15 m=1
R_D643 VSS a_1761_35407# 1e15 m=1
R_D644 VSS a_1761_52815# 1e15 m=1
R_D645 VSS a_2775_46025# 1e15 m=1
R_D646 VSS a_1586_51335# 1e15 m=1
R_D647 VSS a_2606_41079# 1e15 m=1
R_D648 VSS a_11067_13095# 1e15 m=1
R_D649 VSS a_12355_15055# 1e15 m=1
R_D65 VSS a_12899_3311# 1e15 m=1
R_D650 VSS a_1761_30511# 1e15 m=1
R_D651 VSS a_9135_27239# 1e15 m=1
R_D652 VSS config_1_in[2] 1e15 m=1
R_D653 VSS a_13643_28327# 1e15 m=1
R_D654 VSS a_1770_14441# 1e15 m=1
R_D655 VSS a_2606_41079# 1e15 m=1
R_D656 VSS a_11067_47695# 1e15 m=1
R_D657 VSS a_26523_28111# 1e15 m=1
R_D658 VSS a_6559_59663# 1e15 m=1
R_D659 VSS a_23395_52047# 1e15 m=1
R_D66 VSS a_18979_30287# 1e15 m=1
R_D660 VSS a_11067_46823# 1e15 m=1
R_D661 VSS a_20359_29199# 1e15 m=1
R_D662 VSS a_19807_28111# 1e15 m=1
R_D663 VSS a_6095_44807# 1e15 m=1
R_D664 VSS a_7939_30503# 1e15 m=1
R_D665 VSS a_20635_29415# 1e15 m=1
R_D666 VSS a_4351_67279# 1e15 m=1
R_D667 VSS a_1586_21959# 1e15 m=1
R_D668 VSS a_3339_32463# 1e15 m=1
R_D669 VSS a_6559_22671# 1e15 m=1
R_D67 VSS a_2143_15271# 1e15 m=1
R_D670 VSS a_7295_44647# 1e15 m=1
R_D671 VSS a_11067_67279# 1e15 m=1
R_D672 VSS a_12473_37429# 1e15 m=1
R_D673 VSS a_2012_33927# 1e15 m=1
R_D674 VSS a_1761_40847# 1e15 m=1
R_D675 VSS a_7841_12167# 1e15 m=1
R_D676 VSS a_11067_13095# 1e15 m=1
R_D677 VSS a_12355_65103# 1e15 m=1
R_D678 VSS a_13643_28327# 1e15 m=1
R_D679 VSS a_3247_20495# 1e15 m=1
R_D68 VSS a_2775_46025# 1e15 m=1
R_D680 VSS a_11803_55311# 1e15 m=1
R_D681 VSS a_4339_64521# 1e15 m=1
R_D682 VSS a_20635_29415# 1e15 m=1
R_D683 VSS a_1689_10396# 1e15 m=1
R_D684 VSS config_1_in[9] 1e15 m=1
R_D685 VSS a_4443_46607# 1e15 m=1
R_D686 VSS a_2235_30503# 1e15 m=1
R_D687 VSS a_8531_70543# 1e15 m=1
R_D688 VSS a_3668_56311# 1e15 m=1
R_D689 VSS a_3668_56311# 1e15 m=1
R_D69 VSS a_8583_33551# 1e15 m=1
R_D690 VSS a_6467_55527# 1e15 m=1
R_D691 VSS config_1_in[8] 1e15 m=1
R_D692 VSS a_22843_29415# 1e15 m=1
R_D693 VSS a_7571_26151# 1e15 m=1
R_D694 VSS a_6559_22671# 1e15 m=1
R_D695 VSS a_6831_63303# 1e15 m=1
R_D696 VSS a_1761_25071# 1e15 m=1
R_D697 VSS a_10515_63143# 1e15 m=1
R_D698 VSS a_1586_18695# 1e15 m=1
R_D699 VSS a_5915_30287# 1e15 m=1
R_D7 VSS config_2_in[2] 1e15 m=1
R_D70 VSS a_2235_30503# 1e15 m=1
R_D700 VSS a_26523_29199# 1e15 m=1
R_D701 VSS a_11067_46823# 1e15 m=1
R_D702 VSS a_11067_66191# 1e15 m=1
R_D703 VSS a_5831_39189# 1e15 m=1
R_D704 VSS a_4758_45369# 1e15 m=1
R_D705 VSS a_13669_37429# 1e15 m=1
R_D706 VSS a_2787_32679# 1e15 m=1
R_D707 VSS a_6559_22671# 1e15 m=1
R_D708 VSS a_5915_30287# 1e15 m=1
R_D709 VSS a_2959_47113# 1e15 m=1
R_D71 VSS a_2606_41079# 1e15 m=1
R_D710 VSS a_1689_10396# 1e15 m=1
R_D711 VSS a_12447_29199# 1e15 m=1
R_D712 VSS a_2411_26133# 1e15 m=1
R_D713 VSS a_12447_29199# 1e15 m=1
R_D714 VSS a_20635_29415# 1e15 m=1
R_D715 VSS a_5915_30287# 1e15 m=1
R_D716 VSS a_22015_28111# 1e15 m=1
R_D717 VSS a_1586_21959# 1e15 m=1
R_D718 VSS a_7295_44647# 1e15 m=1
R_D719 VSS a_2191_68565# 1e15 m=1
R_D72 VSS a_18979_30287# 1e15 m=1
R_D720 VSS a_7939_30503# 1e15 m=1
R_D721 VSS a_1761_22895# 1e15 m=1
R_D722 VSS a_23395_32463# 1e15 m=1
R_D723 VSS a_19807_28111# 1e15 m=1
R_D724 VSS a_1761_34319# 1e15 m=1
R_D725 VSS a_22015_28111# 1e15 m=1
R_D726 VSS a_7479_54439# 1e15 m=1
R_D727 VSS a_2099_59861# 1e15 m=1
R_D728 VSS a_1761_27791# 1e15 m=1
R_D729 VSS config_1_in[13] 1e15 m=1
R_D73 VSS a_12447_29199# 1e15 m=1
R_D730 VSS a_7862_34025# 1e15 m=1
R_D731 VSS a_3668_56311# 1e15 m=1
R_D732 VSS a_34482_29941# 1e15 m=1
R_D733 VSS a_8491_41383# 1e15 m=1
R_D734 VSS a_8123_56399# 1e15 m=1
R_D735 VSS a_1586_18695# 1e15 m=1
R_D736 VSS a_22291_29415# 1e15 m=1
R_D737 VSS a_11067_66191# 1e15 m=1
R_D738 VSS a_13097_36367# 1e15 m=1
R_D739 VSS a_8583_33551# 1e15 m=1
R_D74 VSS a_4351_67279# 1e15 m=1
R_D740 VSS a_1768_13103# 1e15 m=1
R_D741 VSS a_21187_29415# 1e15 m=1
R_D742 VSS a_6559_59663# 1e15 m=1
R_D743 VSS a_10515_22671# 1e15 m=1
R_D744 VSS a_10680_52245# 1e15 m=1
R_D745 VSS a_1761_25071# 1e15 m=1
R_D746 VSS a_10515_63143# 1e15 m=1
R_D747 VSS a_26523_29199# 1e15 m=1
R_D748 VSS a_11067_46823# 1e15 m=1
R_D749 VSS a_2143_15271# 1e15 m=1
R_D75 VSS a_2419_48783# 1e15 m=1
R_D750 VSS a_24959_30503# 1e15 m=1
R_D751 VSS a_7571_29199# 1e15 m=1
R_D752 VSS a_6559_22671# 1e15 m=1
R_D753 VSS a_4351_67279# 1e15 m=1
R_D754 VSS a_17507_52047# 1e15 m=1
R_D755 VSS a_4443_46607# 1e15 m=1
R_D756 VSS a_6835_46823# 1e15 m=1
R_D757 VSS a_4443_46607# 1e15 m=1
R_D758 VSS a_1803_20719# 1e15 m=1
R_D759 VSS a_2021_22325# 1e15 m=1
R_D76 VSS a_2411_26133# 1e15 m=1
R_D760 VSS a_4191_33449# 1e15 m=1
R_D761 VSS a_2959_47113# 1e15 m=1
R_D762 VSS a_4339_64521# 1e15 m=1
R_D763 VSS a_8123_56399# 1e15 m=1
R_D764 VSS a_12357_37999# 1e15 m=1
R_D765 VSS a_7862_34025# 1e15 m=1
R_D766 VSS a_3339_43023# 1e15 m=1
R_D767 VSS a_2411_26133# 1e15 m=1
R_D768 VSS a_6559_59663# 1e15 m=1
R_D769 VSS a_3339_30503# 1e15 m=1
R_D77 VSS a_2419_48783# 1e15 m=1
R_D770 VSS a_7841_12167# 1e15 m=1
R_D771 VSS a_2143_15271# 1e15 m=1
R_D772 VSS a_5682_69367# 1e15 m=1
R_D773 VSS config_2_in[7] 1e15 m=1
R_D774 VSS a_27535_30503# 1e15 m=1
R_D775 VSS a_7862_34025# 1e15 m=1
R_D776 VSS a_4351_67279# 1e15 m=1
R_D777 VSS inn_analog 1e15 m=1
R_D778 VSS a_21371_52263# 1e15 m=1
R_D779 VSS a_2840_66103# 1e15 m=1
R_D78 VSS a_7841_12167# 1e15 m=1
R_D780 VSS a_15607_46805# 1e15 m=1
R_D781 VSS a_11251_59879# 1e15 m=1
R_D782 VSS a_2840_66103# 1e15 m=1
R_D783 VSS a_12355_15055# 1e15 m=1
R_D784 VSS a_43362_28879# 1e15 m=1
R_D785 VSS a_13909_41923# 1e15 m=1
R_D786 VSS a_5363_30503# 1e15 m=1
R_D787 VSS a_2235_30503# 1e15 m=1
R_D788 VSS a_1768_16367# 1e15 m=1
R_D789 VSS a_1586_21959# 1e15 m=1
R_D79 VSS a_12907_27023# 1e15 m=1
R_D790 VSS a_1689_10396# 1e15 m=1
R_D791 VSS a_16955_52047# 1e15 m=1
R_D792 VSS a_2004_42453# 1e15 m=1
R_D793 VSS a_18703_29199# 1e15 m=1
R_D794 VSS a_41261_28335# 1e15 m=1
R_D795 VSS a_4674_40277# 1e15 m=1
R_D796 VSS a_2775_46025# 1e15 m=1
R_D797 VSS a_10055_58791# 1e15 m=1
R_D798 VSS a_5915_30287# 1e15 m=1
R_D799 VSS a_2840_66103# 1e15 m=1
R_D8 VSS a_8531_70543# 1e15 m=1
R_D80 VSS a_18979_30287# 1e15 m=1
R_D800 VSS a_8491_41383# 1e15 m=1
R_D801 VSS a_2143_15271# 1e15 m=1
R_D802 VSS a_3987_19623# 1e15 m=1
R_D803 VSS a_4811_34855# 1e15 m=1
R_D804 VSS a_5915_30287# 1e15 m=1
R_D805 VSS a_11067_63143# 1e15 m=1
R_D806 VSS a_2787_30503# 1e15 m=1
R_D807 VSS a_11067_13095# 1e15 m=1
R_D808 VSS a_25787_28327# 1e15 m=1
R_D809 VSS a_8491_57487# 1e15 m=1
R_D81 VSS config_2_in[10] 1e15 m=1
R_D810 VSS a_20359_29199# 1e15 m=1
R_D811 VSS a_4339_64521# 1e15 m=1
R_D812 VSS a_14831_50095# 1e15 m=1
R_D813 VSS a_2872_44111# 1e15 m=1
R_D814 VSS a_7571_29199# 1e15 m=1
R_D815 VSS a_4215_51157# 1e15 m=1
R_D816 VSS a_12447_29199# 1e15 m=1
R_D817 VSS a_12473_42869# 1e15 m=1
R_D818 VSS a_12381_43957# 1e15 m=1
R_D819 VSS a_2419_48783# 1e15 m=1
R_D82 VSS a_21187_29415# 1e15 m=1
R_D820 VSS a_4119_70741# 1e15 m=1
R_D821 VSS a_1761_52815# 1e15 m=1
R_D822 VSS a_2787_32679# 1e15 m=1
R_D823 VSS a_8295_47388# 1e15 m=1
R_D824 VSS a_13067_38517# 1e15 m=1
R_D825 VSS config_1_in[6] 1e15 m=1
R_D826 VSS a_1586_51335# 1e15 m=1
R_D827 VSS a_1689_10396# 1e15 m=1
R_D828 VSS a_2787_32679# 1e15 m=1
R_D829 VSS a_2411_26133# 1e15 m=1
R_D83 VSS start_conversion_in 1e15 m=1
R_D830 VSS a_18979_30287# 1e15 m=1
R_D831 VSS a_34482_29941# 1e15 m=1
R_D832 VSS a_27535_30503# 1e15 m=1
R_D833 VSS a_5831_39189# 1e15 m=1
R_D834 VSS a_1586_18695# 1e15 m=1
R_D835 VSS a_6467_55527# 1e15 m=1
R_D836 VSS a_27535_30503# 1e15 m=1
R_D837 VSS a_2339_38129# 1e15 m=1
R_D838 VSS a_10055_58791# 1e15 m=1
R_D839 VSS a_12355_15055# 1e15 m=1
R_D84 VSS a_1803_19087# 1e15 m=1
R_D840 VSS a_15607_46805# 1e15 m=1
R_D85 VSS a_4339_64521# 1e15 m=1
R_D86 VSS a_26523_29199# 1e15 m=1
R_D87 VSS a_12725_44527# 1e15 m=1
R_D88 VSS a_15607_46805# 1e15 m=1
R_D89 VSS a_8491_57487# 1e15 m=1
R_D9 VSS a_13123_38231# 1e15 m=1
R_D90 VSS a_3987_19623# 1e15 m=1
R_D91 VSS a_24959_30503# 1e15 m=1
R_D92 VSS a_11067_63143# 1e15 m=1
R_D93 VSS a_10515_63143# 1e15 m=1
R_D94 VSS a_4811_34855# 1e15 m=1
R_D95 VSS a_7571_26151# 1e15 m=1
R_D96 VSS a_1761_44111# 1e15 m=1
R_D97 VSS a_20267_30503# 1e15 m=1
R_D98 VSS a_1586_51335# 1e15 m=1
R_D99 VSS a_11619_56615# 1e15 m=1
R0 VSS dummypin[1] 1e-3 m=1
R1 VSS dummypin[8] 1e-3 m=1
R10 VDD a_82729_53080# 1e-3 m=1
R11 VDD a_82821_19352# 1e-3 m=1
R12 a_17869_27221# VDD 1e-3 m=1
R13 dummypin[7] VSS 1e-3 m=1
R14 VDD a_82821_57432# 1e-3 m=1
R15 VDD a_82821_15000# 1e-3 m=1
R16 a_12809_71285# VSS 1e-3 m=1
R17 a_82729_2197# VDD 1e-3 m=1
R18 a_82729_10901# VDD 1e-3 m=1
R19 a_82729_74005# VDD 1e-3 m=1
R2 VSS a_18007_27441# 1e-3 m=1
R20 a_82729_31573# VDD 1e-3 m=1
R21 VSS dummypin[15] 1e-3 m=1
R22 VSS dummypin[3] 1e-3 m=1
R23 VDD a_12809_23704# 1e-3 m=1
R24 dummypin[9] VSS 1e-3 m=1
R25 VDD a_82821_48728# 1e-3 m=1
R26 VSS a_12809_8945# 1e-3 m=1
R27 VSS dummypin[2] 1e-3 m=1
R28 VSS a_18835_52465# 1e-3 m=1
R29 a_12947_8725# VDD 1e-3 m=1
R3 a_82729_69653# VDD 1e-3 m=1
R30 dummypin[10] VSS 1e-3 m=1
R31 VSS a_12947_56817# 1e-3 m=1
R32 dummypin[0] VSS 1e-3 m=1
R33 dummypin[6] VSS 1e-3 m=1
R34 dummypin[4] VSS 1e-3 m=1
R35 a_18602_55312# VDD 1e-3 m=1
R36 VDD a_82821_28056# 1e-3 m=1
R37 a_82729_6549# VDD 1e-3 m=1
R38 VSS dummypin[14] 1e-3 m=1
R39 VDD a_82821_23704# 1e-3 m=1
R4 dummypin[11] VSS 1e-3 m=1
R40 VDD a_12947_71576# 1e-3 m=1
R41 a_82729_65301# VDD 1e-3 m=1
R42 VDD a_82821_61784# 1e-3 m=1
R43 VSS dummypin[13] 1e-3 m=1
R5 a_12947_23413# VSS 1e-3 m=1
R6 a_12809_56597# VDD 1e-3 m=1
R7 VDD a_82729_78104# 1e-3 m=1
R8 dummypin[5] VSS 1e-3 m=1
R9 dummypin[12] VSS 1e-3 m=1
X0 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=4.54474e+15p pd=2.80061e+10u as=0p ps=0u w=550000u l=2.89e+06u M=254
X1 VDD a_3143_22364# a_4807_27613# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.78423e+15p pd=2.64739e+10u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10 VDD a_7644_46805# a_8126_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X100 VDD a_12877_16911# a_27314_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1000 a_19374_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10000 a_34342_16886# a_16362_16520# a_34434_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10001 a_14859_43447# a_14919_43421# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X10002 a_37846_62516# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10003 VDD a_12981_59343# a_41370_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10004 a_10075_55862# a_7479_54439# a_10003_55862# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X10005 VDD a_35932_41953# a_36520_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10006 vcm_commonmode a_16362_57174# a_18370_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10007 a_38450_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10008 a_24302_72234# VSS a_24394_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10009 VSS a_12727_58255# a_26706_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1001 a_8295_47388# a_10526_22057# a_11390_21807# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X10010 a_22386_55166# VDD a_22294_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10011 VSS a_11067_67279# a_26706_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10012 a_23694_16886# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10013 a_33830_7452# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10014 a_19780_37253# a_18811_36965# a_19743_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10015 a_9983_18870# a_7377_18012# a_9983_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10016 a_21290_10862# a_16362_10496# a_21382_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10017 a_1681_5175# a_1591_7119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10018 VSS a_9215_61127# a_2794_62697# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10019 VDD VDD a_43378_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1002 a_49494_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10020 a_35742_69222# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10021 VDD a_11067_21583# a_27314_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10022 a_26447_42895# a_12549_44212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10023 VDD a_12947_71576# a_31330_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10024 a_7749_20291# a_6816_19355# a_7653_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10025 a_22411_34473# a_21479_34239# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X10026 a_4809_18785# a_4591_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X10027 a_2101_12342# a_1929_12131# a_1887_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X10028 VSS a_24029_39355# a_36579_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X10029 a_31422_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1003 a_21071_37782# a_14293_37455# a_20612_37607# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10030 a_6934_43567# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10031 vcm_commonmode a_16362_23548# a_37446_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10032 a_41462_21540# a_16746_21538# a_41370_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10033 a_36350_58178# a_16362_58178# a_36442_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10034 VDD a_12727_15529# a_17274_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10035 a_20682_9858# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10036 VSS a_7580_61751# a_7837_68591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X10037 a_25702_7850# VDD a_25306_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10038 VDD a_29269_44545# a_30264_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10039 a_18695_47349# a_18539_47617# a_18840_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X1004 a_36842_17492# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10040 VDD a_3339_32463# a_18162_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10041 a_39758_68218# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10042 a_36350_17890# a_12899_10927# a_36842_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10043 a_28410_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10044 VSS a_12546_22351# a_30722_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10045 a_8357_48246# a_6831_63303# a_8143_48246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10046 a_25306_11866# a_16362_11500# a_25398_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10047 a_41783_27247# a_20635_29415# a_9135_27239# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X10048 a_35553_29199# a_15607_46805# a_35263_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10049 a_40858_15484# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1005 a_36746_23914# a_10515_23975# a_36350_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10050 VDD a_12899_10927# a_43378_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10051 a_27183_36965# a_25300_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10052 VSS a_9184_13255# a_7999_13083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10053 a_26413_31055# a_26065_31171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X10054 a_44474_12504# a_16746_12502# a_44382_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10055 a_18770_10464# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10056 VSS a_10515_22671# a_33734_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10057 a_41370_7850# VSS a_41462_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10058 VDD a_10394_19605# a_8933_22583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10059 VDD a_22176_47919# a_22351_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1006 a_34342_18894# a_16362_18528# a_34434_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10060 a_27406_22544# a_16746_22542# a_27314_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10061 vcm_commonmode a_16362_70226# a_36442_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10062 a_44382_69222# a_16362_69222# a_44474_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10063 VSS a_12257_56623# a_46786_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10064 VSS a_5239_45717# a_5173_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10065 VSS a_23540_48981# a_23487_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X10066 VDD a_17488_48731# a_18430_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10067 a_33681_49373# a_33515_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10068 a_17274_7850# VSS a_17366_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10069 VDD a_12970_34191# a_13515_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1007 VDD a_12877_14441# a_40366_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10070 a_41370_11866# a_10055_58791# a_41862_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10071 VSS a_12983_63151# a_29718_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10072 a_26706_64202# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10073 a_6422_11293# a_5345_10927# a_6260_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10074 a_48490_11500# a_16746_11498# a_48398_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10075 a_27406_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10076 VDD a_12727_58255# a_34342_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10077 a_31186_48169# a_27869_50095# a_31114_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10078 VSS a_12447_29199# a_40233_31605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10079 VDD a_12895_13967# a_47394_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1008 VSS a_1586_45431# a_6559_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10080 a_31330_63198# a_16362_63198# a_31422_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10081 VSS a_12901_58799# a_19678_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10082 a_41462_7484# VDD a_41370_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10083 a_23643_41569# a_23789_39100# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10084 VDD a_7050_53333# a_17600_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10085 a_21382_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10086 a_23694_57174# a_10515_22671# a_23298_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10087 VDD a_1591_63151# a_2835_62215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10088 a_17766_16488# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10089 VSS a_2292_43291# a_4761_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1009 a_49798_64202# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10090 vcm_commonmode a_16362_68218# a_30418_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10091 a_10075_55535# a_9821_55862# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10092 a_35463_44031# a_33856_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10093 a_2295_33609# a_1849_33237# a_2199_33609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10094 a_35346_67214# a_12983_63151# a_35838_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10095 vcm_commonmode a_16362_10496# a_18370_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10096 a_20927_35877# a_19780_37253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10097 VDD a_2835_62215# a_2787_62063# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10098 VSS a_1959_26703# a_2099_59861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X10099 VSS a_14289_29687# a_14646_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X101 a_24794_10464# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1010 a_16270_24918# VSS a_16762_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10100 VSS a_6831_63303# a_27388_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X10101 a_48398_66210# a_10975_66407# a_48890_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10102 vcm_commonmode a_16362_9492# a_22386_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10103 a_6913_64239# a_6375_64489# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10104 a_5213_70223# a_4935_70561# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10105 a_2104_52271# a_1987_52484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10106 a_35742_22910# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10107 vcm_commonmode a_16362_59182# a_33430_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10108 a_32426_9492# a_16746_9490# a_32334_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10109 a_42770_23914# a_10515_23975# a_42374_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1011 a_10515_22671# a_15617_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X10110 VSS a_11053_69135# a_11989_68367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X10111 a_7621_18038# a_6816_19355# a_7407_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X10112 VDD a_20881_28111# a_24473_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10113 a_32952_29199# a_12907_27023# a_32649_28853# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10114 VDD a_5671_21495# a_10394_19605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10115 a_33656_43439# a_33479_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10116 a_42866_56492# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10117 a_22294_24918# VSS a_22786_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10118 a_24387_47375# a_23763_47381# a_24279_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10119 a_9503_68841# a_8782_65015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1012 VDD a_7293_49525# a_7183_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X10120 VDD a_12516_7093# a_28318_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10121 a_25798_66532# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10122 a_3392_73853# a_3275_73658# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10123 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10124 a_14097_31375# a_9765_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10125 VDD a_12985_19087# a_47394_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10126 a_32730_15882# a_12877_14441# a_32334_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10127 a_4395_49007# a_3325_49551# a_4032_49159# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X10128 a_28410_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10129 a_25306_56170# a_16362_56170# a_25398_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1013 a_20778_22512# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10130 VSS a_19517_31751# a_18328_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10131 a_39758_21906# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10132 a_7265_56053# a_7803_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X10133 a_22193_49007# a_21003_49007# a_22084_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X10134 VSS VDD a_37750_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10135 a_46882_55488# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10136 a_6637_20407# a_5825_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10137 VSS a_11719_28023# a_11711_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.2575e+11p ps=3.91e+06u w=650000u l=150000u
X10138 VDD a_27155_40871# a_15459_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X10139 a_10053_62581# a_9835_62985# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1014 a_49798_22910# a_11067_21583# a_49402_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10140 a_30326_72234# VDD a_30818_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10141 a_41766_70226# a_12901_66665# a_41370_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10142 a_12165_60975# a_10975_60975# a_12056_60975# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X10143 a_33830_58500# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10144 VSS a_35036_34191# a_35142_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10145 a_29814_65528# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10146 a_26310_62194# a_12355_15055# a_26802_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10147 a_33864_28111# a_15607_46805# a_33761_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10148 a_30818_60508# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10149 VSS a_10055_58791# a_33734_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1015 a_47394_21906# a_11067_21583# a_47886_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10150 a_29322_55166# VSS a_29414_55166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10151 vcm_commonmode a_16362_17524# a_42466_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10152 a_3571_9334# a_1761_8751# a_3112_9527# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X10153 a_2215_12559# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10154 a_7067_30663# a_2787_32679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10155 VSS a_34062_47607# a_33868_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10156 a_28410_71230# a_16746_71232# a_28318_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10157 VSS a_3143_66972# a_7060_61225# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10158 a_24331_34239# a_20715_34717# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10159 VSS a_12985_16367# a_46786_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1016 a_3484_61493# a_3938_61493# a_3876_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X10160 a_19774_57496# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10161 a_6260_74031# a_5179_74031# a_5913_74273# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10162 VDD VSS a_23298_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10163 VSS a_1586_18695# a_7571_16917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10164 a_29322_14878# a_12877_14441# a_29814_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10165 VSS a_12985_7663# a_29718_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10166 a_44778_61190# a_12355_15055# a_44382_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10167 a_45386_9858# a_16362_9492# a_45478_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10168 a_7294_22467# a_5839_22351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10169 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1017 a_47394_17890# a_16362_17524# a_47486_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10170 a_14131_44135# a_3339_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10171 a_27937_27247# a_27659_27275# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X10172 VSS a_12877_16911# a_19678_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10173 a_23694_10862# a_12546_22351# a_23298_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10174 a_6739_59049# a_6880_58773# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10175 VSS a_4032_49159# a_2467_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10176 vcm_commonmode a_16362_21540# a_30418_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10177 VDD a_7925_72399# a_9183_72007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10178 a_46482_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10179 a_48794_60186# a_12981_59343# a_48398_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1018 a_36442_70226# a_16746_70228# a_36350_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10180 VSS a_12899_11471# a_45782_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10181 a_48794_19898# a_12895_13967# a_48398_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10182 a_5924_69135# a_5295_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10183 VDD a_17863_36595# a_17889_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X10184 vcm_commonmode a_16362_18528# a_19374_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10185 a_2250_54813# a_2124_54715# a_1846_54699# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X10186 VDD a_11067_67279# a_33338_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10187 a_6559_59663# a_26218_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10188 a_12983_63151# a_12710_63151# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10189 a_23390_16520# a_16746_16518# a_23298_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1019 a_39758_56170# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10190 vcm_commonmode a_16362_13508# a_20378_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10191 a_32826_18496# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10192 VDD a_1761_37039# a_31131_35281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10193 a_33989_35303# a_34297_35516# a_33963_35507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10194 a_36442_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10195 VDD a_32181_36893# a_31787_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10196 a_27016_29587# a_27169_30083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10197 a_36432_42919# a_35463_42943# a_36395_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10198 a_7255_10357# a_7458_10515# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10199 VDD a_30412_34337# a_30816_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X102 a_28152_40517# a_27183_40229# a_28056_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X1020 a_17763_43413# a_13005_43983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10200 vcm_commonmode a_16362_12504# a_33430_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10201 vcm_commonmode a_16362_63198# a_45478_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10202 a_46390_59182# a_12901_58799# a_46882_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10203 a_6720_15279# a_5639_15279# a_6373_15521# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X10204 a_22690_58178# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10205 a_2776_41167# a_2339_38129# a_2473_40821# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10206 a_34342_24918# VSS a_34434_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10207 a_37846_70548# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10208 VSS a_21387_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10209 a_8297_25071# a_6559_22671# a_8215_25071# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1021 a_31184_40517# a_30311_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10210 a_13669_37429# a_31083_36395# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X10211 VSS a_28524_47919# a_30485_49257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10212 a_34434_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10213 VSS a_34395_31287# a_33798_31145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10214 a_13980_35077# a_13107_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10215 VDD a_1586_9991# a_1591_9839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10216 a_34738_69222# a_12516_7093# a_34342_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10217 a_37354_60186# a_16362_60186# a_37446_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10218 a_16891_36649# a_15959_36415# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10219 a_22386_63198# a_16746_63200# a_22294_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1022 a_5173_45743# a_3983_45743# a_5064_45743# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X10220 a_19127_43439# a_18950_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10221 a_47486_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10222 VSS VDD a_48794_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10223 a_40316_28111# a_13643_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10224 VDD a_10873_27497# a_17691_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10225 VSS a_28599_28023# a_24740_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10226 VSS a_2292_17179# a_3629_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X10227 a_22922_30287# a_5915_35943# a_22836_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10228 a_2647_35951# a_2216_28309# a_2284_36103# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10229 a_12479_8545# a_11067_67279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1023 a_37354_13874# a_12727_15529# a_37846_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10230 vcm_commonmode a_16362_64202# a_49494_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10231 a_30089_41835# a_30023_41959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10232 a_38754_68218# a_12901_66959# a_38358_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10233 a_8061_58575# a_8199_58229# a_8152_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10234 VSS a_12355_65103# a_35742_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10235 a_29718_9858# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10236 vcm_commonmode a_16362_56170# a_39454_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10237 VSS a_3983_68591# a_1923_73087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X10238 VSS a_20881_28111# a_23734_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10239 a_2215_18909# a_1591_18543# a_2107_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X1024 a_8162_53609# a_7749_55535# a_8005_53333# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.65e+11p pd=7.93e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10240 VDD a_26523_28111# a_36448_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10241 a_44778_15882# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10242 a_29391_44031# a_28152_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10243 VDD a_5064_48841# a_5239_48767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10244 a_42985_46831# a_18979_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10245 a_7289_38127# a_4314_40821# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10246 VDD a_4719_51183# a_4215_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10247 a_26402_64202# a_16746_64204# a_26310_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10248 a_6737_60431# a_3143_66972# a_6737_60751# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X10249 a_5800_71855# a_4885_71855# a_5453_72097# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X1025 VSS a_37888_34191# a_37994_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10250 VSS a_2143_15271# a_3983_16617# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10251 VSS a_12947_23413# a_31726_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10252 VSS a_4674_40277# a_19517_31751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10253 a_28410_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10254 a_4676_47607# a_4563_32900# a_4818_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X10255 VDD a_12355_15055# a_35346_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10256 a_31330_56170# a_12947_56817# a_31822_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10257 a_40458_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10258 VDD a_12727_13353# a_39362_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10259 a_31171_27412# a_31263_27221# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1026 a_41862_11468# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10260 a_16362_56170# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X10261 a_17670_17890# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10262 a_37885_43777# a_12357_37999# a_37799_43777# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X10263 a_39396_32143# a_38239_32375# a_39223_32463# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.55e+11p pd=2.51e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X10264 VSS a_12727_13353# a_21686_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10265 a_31873_37253# a_31847_36893# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10266 VSS a_21233_44220# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10267 a_40762_9858# a_12985_19087# a_40366_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10268 a_16832_44007# a_15959_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10269 a_41335_29423# a_39727_27765# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1027 VSS a_11067_13095# a_26706_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10270 VSS clk_vcm a_77972_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10271 a_43774_62194# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10272 a_5730_12265# a_1929_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X10273 a_7039_65469# a_1586_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10274 VDD a_4758_45369# a_4721_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10275 a_26706_72234# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10276 a_8127_39465# a_7948_38377# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10277 VSS a_12516_7093# a_30722_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10278 a_22294_58178# a_10515_22671# a_22786_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10279 VSS a_2319_63388# a_2250_63517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1028 VSS a_12191_37999# a_12357_37999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X10280 a_7850_13967# a_7797_13885# a_7623_13621# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=1.9825e+11p ps=1.91e+06u w=650000u l=150000u
X10281 VDD a_12727_67753# a_34342_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10282 a_22690_11866# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10283 a_23593_41831# a_23901_42044# a_23567_42035# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10284 a_19282_10862# a_16362_10496# a_19374_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10285 a_3705_73461# a_3487_73865# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10286 a_44874_24520# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10287 a_11714_14557# a_10956_14459# a_11151_14428# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10288 VSS a_1586_45431# a_7387_48469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10289 a_34434_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1029 a_7295_25321# a_5211_24759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10290 VSS a_12355_15055# a_20682_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10291 VSS a_1643_59317# a_1591_59343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10292 a_17366_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10293 a_19678_55166# VSS a_19282_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10294 a_34738_64202# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10295 a_47486_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10296 a_6788_30287# a_6752_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X10297 VDD a_2473_34293# a_4053_35523# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X10298 a_34738_22910# a_11067_21583# a_34342_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10299 VDD VSS a_21290_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X103 a_9405_56623# a_5254_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X1030 a_24794_21508# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10300 a_31691_32143# a_31440_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10301 a_4812_13879# a_6435_10901# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X10302 a_48890_23516# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10303 a_1916_33927# a_1915_35015# a_2058_34102# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X10304 a_45386_20902# a_12985_7663# a_45878_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10305 a_45386_16886# a_16362_16520# a_45478_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10306 a_48490_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10307 a_3594_15955# a_3872_15939# a_3828_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10308 a_37465_50095# a_36821_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10309 VDD a_1689_10396# a_2101_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1031 a_24394_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10310 VSS a_24800_41953# a_23901_42044# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X10311 VDD a_2419_55687# a_2419_55535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X10312 a_38850_15484# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10313 a_35346_12870# a_12877_16911# a_35838_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10314 a_38754_21906# a_12985_7663# a_38358_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10315 a_6984_26409# a_5211_24759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10316 VDD a_12877_16911# a_42374_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10317 a_27710_66210# a_12983_63151# a_27314_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10318 VDD a_12947_8725# a_23298_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10319 a_8561_31375# a_2235_30503# a_8215_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X1032 a_21290_14878# a_16362_14512# a_21382_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10320 a_18278_22910# a_10515_23975# a_18770_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10321 a_25447_36919# a_24515_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10322 a_4311_52245# a_4514_52523# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10323 a_26319_41781# a_12641_42036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10324 a_22786_20504# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10325 VDD a_10515_23975# a_25306_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10326 a_22386_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10327 a_5515_32661# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10328 a_49402_15882# a_16362_15516# a_49494_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10329 vcm_commonmode a_16362_8488# a_36442_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1033 a_38867_38591# a_38101_38565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10330 a_25306_64202# a_16362_64202# a_25398_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10331 a_46786_69222# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10332 VSS a_4842_45467# a_4788_45565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10333 a_5755_14709# a_6895_15253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10334 a_16824_28309# a_17278_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X10335 vcm_commonmode VSS a_35438_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10336 a_15290_30761# a_10506_29967# a_15548_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X10337 VDD a_26319_42869# a_19004_40413# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10338 vcm_commonmode a_16362_69222# a_24394_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10339 a_39362_11866# a_10055_58791# a_39854_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1034 a_27314_65206# a_16362_65206# a_27406_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10340 a_8753_19319# a_7377_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10341 a_5449_25071# a_5085_24759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X10342 vcm_commonmode a_16362_23548# a_48490_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10343 a_12549_44212# a_12671_43222# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10344 a_5140_71855# a_5023_72068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10345 VSS a_4771_42167# a_2539_42106# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10346 a_33830_66532# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10347 VDD a_12727_15529# a_28318_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10348 a_26310_70226# a_12516_7093# a_26802_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10349 VSS a_12901_58799# a_40762_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1035 VDD a_12585_39069# a_12191_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X10350 a_26402_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10351 a_23298_12870# a_16362_12504# a_23390_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10352 a_11645_9839# a_11266_10205# a_11573_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10353 a_6519_65301# a_6722_65579# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10354 VSS a_1586_69367# a_7755_74581# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10355 a_29322_63198# a_16362_63198# a_29414_63198# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10356 VSS rst_n a_1591_25615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10357 a_12549_35836# a_13867_35606# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10358 a_2589_55535# a_2419_55535# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10359 vcm_commonmode a_16362_15516# a_38450_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1036 VDD a_19028_35823# a_19134_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10360 a_5094_68086# a_2843_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X10361 VDD a_2744_46983# a_2467_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10362 a_42466_13508# a_16746_13506# a_42374_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10363 a_12954_50639# a_11877_50645# a_12792_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10364 a_21290_8854# a_16362_8488# a_21382_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10365 a_22260_38567# a_21387_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10366 a_5414_39215# a_3949_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10367 VSS a_19807_28111# a_35539_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X10368 a_25398_23548# a_16746_23546# a_25306_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10369 a_10400_62985# a_9485_62613# a_10053_62581# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X1037 a_39454_61190# a_16746_61192# a_39362_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10370 VDD a_5043_19306# a_4379_18756# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X10371 a_6825_29673# a_5441_27791# a_6743_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X10372 a_34342_62194# a_12355_15055# a_34834_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10373 VDD a_9379_15039# a_9366_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10374 a_12631_28585# a_9179_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10375 a_15828_38695# a_16043_38825# a_15970_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X10376 VDD a_2657_60949# a_2605_60975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10377 VDD a_7461_27247# a_8373_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.85e+11p ps=3.57e+06u w=1e+06u l=150000u
X10378 a_9740_62973# a_7676_61493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10379 a_29814_10464# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1038 a_31422_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10380 VSS a_10515_22671# a_44778_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10381 a_18959_50639# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X10382 a_41766_55166# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10383 VSS a_7571_26151# a_12082_25077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10384 VSS a_2292_17179# a_2369_12925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10385 VSS a_12727_67753# a_27710_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10386 a_1761_6031# a_1591_6031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10387 a_47394_61190# a_12981_59343# a_47886_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10388 VDD a_12725_44527# a_30835_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10389 VDD a_7244_39189# a_7847_39872# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1039 vcm_commonmode a_16362_17524# a_36442_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10390 a_32887_42405# a_32121_42369# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10391 a_12631_30511# a_12161_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10392 VSS a_4500_45289# a_4458_45565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10393 VDD a_7377_18012# a_8689_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X10394 a_38358_19898# a_11067_67279# a_38850_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10395 VSS a_1586_40455# a_6559_49557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10396 VSS a_17187_31287# a_16087_31751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10397 a_17191_32117# a_17394_32275# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10398 a_21382_8488# a_16746_8486# a_21290_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10399 a_21686_58178# a_12901_58799# a_21290_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X104 VDD a_7862_34025# a_27139_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1040 a_25605_32259# a_25321_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X10400 a_7159_22583# a_5839_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X10401 a_37926_51727# a_37459_51183# a_6467_55527# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X10402 a_35742_71230# a_12947_71576# a_35346_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10403 VDD a_12355_65103# a_27314_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10404 VSS a_28446_31375# a_29915_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X10405 a_24794_61512# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10406 VSS a_26397_51183# a_32507_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X10407 a_38288_32143# a_32367_28309# a_38115_32463# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X10408 a_5313_43567# a_5269_43809# a_5147_43567# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10409 a_32426_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1041 VSS a_35647_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10410 a_19374_14512# a_16746_14510# a_19282_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10411 a_33363_30305# a_19626_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10412 a_2571_72040# a_2843_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10413 VDD a_3247_20495# a_7621_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10414 VDD a_9123_55223# a_3780_56347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10415 VSS a_1689_10396# a_2108_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10416 a_46390_67214# a_12983_63151# a_46882_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10417 a_6422_74397# a_5345_74031# a_6260_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10418 VDD a_12257_56623# a_17274_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10419 VDD a_35217_44509# a_34823_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1042 a_40458_15516# a_16746_15514# a_40366_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10420 a_19594_35823# a_19417_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10421 VDD a_3949_41935# a_4578_40455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10422 a_11137_9839# a_10659_9813# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10423 a_16035_31375# a_15851_27791# a_15941_31375# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X10424 a_40762_24918# VSS a_40366_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10425 a_28810_60508# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10426 a_34434_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10427 a_77451_38925# a_75794_40594# vcm_commonmode VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X10428 VDD a_4674_40277# a_5831_39189# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10429 a_40858_57496# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1043 VDD a_12727_13353# a_17274_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10430 a_46786_22910# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10431 a_26417_40193# a_25987_41317# a_26860_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10432 a_9740_69501# a_9503_68841# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X10433 vcm_commonmode a_16362_22544# a_24394_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10434 VSS a_8117_12559# a_8056_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10435 a_33338_24918# a_12899_2767# a_33830_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10436 a_23298_57174# a_16362_57174# a_23390_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10437 a_36264_30511# a_26523_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10438 VDD a_23567_43123# a_23593_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10439 VSS a_12899_10927# a_39758_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1044 a_25702_9858# a_12985_19087# a_25306_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10440 a_4497_29673# a_4095_29423# a_4333_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X10441 vcm_commonmode VSS a_49494_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10442 a_43774_15882# a_12877_14441# a_43378_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10443 VSS a_12877_16911# a_40762_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10444 a_30928_52271# a_29361_51727# a_30625_52245# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X10445 a_20713_36929# a_20927_35877# a_21859_35831# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X10446 a_7862_10383# a_7775_10625# a_7458_10515# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X10447 VSS a_35647_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10448 VDD a_12899_11471# a_30326_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10449 a_12749_51183# a_12683_51329# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1045 vcm_commonmode VSS a_49494_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10450 a_2012_45565# a_1867_45743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10451 a_10899_28879# a_10648_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X10452 VDD a_19780_39429# a_19684_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10453 VSS a_15443_29941# a_14354_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10454 VDD a_10391_49855# a_6831_63303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X10455 a_43470_62194# a_16746_62196# a_43378_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10456 a_44874_58500# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10457 vcm_commonmode a_16362_18528# a_40458_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10458 VDD a_12677_40157# a_12283_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10459 VDD a_3325_18543# a_5175_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1046 a_10835_54269# a_10680_52245# a_10472_54135# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X10460 a_26402_72234# VDD a_26310_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10461 VSS a_20535_51727# a_21267_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10462 a_47790_14878# a_12727_15529# a_47394_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10463 VSS a_10055_58791# a_44778_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10464 a_10659_9813# a_10862_10091# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10465 a_28426_29941# a_28680_30057# a_28638_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10466 VSS a_35033_42044# a_34725_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10467 a_8950_13763# a_1929_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10468 VSS a_3112_9527# a_3063_9295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10469 a_27314_15882# a_12727_13353# a_27806_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1047 a_6372_38279# a_7061_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X10470 VSS a_11067_21583# a_27710_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10471 a_20514_28111# a_15661_29199# a_20442_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X10472 a_13445_51335# a_13445_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10473 VDD a_2686_70223# a_7063_70313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10474 VSS a_5239_65301# a_5682_69367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X10475 a_31822_13476# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10476 VSS a_35969_28111# a_36459_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10477 a_21675_43447# a_20743_43493# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10478 a_20286_9858# a_12546_22351# a_20778_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10479 a_6985_25615# a_4571_26677# a_7343_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X1048 VDD a_6611_14967# a_5465_14967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10480 a_4065_13103# a_2873_13879# a_3843_13880# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10481 a_10197_18870# a_7377_18012# a_9983_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X10482 a_4581_60797# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10483 a_8491_57487# a_10680_52245# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X10484 VDD a_12901_58799# a_21290_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10485 VDD a_3339_30503# a_26350_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10486 VSS a_12727_15529# a_17670_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10487 a_21686_11866# a_12985_16367# a_21290_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10488 a_30818_9460# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10489 a_30418_17524# a_16746_17522# a_30326_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1049 VSS a_9751_25071# a_11163_25321# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X10490 VDD a_36392_43677# a_35493_43421# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X10491 a_26523_28111# a_35907_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10492 a_75199_40594# a_75111_40050# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10493 a_41370_70226# a_16362_70226# a_41462_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10494 VDD a_10575_69439# a_10562_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10495 a_22294_66210# a_10975_66407# a_22786_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10496 a_33734_64202# a_12355_65103# a_33338_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10497 vcm_commonmode a_16362_60186# a_17366_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10498 vcm_commonmode a_16362_19532# a_17366_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10499 a_1757_29973# a_1591_29973# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X105 a_39799_38825# a_38867_38591# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X1050 a_18370_10496# a_16746_10494# a_18278_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10500 VDD a_4220_57685# a_2944_57960# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10501 a_34434_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10502 VSS a_32371_32117# a_23395_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10503 a_4499_48841# a_3983_48469# a_4404_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X10504 vcm_commonmode a_16362_13508# a_31422_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10505 VDD a_11067_67279# a_44382_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10506 a_19678_63198# a_15439_49525# a_19282_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10507 a_26523_29199# a_26350_28585# a_27214_28335# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X10508 a_34738_72234# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10509 a_21095_51727# a_19478_51959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X1051 a_27806_12472# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10510 a_47486_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10511 a_10473_11809# a_10317_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10512 a_46882_8456# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10513 a_42770_8854# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10514 a_8197_15279# a_7841_12167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10515 VSS a_2787_30503# a_24223_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10516 a_33734_58178# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10517 a_33603_47081# a_22291_29415# a_33385_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10518 a_47790_71230# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10519 a_46482_69222# a_16746_69224# a_46390_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1052 a_25306_13874# a_16362_13508# a_25398_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10520 vcm_commonmode a_16362_66210# a_43470_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10521 VDD a_10055_58791# a_34342_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10522 a_37287_51433# a_37307_51339# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X10523 a_41872_29423# a_41335_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X10524 a_45386_24918# VSS a_45478_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10525 a_4157_32259# a_1915_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10526 a_8143_44982# a_7295_44647# a_8071_44982# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X10527 a_45478_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10528 a_48398_60186# a_16362_60186# a_48490_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10529 VSS a_12985_19087# a_28714_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1053 a_1895_14906# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10530 VSS a_12981_59343# a_41766_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10531 a_3877_57167# a_3521_57283# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10532 a_19559_43177# a_18627_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10533 a_1761_44111# a_1591_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10534 a_29322_56170# a_12947_56817# a_29814_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10535 VSS a_4219_34551# a_3187_34293# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10536 a_38450_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10537 a_75162_40202# a_75258_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10538 a_10103_11079# a_9484_11989# a_10337_10927# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10539 a_23849_30511# a_22151_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1054 VDD a_12546_22351# a_31330_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10540 VSS a_12901_66665# a_24698_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10541 a_11617_66415# a_11521_66567# a_9513_65301# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X10542 a_4404_65327# a_4287_65540# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10543 a_20378_66210# a_16746_66212# a_20286_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10544 vcm_commonmode a_16362_65206# a_47486_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10545 VDD a_12985_16367# a_38358_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10546 a_6451_22895# a_6007_23145# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10547 a_22386_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10548 VDD a_32970_31145# a_40323_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10549 a_49402_23914# a_16362_23548# a_49494_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1055 a_48890_66532# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10550 a_38704_52047# a_35568_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X10551 a_22531_51017# a_22181_50645# a_22436_51005# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X10552 a_25398_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10553 vcm_commonmode a_16362_57174# a_37446_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10554 a_13097_35279# a_12831_35645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10555 a_41167_42943# a_37551_42333# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10556 a_49798_68218# a_12901_66959# a_49402_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10557 VSS a_5963_20149# a_8583_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.565e+11p ps=5.92e+06u w=650000u l=150000u
X10558 a_41462_55166# VDD a_41370_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10559 a_42770_16886# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1056 a_45386_63198# a_12981_62313# a_45878_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10560 VDD a_10825_29688# a_10761_29745# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.344e+11p ps=1.48e+06u w=420000u l=150000u
X10561 a_10614_52598# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X10562 VSS a_12516_7093# a_28714_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10563 a_40366_10862# a_16362_10496# a_40458_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10564 a_33049_28585# a_24959_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10565 a_24394_65206# a_16746_65208# a_24302_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10566 ctopn a_8583_33551# ctopn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u M=2
X10567 VDD a_2235_30503# a_25462_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X10568 a_23298_20902# a_16362_20536# a_23390_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10569 a_26402_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1057 VDD a_4717_65569# a_4607_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X10570 VDD a_12981_62313# a_33338_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10571 VSS a_6224_73095# a_7289_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X10572 VDD a_2122_19087# a_2228_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10573 VSS a_12355_15055# a_18674_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10574 VSS a_23789_39100# a_24208_39453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10575 a_25306_7850# VDD a_25798_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10576 VDD a_12355_15055# a_46390_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10577 a_22690_60186# a_12981_59343# a_22294_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10578 a_22690_19898# a_12895_13967# a_22294_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10579 a_2216_42997# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1058 a_36442_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10580 VSS a_28152_40517# a_28115_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X10581 a_2467_29397# a_2347_28918# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10582 vcm_commonmode a_16362_8488# a_44474_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10583 a_27406_56170# a_16746_56172# a_27314_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10584 a_7953_13967# a_7917_13885# a_7850_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10585 a_16891_35561# a_15959_35327# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10586 a_28714_17890# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10587 a_19678_7850# VDD a_19282_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10588 a_34342_70226# a_12516_7093# a_34834_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10589 a_6106_34863# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1059 a_12725_44527# a_12559_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X10590 a_3670_42301# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10591 VSS a_12727_13353# a_32730_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10592 a_31726_7850# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10593 a_41766_63198# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10594 a_38358_68218# a_16362_68218# a_38450_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10595 VSS a_10382_58487# a_10331_58255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10596 VDD a_15439_49525# a_19282_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10597 a_21490_28585# a_20747_27765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X10598 a_44382_11866# a_16362_11500# a_44474_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10599 a_20286_59182# a_12901_58799# a_20778_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X106 a_6094_67825# a_6156_67477# a_6093_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.323e+11p ps=1.47e+06u w=420000u l=150000u
X1060 a_2012_23805# a_1867_23983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X10600 VDD a_4811_34855# a_23498_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10601 vcm_commonmode a_16362_62194# a_32426_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10602 a_33430_23548# a_16746_23546# a_33338_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10603 a_33338_58178# a_10515_22671# a_33830_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10604 VDD a_6224_73095# a_7761_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10605 VDD a_24800_35425# a_25204_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10606 a_12135_69109# a_11955_69653# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10607 a_17103_49007# a_16753_49007# a_17008_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X10608 a_33734_11866# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10609 a_46482_22544# a_16746_22542# a_46390_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1061 a_44474_14512# a_16746_14510# a_44382_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10610 VSS a_13837_38772# a_15129_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X10611 VSS a_2952_66139# a_7479_67075# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10612 a_24773_48463# a_24209_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u
X10613 a_7251_43894# a_7000_43541# a_6792_43719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10614 VDD VDD a_27314_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10615 a_45478_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10616 VSS config_2_in[8] a_1591_41935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10617 a_7708_46287# a_7494_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10618 a_21382_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10619 a_8143_44655# a_7889_44982# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1062 a_25764_51183# a_24683_51183# a_25417_51425# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X10620 VDD config_2_in[6] a_1591_39215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X10621 a_4702_32143# a_4263_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X10622 VSS a_12983_63151# a_48794_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10623 a_45782_64202# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10624 VDD a_1586_40455# a_1591_43029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10625 a_43378_21906# a_11067_21583# a_43870_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10626 VSS a_1923_59583# a_11753_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10627 a_14049_42869# a_13716_43047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10628 a_43378_17890# a_16362_17524# a_43470_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10629 a_5113_64061# a_4734_63695# a_5041_64061# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1063 vcm_commonmode a_16362_11500# a_41462_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10630 a_35438_7484# VDD a_35346_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10631 a_35932_38689# a_35647_39141# a_36520_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10632 VSS a_12901_58799# a_38754_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10633 a_35742_56170# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10634 VDD a_3949_41935# a_4706_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X10635 a_42770_57174# a_10515_22671# a_42374_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10636 a_36842_16488# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10637 a_7578_46831# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10638 VDD a_7050_53333# a_17210_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X10639 a_4446_40553# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X1064 a_24515_43493# a_20899_44211# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10640 a_18674_66210# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10641 a_25702_67214# a_12727_67753# a_25306_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10642 VSS a_11067_13095# a_22690_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10643 a_14258_44527# a_14081_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10644 a_8031_24527# a_4351_26703# a_8113_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10645 VSS a_31741_30485# a_30891_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X10646 VDD a_22151_29941# a_22243_30491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10647 a_49894_15484# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10648 vcm_commonmode a_16362_10496# a_37446_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10649 a_49798_21906# a_12985_7663# a_49402_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1065 a_8176_74941# a_8059_74746# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10650 a_46390_12870# a_12877_16911# a_46882_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10651 a_20778_21508# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10652 a_20378_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10653 VSS a_11067_23759# a_16362_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X10654 a_23298_65206# a_16362_65206# a_23390_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10655 a_2834_66781# a_1757_66415# a_2672_66415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10656 a_35438_61190# a_16746_61192# a_35346_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10657 a_2325_14709# a_2107_15113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10658 a_17799_38591# a_17033_38565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X10659 vcm_commonmode VSS a_33430_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1066 a_3118_33597# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X10660 a_39758_55166# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10661 a_39758_13874# a_12877_16911# a_39362_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10662 a_23481_31171# a_14646_29423# a_23385_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X10663 a_5411_12791# a_1929_12131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10664 a_4952_68279# a_5167_68060# a_5094_68086# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X10665 vcm_commonmode VSS a_46482_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10666 a_24515_34789# a_20623_36595# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10667 a_20378_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10668 VDD a_12877_14441# a_26310_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10669 VSS a_32029_38565# a_33543_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X1067 vcm_commonmode a_16362_56170# a_30418_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10670 a_21290_13874# a_16362_13508# a_21382_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10671 VDD a_12516_7093# a_47394_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10672 a_44874_66532# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10673 VSS a_2317_28892# a_5087_23145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10674 a_41370_63198# a_12981_62313# a_41862_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10675 a_39454_60186# a_16746_60188# a_39362_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10676 vcm_commonmode a_16362_16520# a_36442_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10677 a_39454_19532# a_16746_19530# a_39362_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10678 VSS VSS a_16666_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10679 a_8916_19203# a_7377_18012# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1068 a_12605_55311# a_12371_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X10680 a_40458_14512# a_16746_14510# a_40366_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10681 a_44382_56170# a_16362_56170# a_44474_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10682 VDD a_6373_15521# a_6263_15645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10683 VSS a_2411_19605# a_2369_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10684 VDD a_22632_42919# a_22536_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X10685 a_30722_61190# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10686 a_29322_9858# a_12546_22351# a_29814_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10687 VSS a_30035_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10688 a_27314_66210# a_16362_66210# a_27406_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10689 a_27806_11468# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1069 a_40858_19500# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10690 a_7910_38671# a_5631_38127# a_8177_38991# VSS sky130_fd_pr__nfet_01v8 ad=1.9825e+11p pd=1.91e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X10691 a_4883_33053# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X10692 a_17766_68540# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10693 VDD a_12983_63151# a_21290_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10694 a_48890_65528# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10695 a_45386_62194# a_12355_15055# a_45878_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10696 a_2375_48084# a_2467_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X10697 a_6926_70339# a_2952_66139# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X10698 a_3357_67257# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10699 a_21382_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X107 a_48794_59182# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1070 a_27406_24552# VDD a_27314_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10700 VSS a_7221_43541# a_7155_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10701 vcm_commonmode VSS a_30418_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10702 VSS a_42941_32143# a_41842_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X10703 a_38850_57496# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10704 VSS a_4584_20407# a_3799_20407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10705 VDD VSS a_42374_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10706 a_33734_72234# VDD a_33338_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10707 VDD a_7039_65469# a_7000_65595# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10708 VSS a_12985_7663# a_48794_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10709 VDD a_12985_19087# a_40366_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1071 a_24473_31171# a_15548_30761# a_24401_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10710 a_18278_64202# a_11067_13095# a_18770_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10711 VDD a_10975_66407# a_25306_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10712 a_22786_62516# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10713 VSS a_6327_14343# a_6277_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10714 a_12723_13647# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X10715 a_46786_71230# a_12947_71576# a_46390_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10716 VSS a_12877_16911# a_38754_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10717 a_42770_10862# a_12546_22351# a_42374_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10718 VDD a_19807_28111# a_31522_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10719 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1072 a_10055_58791# a_7000_43541# a_12263_48783# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X10720 a_25702_20902# a_11067_67279# a_25306_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10721 VDD a_12889_39889# a_12831_39997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X10722 a_16928_44007# a_15959_44031# a_16832_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10723 VDD a_12257_56623# a_28318_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10724 VDD a_9135_29423# a_9135_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10725 a_20682_69222# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10726 a_16746_15514# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X10727 a_8583_22671# a_8933_22583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10728 VSS a_4811_34855# a_34016_31849# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10729 a_45478_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1073 VDD a_12257_56623# a_42374_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10730 VSS a_41636_37601# a_42283_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X10731 VSS a_11495_16341# a_11429_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10732 a_35598_49551# a_35568_49525# a_35224_49871# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X10733 vcm_commonmode a_16362_23548# a_22386_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10734 a_36711_29199# a_32823_29397# a_36615_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10735 a_38213_47081# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X10736 a_30679_43493# a_29913_43457# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10737 a_25759_32259# a_25321_29673# a_25687_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10738 a_21290_58178# a_16362_58178# a_21382_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10739 a_35346_71230# a_16362_71230# a_35438_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1074 VSS a_10409_18543# a_10791_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X10740 VSS a_12895_13967# a_37750_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10741 a_32795_36415# a_31280_36165# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10742 a_41766_16886# a_12727_13353# a_41370_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10743 VSS a_35647_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10744 a_24698_68218# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10745 a_5132_58255# a_4918_58255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X10746 a_1925_18231# a_2021_17973# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10747 VSS a_8275_43255# a_8171_43541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10748 a_21290_17890# a_12899_10927# a_21782_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10749 a_2163_64381# a_1586_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1075 VDD a_5535_18012# a_10786_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X10750 VDD a_4308_45431# a_4259_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10751 a_28410_17524# a_16746_17522# a_28318_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10752 a_7571_22057# a_5085_23047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X10753 a_24394_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10754 a_7365_46653# a_6655_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X10755 a_41462_63198# a_16746_63200# a_41370_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10756 a_39362_70226# a_16362_70226# a_39454_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10757 a_42866_59504# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10758 a_38754_14878# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10759 vcm_commonmode a_16362_70226# a_21382_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1076 VSS a_41820_41501# a_40921_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X10760 a_27710_59182# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10761 VSS a_12257_56623# a_31726_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10762 a_8461_32937# a_2787_32679# a_8307_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10763 a_15129_38543# a_14859_38909# a_15039_38909# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10764 VDD a_12901_66665# a_33338_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10765 a_25306_16886# a_12899_11471# a_25798_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10766 a_35550_27791# a_35616_27765# a_35383_28111# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10767 VSS a_1586_45431# a_9779_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10768 a_4406_37949# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10769 a_5905_57711# a_1823_65853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1077 VDD a_12983_63151# a_25306_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10770 a_5173_44655# a_4842_45467# a_5185_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10771 a_52778_39936# a_52590_39936# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10772 a_33430_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10773 vcm_commonmode a_16362_13508# a_29414_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10774 a_10151_21379# a_7377_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10775 a_5594_36727# a_5691_36727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10776 VDD a_11067_13095# a_12877_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X10777 a_16362_70226# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X10778 a_30665_30511# a_30790_30663# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X10779 a_43680_29941# a_26523_29199# a_44273_30287# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1078 a_22786_63520# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10780 a_14625_30761# a_10506_29967# a_14553_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X10781 a_8636_63669# a_4339_64521# a_8856_64015# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X10782 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10783 a_1586_21959# a_1643_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10784 VSS a_35815_31751# a_16863_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X10785 VDD a_2939_52245# a_2926_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10786 VDD a_23567_42035# a_23593_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10787 VDD a_12947_71576# a_19282_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10788 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X10789 a_9253_24011# a_6559_22671# a_9167_24011# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1079 a_49402_62194# a_12355_15055# a_49894_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10790 a_20286_67214# a_12983_63151# a_20778_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10791 a_12203_54475# a_12202_54599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10792 VDD VDD a_45386_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10793 VSS a_23271_50943# a_23205_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X10794 VSS VDD a_41766_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X10795 a_5013_20473# a_3247_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10796 a_6260_74031# a_5345_74031# a_5913_74273# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X10797 a_19374_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10798 a_8494_10383# a_7736_10499# a_7931_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10799 VSS a_26319_35253# a_15968_36061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X108 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u M=564
X1080 a_17366_16520# a_16746_16518# a_17274_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10800 a_33338_66210# a_10975_66407# a_33830_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10801 a_34738_9858# a_12985_19087# a_34342_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10802 a_44778_64202# a_12355_65103# a_44382_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10803 vcm_commonmode a_16362_60186# a_28410_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10804 vcm_commonmode a_16362_19532# a_28410_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10805 a_18370_66210# a_16746_66212# a_18278_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10806 a_6661_42255# a_6607_42167# a_6579_42255# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10807 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=5.1e+06u w=1.89e+07u
X10808 VDD a_19780_38341# a_19684_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10809 a_20682_22910# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1081 a_16746_67216# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X10810 a_45478_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10811 a_17274_21906# a_16362_21540# a_17366_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10812 a_22690_9858# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10813 a_34738_56170# a_12257_56623# a_34342_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10814 a_27710_7850# VDD a_27314_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10815 a_45782_72234# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10816 vcm_commonmode a_16362_67214# a_41462_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10817 a_3789_28995# a_1915_35015# a_3707_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10818 VSS a_7000_43541# a_13461_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X10819 VSS a_11855_51959# a_11801_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1082 VSS a_17682_50095# a_32580_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X10820 a_12227_51017# a_11711_50645# a_12132_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X10821 VSS a_12546_22351# a_32730_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10822 VSS a_7244_39189# a_7188_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10823 VDD a_28295_31287# a_28089_31157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5795e+11p ps=2.99e+06u w=420000u l=150000u
X10824 a_24937_39306# a_1761_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X10825 VSS a_6831_63303# a_30125_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10826 VSS a_7939_30503# a_27169_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10827 a_24698_21906# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10828 VDD a_32367_28309# a_38288_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10829 a_5357_62313# a_3016_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X1083 a_8203_23145# a_8105_21263# a_7841_22895# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X10830 a_27314_57174# a_12257_56623# a_27806_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10831 a_43378_7850# VSS a_43470_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10832 a_36442_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10833 a_38754_55166# VSS a_38358_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10834 a_2399_47375# a_1775_47381# a_2291_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X10835 a_31822_55488# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10836 VSS VDD a_22690_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10837 a_11599_55901# a_10975_55535# a_11491_55535# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X10838 a_5483_11140# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10839 a_49494_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1084 a_22786_8456# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10840 VSS a_34759_31029# a_41397_30333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10841 a_10472_52423# a_10687_52553# a_10614_52598# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X10842 a_19282_7850# VSS a_19374_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10843 VSS a_28881_52271# a_34895_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10844 VDD a_12985_16367# a_49402_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10845 VDD VSS a_40366_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10846 VDD a_12901_66959# a_39362_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10847 a_27710_12870# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10848 a_39758_63198# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10849 vcm_commonmode a_16362_58178# a_35438_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1085 a_25015_48437# a_25019_47679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10850 VSS a_12985_16367# a_31726_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10851 VDD a_33486_34191# a_34859_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10852 a_29414_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10853 VDD a_5839_22351# a_6257_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10854 VDD a_37076_37253# a_36980_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10855 VDD a_3173_46805# a_3203_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10856 vcm_commonmode a_16362_68218# a_18370_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10857 vcm_commonmode a_16362_57174# a_48490_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10858 a_19113_51005# a_19069_50613# a_18947_51017# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X10859 a_43470_7484# VDD a_43378_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1086 VSS a_21041_37429# a_20975_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10860 a_32769_29423# a_4811_34855# a_30790_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10861 VDD a_4811_34855# a_32319_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10862 a_37354_22910# a_10515_23975# a_37846_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X10863 a_41370_71230# a_12901_66665# a_41862_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10864 a_14258_34191# a_14081_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10865 a_41862_20504# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10866 a_41462_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10867 a_2834_38671# a_1757_38677# a_2672_39049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10868 VDD a_12981_62313# a_44382_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10869 a_44382_64202# a_16362_64202# a_44474_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1087 VDD a_14919_43421# a_14945_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10870 a_18829_29423# a_18551_29451# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X10871 vcm_commonmode a_16362_9492# a_24394_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10872 VSS a_12355_15055# a_29718_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10873 a_25398_57174# a_16746_57176# a_25306_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10874 a_26706_18894# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10875 a_31422_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10876 VSS a_12899_11471# a_30722_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10877 a_45386_70226# a_12516_7093# a_45878_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10878 VDD a_12727_15529# a_47394_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10879 VSS a_22351_47893# a_7571_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X1088 a_12407_54965# a_12481_54447# a_12605_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X10880 VDD a_2419_48783# a_2971_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10881 a_2169_74913# a_1586_69367# a_2083_74913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X10882 a_42374_12870# a_16362_12504# a_42466_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10883 a_9513_65301# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10884 a_8638_65103# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.7125e+11p pd=4.05e+06u as=0p ps=0u w=650000u l=150000u
X10885 a_21382_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10886 a_31127_29423# a_30790_30663# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10887 VSS a_12901_66959# a_42770_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10888 a_7583_12265# a_1929_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X10889 vcm_commonmode a_16362_63198# a_30418_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1089 VDD a_7467_61751# a_3938_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X10890 a_31330_59182# a_12901_58799# a_31822_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10891 a_28671_30539# a_28670_30663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10892 a_23096_51017# a_22015_50645# a_22749_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10893 a_31223_36369# a_1761_39215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10894 VSS a_19576_51701# a_22169_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10895 a_44474_23548# a_16746_23546# a_44382_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10896 a_22291_29415# a_36401_46859# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u M=2
X10897 a_18278_72234# VDD a_18770_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10898 vcm_commonmode a_16362_20536# a_41462_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10899 a_18770_21508# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X109 VSS a_12727_67753# a_22690_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1090 a_10678_14443# a_10956_14459# a_10912_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X10900 a_3487_37961# a_3137_37589# a_3392_37949# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X10901 a_18370_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10902 a_22786_70548# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10903 a_48890_10464# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10904 a_2012_21807# a_1867_21263# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10905 VDD a_7213_62215# a_7171_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10906 a_4968_60405# a_5421_60137# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X10907 a_22294_60186# a_16362_60186# a_22386_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10908 VSS a_12727_67753# a_46786_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10909 a_43774_65206# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1091 a_41462_9492# a_16746_9490# a_41370_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10910 a_34434_15516# a_16746_15514# a_34342_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10911 VSS a_5039_42167# a_11067_66191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X10912 a_32426_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10913 VSS a_2805_22869# a_2739_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10914 VDD a_2451_72373# a_2409_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X10915 a_41370_18894# a_16362_18528# a_41462_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10916 a_28884_41831# a_28011_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10917 a_5295_69135# a_5213_70223# a_5489_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X10918 a_16832_36391# a_15959_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10919 a_10296_55535# a_7479_54439# a_10075_55862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1092 a_6735_36611# a_4314_40821# a_6653_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10920 a_15697_28335# a_14273_27791# a_15788_28335# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=0p ps=0u w=650000u l=150000u
X10921 a_15851_27791# a_14273_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10922 a_2847_71615# a_2672_71689# a_3026_71677# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X10923 a_19282_13874# a_16362_13508# a_19374_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10924 VDD a_12546_22351# a_25306_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10925 VDD a_24893_37429# a_24837_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X10926 a_40762_58178# a_12901_58799# a_40366_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10927 a_16746_23546# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X10928 a_39362_63198# a_12981_62313# a_39854_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10929 VSS a_12901_58799# a_49798_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1093 a_37750_72234# VDD a_37354_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10930 a_23694_68218# a_12901_66959# a_23298_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10931 VSS a_12355_65103# a_20682_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10932 a_12712_62313# a_11067_63143# a_12621_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X10933 a_43870_61512# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10934 a_46786_56170# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10935 a_47394_9858# a_16362_9492# a_47486_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10936 a_42224_39429# a_41351_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X10937 a_38450_14512# a_16746_14510# a_38358_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10938 vcm_commonmode a_16362_11500# a_35438_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10939 a_5671_21495# a_11495_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X1094 a_7097_40303# a_6671_40630# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10940 a_47886_16488# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10941 VSS a_4227_37887# a_4161_37961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X10942 a_13335_27497# a_11866_27791# a_13241_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X10943 a_10301_66237# a_9513_65301# a_10229_66237# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X10944 vcm_commonmode a_16362_56170# a_24394_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10945 a_34834_19500# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10946 vcm_commonmode a_16362_21540# a_18370_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10947 vcm_commonmode a_16362_10496# a_48490_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10948 a_4496_18543# a_4379_18756# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10949 a_2405_19087# a_2228_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1095 a_18456_47375# a_17787_47349# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X10950 VDD a_19492_52245# a_12659_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X10951 a_26514_47375# a_26259_47491# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X10952 a_4503_21523# a_4839_21495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X10953 a_2325_23413# a_2107_23817# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X10954 VDD a_18045_38017# a_19224_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X10955 a_26706_59182# a_12727_58255# a_26310_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10956 a_1761_6031# a_1591_6031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X10957 a_9215_61127# a_8500_58799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10958 VDD a_12355_15055# a_20286_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10959 a_21516_47919# a_19788_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1096 a_26802_62516# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10960 a_7457_56053# a_6927_56873# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10961 a_7758_65693# a_7000_65595# a_7195_65564# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X10962 a_2520_16911# a_2040_17289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10963 a_6725_45205# a_6559_45205# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10964 VDD a_12727_13353# a_24302_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10965 a_38358_69222# a_12901_66959# a_38850_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10966 a_42866_67536# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10967 a_25398_10496# a_16746_10494# a_25306_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10968 VSS a_20927_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X10969 a_1823_53885# a_2939_52245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1097 VDD a_4035_54965# a_1823_58773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10970 a_11173_12015# a_11138_12267# a_10935_11989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X10971 a_42374_57174# a_16362_57174# a_42466_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10972 a_25306_67214# a_16362_67214# a_25398_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X10973 VSS VSS a_27710_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10974 a_10984_58487# a_11080_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10975 a_13047_29575# a_6459_30511# a_13516_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X10976 a_35932_37601# a_35647_38053# a_36520_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X10977 a_2737_68413# a_2693_68021# a_2571_68425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X10978 VSS a_10515_23975# a_42770_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10979 a_39454_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1098 a_31330_67214# a_16362_67214# a_31422_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X10980 a_2289_35113# a_1915_35015# a_2217_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X10981 VSS a_25015_48437# a_26273_48801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10982 a_2203_45577# a_1757_45205# a_2107_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10983 VSS a_12755_51562# a_13735_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X10984 VDD a_3016_60949# a_5905_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10985 a_11307_57711# a_10791_57711# a_11212_57711# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X10986 a_35742_17890# a_12899_11471# a_35346_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X10987 a_13239_29575# a_12965_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X10988 a_32426_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10989 a_4500_45289# a_4443_46607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 VDD a_12981_59343# a_30326_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X10990 a_16191_38543# a_16043_38825# a_15828_38695# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X10991 VDD a_3305_38671# a_6607_39991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10992 VDD a_7815_45503# a_7802_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10993 VSS a_11067_21583# a_46786_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10994 VSS a_20592_46983# a_20543_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10995 a_26985_31605# a_25321_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X10996 a_4037_58773# a_3141_59887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10997 a_2856_47753# a_1775_47381# a_2509_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10998 a_49894_57496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X10999 a_44778_72234# VDD a_44382_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u M=777
X110 a_42374_61190# a_12981_59343# a_42866_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1100 a_18162_31055# a_13353_30511# a_18162_31375# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X11000 a_19282_58178# a_16362_58178# a_19374_58178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11001 a_30326_20902# a_12985_7663# a_30818_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11002 a_30326_16886# a_16362_16520# a_30418_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11003 VDD a_12901_58799# a_40366_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11004 VDD a_77972_39480# a_77664_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11005 VSS a_12727_15529# a_36746_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11006 VSS a_24893_37429# a_24837_37782# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11007 a_40762_11866# a_12985_16367# a_40366_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11008 a_22084_49007# a_21169_49007# a_21737_49249# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11009 a_19282_17890# a_12899_10927# a_19774_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1101 a_9465_53903# a_7155_55509# a_9031_54135# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X11010 VSS a_12947_23413# a_19678_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11011 a_7725_72765# a_6453_71855# a_7653_72765# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11012 a_14088_37455# a_13097_37455# a_13867_37782# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11013 a_23790_15484# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11014 a_4866_13967# a_4812_13879# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.7125e+11p pd=4.05e+06u as=0p ps=0u w=650000u l=150000u
X11015 VSS a_12877_16911# a_49798_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11016 a_23694_21906# a_12985_7663# a_23298_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11017 VSS a_21049_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X11018 a_12056_60975# a_11141_60975# a_11709_61217# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11019 VDD a_12407_54965# a_11710_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1102 a_43680_29941# a_41597_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X11020 a_20286_12870# a_12877_16911# a_20778_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11021 a_12805_68367# a_11710_58487# a_11947_68279# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11022 VDD a_10515_22671# a_26310_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11023 VDD a_22632_41831# a_22536_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X11024 a_7999_40553# a_5363_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11025 a_4425_32687# a_4259_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11026 a_6010_56989# a_5252_56891# a_5447_56860# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11027 vcm_commonmode a_16362_70226# a_19374_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11028 a_31726_69222# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11029 vcm_commonmode a_16362_18528# a_49494_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1103 a_45478_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11030 vcm_commonmode VSS a_20378_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11031 a_26706_12870# a_10055_58791# a_26310_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11032 a_38754_63198# a_15439_49525# a_38358_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11033 VSS a_12727_58255# a_35742_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11034 a_42770_9858# a_12985_19087# a_42374_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11035 a_24302_11866# a_10055_58791# a_24794_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11036 a_36746_8854# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11037 VSS a_11067_67279# a_35742_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11038 VSS a_51330_39932# a_52590_39198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.55e+11p ps=1.62e+06u w=500000u l=150000u
X11039 VSS a_40383_29575# a_28841_29575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1104 a_2805_22869# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11040 a_4273_55357# a_4238_55123# a_4035_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11041 vcm_commonmode a_16362_23548# a_33430_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11042 a_28423_52245# a_28248_52271# a_28602_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11043 a_46390_71230# a_16362_71230# a_46482_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11044 VDD a_12727_58255# a_17274_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11045 a_21041_37429# a_18127_35797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11046 a_7295_44647# a_17651_30485# a_17589_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11047 a_2369_21807# a_2325_22049# a_2203_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11048 VDD a_9828_56311# a_9599_57141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11049 a_26402_18528# a_16746_18526# a_26310_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1105 VSS a_12587_51335# a_11855_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11050 VDD a_11067_21583# a_36350_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11051 a_4988_67753# a_3325_69135# a_4906_67509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11052 vcm_commonmode a_16362_15516# a_23390_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11053 a_17939_43745# a_13716_43047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11054 VSS a_21233_44220# a_20925_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11055 a_11898_10205# a_11140_10107# a_11335_10076# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11056 a_4811_34855# a_23195_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X11057 a_7841_29673# a_5087_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11058 a_40458_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11059 a_7002_21263# a_2339_38129# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1106 a_7933_51433# a_2840_66103# a_7933_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X11060 VSS a_4311_52245# a_1823_63677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11061 a_1846_54699# a_2163_54589# a_2121_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11062 VDD a_18979_30287# a_30190_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X11063 a_4711_54965# a_4516_55107# a_5021_55357# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X11064 VSS a_12901_66665# a_43774_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11065 a_7494_46287# a_7407_46529# a_7090_46419# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X11066 a_32334_61190# a_12981_59343# a_32826_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11067 a_41462_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11068 a_26495_35253# a_12381_35836# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11069 vcm_commonmode a_16362_14512# a_27406_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1107 a_12985_7663# a_12815_7663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11070 VDD a_12901_66665# a_44382_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11071 a_37446_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11072 VDD a_3705_73461# a_3595_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11073 a_23298_19898# a_11067_67279# a_23790_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11074 a_44474_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11075 a_27406_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11076 vcm_commonmode a_16362_67214# a_39454_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11077 a_20682_71230# a_12947_71576# a_20286_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11078 VDD a_11763_57399# a_11080_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X11079 a_43470_65206# a_16746_65208# a_43378_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1108 VDD a_1923_59583# a_2464_64605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X11080 a_7061_34319# a_6883_37019# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11081 a_11943_69367# a_12039_69367# a_12341_69455# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X11082 VDD a_1761_52815# a_12559_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11083 a_42374_20902# a_16362_20536# a_42466_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11084 a_27429_35301# a_27183_34789# a_28115_34743# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X11085 VDD a_12947_8725# a_25306_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11086 VSS a_12985_19087# a_21686_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11087 a_17366_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11088 a_31330_67214# a_12983_63151# a_31822_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11089 a_33430_57174# a_16746_57176# a_33338_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1109 a_21290_59182# a_16362_59182# a_21382_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11090 a_34738_18894# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11091 a_8289_15529# a_7841_12167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11092 vcm_commonmode a_16362_8488# a_38450_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11093 a_1761_44111# a_1591_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11094 a_7749_45577# a_6559_45205# a_7640_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11095 VSS a_6831_63303# a_30520_50345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11096 a_16362_67214# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11097 a_31726_8854# a_12947_8725# a_31330_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11098 VSS a_11151_14428# a_11082_14557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11099 a_46482_56170# a_16746_56172# a_46390_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X111 a_35765_29967# a_32970_31145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1110 a_8671_22671# a_4798_23759# a_8671_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=4.1e+11p ps=2.82e+06u w=1e+06u l=150000u
X11100 a_47790_17890# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11101 VDD a_1643_63125# a_1591_63151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11102 a_7921_26703# a_5085_23047# a_7837_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11103 VSS a_2292_43291# a_7337_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11104 a_29414_66210# a_16746_66212# a_29322_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11105 VDD a_1586_45431# a_9779_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X11106 a_31726_22910# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11107 VDD a_35815_31751# a_35431_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11108 a_18933_47741# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11109 a_28318_21906# a_16362_21540# a_28410_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1111 a_35742_24918# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11110 a_26319_38517# a_26495_38517# a_26447_38543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X11111 VDD a_15439_49525# a_38358_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11112 a_9405_10927# a_2004_42453# a_9187_10901# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11113 a_4333_22895# a_3985_22901# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11114 a_27710_61190# a_12355_15055# a_27314_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11115 VSS a_12899_10927# a_24698_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11116 VDD a_2824_70197# a_2960_70565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.226e+11p ps=2.21e+06u w=840000u l=150000u
X11117 a_21041_37429# a_18127_35797# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11118 a_49402_10862# a_16362_10496# a_49494_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11119 a_23298_8854# a_16362_8488# a_23390_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1112 VDD a_4443_46607# a_10299_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11120 a_39362_71230# a_12901_66665# a_39854_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11121 a_34434_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11122 VDD a_24800_44129# a_25388_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X11123 a_5411_59317# a_5091_60981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X11124 a_9835_69513# a_9319_69141# a_9740_69501# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X11125 a_3143_22364# a_2847_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11126 VDD a_23096_51017# a_23271_50943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11127 a_47486_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11128 a_49798_55166# VSS a_49402_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11129 a_3871_10383# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X1113 a_41766_17890# a_12899_11471# a_41370_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11130 VSS a_12899_11471# a_28714_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11131 a_25702_13874# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11132 a_5839_22351# a_5588_22467# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X11133 VDD config_2_in[13] a_1591_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11134 a_26402_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11135 a_37446_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11136 a_14939_31375# a_8197_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11137 a_2360_17277# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11138 vcm_commonmode a_16362_58178# a_46482_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11139 a_9557_57167# a_7155_55509# a_9123_57399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1114 a_6559_37583# a_6683_37815# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=0p ps=0u w=1e+06u l=150000u
X11140 a_29545_35841# a_29207_36415# a_30080_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11141 a_23390_8488# a_16746_8486# a_23298_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11142 a_37750_66210# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11143 a_8005_53333# a_7479_54439# a_8162_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11144 VDD a_2899_28111# a_3301_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11145 VSS a_11067_13095# a_41766_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11146 a_35346_23914# a_12947_23413# a_35838_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11147 a_29322_59182# a_12901_58799# a_29814_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11148 a_35346_19898# a_16362_19532# a_35438_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11149 a_22536_42919# a_21663_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1115 a_24698_69222# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11150 a_24194_35823# a_24017_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11151 vcm_commonmode a_16362_20536# a_39454_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11152 a_42374_65206# a_16362_65206# a_42466_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11153 a_48398_22910# a_10515_23975# a_48890_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11154 a_38358_55166# VSS a_38450_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11155 VSS a_12981_62313# a_27710_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11156 a_2203_21807# a_1757_21807# a_2107_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11157 a_9558_15101# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11158 VSS a_18848_27765# a_17358_31069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X11159 a_37446_71230# a_16746_71232# a_37354_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1116 a_30908_44869# a_31004_44869# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X11160 VDD a_12727_13353# a_32334_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11161 a_17670_69222# a_12516_7093# a_17274_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11162 a_3342_34639# a_2503_34319# a_3063_34319# VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=3.9975e+11p ps=3.83e+06u w=650000u l=150000u
X11163 a_31971_37737# a_32365_37692# a_32031_37683# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11164 VDD a_3668_56311# a_6743_54447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X11165 a_38358_14878# a_12877_14441# a_38850_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11166 VDD a_26495_42869# a_26319_42869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X11167 a_12921_39631# a_12651_39997# a_12831_39997# VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11168 a_33430_10496# a_16746_10494# a_33338_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11169 a_39362_18894# a_16362_18528# a_39454_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1117 a_31077_35307# a_26433_39631# a_30991_35307# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X11170 VDD a_12877_14441# a_45386_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11171 a_42866_12472# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11172 a_1643_54421# a_1846_54699# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11173 a_40366_13874# a_16362_13508# a_40458_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11174 VSS a_2375_29588# a_1895_30138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X11175 a_16362_20536# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11176 a_13067_38517# a_27219_44011# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11177 a_25798_22512# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11178 a_28699_48169# a_26397_51183# a_28607_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X11179 VDD a_17668_49007# a_17843_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1118 a_48794_23914# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11180 VSS a_5085_23047# a_5639_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11181 a_28108_48463# a_27929_48579# a_28192_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X11182 a_32426_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11183 a_6980_42479# a_6863_42692# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11184 VSS a_12355_65103# a_18674_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11185 a_42466_24552# VDD a_42374_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11186 a_38044_44759# a_38140_44501# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11187 VDD a_12899_11471# a_18278_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11188 VDD a_32649_28853# a_31768_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11189 a_32730_71230# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1119 a_11711_32143# a_9367_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X11190 a_5094_68413# a_2843_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11191 a_16362_18528# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11192 a_21831_51183# a_22164_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X11193 a_31422_69222# a_16746_69224# a_31330_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11194 a_46882_11468# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11195 VSS a_7061_34319# a_6372_38279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X11196 a_8369_25071# a_6162_28487# a_8297_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11197 a_36842_68540# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11198 a_30326_24918# VSS a_30418_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11199 VSS a_3714_58345# a_3509_58487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X112 vcm_commonmode a_16362_14512# a_37446_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1120 a_36392_43677# a_35647_42405# a_36520_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11200 a_29814_21508# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11201 VDD a_12983_63151# a_40366_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11202 VDD a_12755_51562# a_12587_51335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11203 a_29414_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11204 a_26310_14878# a_16362_14512# a_26402_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11205 a_5265_24643# a_5211_24759# a_5169_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11206 a_30418_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11207 VDD a_5147_50943# a_5134_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11208 a_4399_48084# a_4491_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11209 a_38315_38053# a_37076_37253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X1121 a_49494_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11210 a_4669_51005# a_4625_50613# a_4503_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11211 a_33338_60186# a_16362_60186# a_33430_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11212 VDD a_76648_40202# a_76461_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11213 a_32580_48783# a_14831_50095# a_32319_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11214 a_45478_15516# a_16746_15514# a_45386_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11215 a_23390_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11216 a_6180_69929# a_5438_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X11217 a_19774_13476# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11218 VDD a_12985_19087# a_34342_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11219 vcm_commonmode a_16362_65206# a_32426_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1122 a_37491_42359# a_37885_42333# a_37551_42333# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11220 VDD a_12985_16367# a_23298_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11221 a_1644_54965# a_1823_54973# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11222 a_41405_32463# a_11067_46823# a_41059_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X11223 a_37354_64202# a_11067_13095# a_37846_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11224 a_3983_50095# a_4031_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11225 a_41862_62516# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11226 a_32494_48463# a_17682_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X11227 a_2685_59933# a_1954_61677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11228 a_8500_58799# a_7871_59049# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11229 a_43445_28335# a_18979_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1123 a_8080_47607# a_8295_47388# a_8222_47414# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X11230 a_22294_9858# a_12546_22351# a_22786_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11231 VSS a_2473_34293# a_4263_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11232 vcm_commonmode a_16362_57174# a_22386_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11233 a_11299_62215# a_11145_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11234 a_49494_14512# a_16746_14510# a_49402_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11235 a_22132_44129# a_24331_44581# a_25204_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11236 VDD a_30485_49257# a_30928_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11237 vcm_commonmode a_16362_11500# a_46482_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11238 a_35517_34954# a_4443_46607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11239 a_32826_9460# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1124 a_39362_71230# a_16362_71230# a_39454_71230# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11240 a_45878_19500# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11241 VDD a_12727_67753# a_17274_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11242 a_40961_31375# a_33694_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11243 a_25879_48169# a_6835_46823# a_25961_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11244 VDD a_12257_56623# a_47394_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11245 VSS a_6372_38279# a_7526_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11246 a_4052_37961# a_2971_37589# a_3705_37557# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11247 VDD a_7162_59575# a_6382_61127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X11248 a_27806_63520# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11249 VDD a_12355_15055# a_31330_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1125 VSS a_1586_66567# a_10975_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11250 VDD a_11872_57711# a_12047_57685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11251 result_out[14] a_1644_74005# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X11252 a_11709_55777# a_11491_55535# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X11253 a_10189_60797# a_10145_60405# a_10023_60809# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11254 a_17670_22910# a_11067_21583# a_17274_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11255 a_20589_49917# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11256 a_40366_58178# a_16362_58178# a_40458_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11257 a_14013_30083# a_12935_31287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11258 a_23298_68218# a_16362_68218# a_23390_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11259 a_35438_64202# a_16746_64204# a_35346_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1126 a_25306_58178# a_16362_58178# a_25398_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11260 a_48890_8456# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11261 a_44778_8854# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11262 a_40366_17890# a_12899_10927# a_40858_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11263 VSS a_12947_23413# a_40762_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11264 a_37446_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11265 a_11803_55311# a_26267_43983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11266 a_38171_34191# a_37994_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11267 a_42224_38341# a_41351_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X11268 a_33734_18894# a_12899_10927# a_33338_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11269 VDD a_8969_42233# a_8999_41974# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1127 a_7187_20719# a_6743_20969# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X11270 VDD a_5915_30287# a_23309_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11271 a_31422_22544# a_16746_22542# a_31330_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11272 VSS a_23749_36929# a_24987_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11273 a_26310_59182# a_16362_59182# a_26402_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11274 vcm_commonmode a_16362_70226# a_40458_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11275 VSS a_24382_41629# a_24561_41583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11276 a_9759_49551# a_9135_49557# a_9651_49929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X11277 a_30418_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11278 a_19311_35823# a_19134_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11279 a_2012_44655# a_1778_42631# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1128 a_38754_15882# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11280 a_46786_17890# a_12899_11471# a_46390_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11281 a_44382_16886# a_12899_11471# a_44874_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11282 a_29718_69222# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11283 VSS a_10472_26159# a_11074_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11284 a_30722_64202# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11285 a_21829_48161# a_21611_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X11286 a_31669_51183# a_2959_47113# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11287 a_26779_50461# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11288 VSS a_12877_14441# a_34738_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11289 VDD a_8079_43732# a_6863_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1129 vcm_commonmode a_16362_71230# a_21382_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11290 VDD a_2952_66139# a_7387_66781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11291 a_11866_27791# a_7369_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11292 vcm_commonmode a_16362_61190# a_43470_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11293 VSS a_21049_34717# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X11294 VSS a_12901_58799# a_23694_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11295 a_20682_56170# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11296 a_17274_18894# a_12895_13967# a_17766_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11297 VSS VSS a_17670_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11298 VSS a_13015_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X11299 vcm_commonmode a_16362_71230# a_26402_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X113 a_46390_16886# a_12899_11471# a_46882_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1130 a_45782_16886# a_12727_13353# a_45386_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11300 a_21782_16488# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11301 VSS a_12727_15529# a_47790_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11302 a_15793_28585# a_15315_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11303 VDD a_5671_21495# a_11887_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11304 VDD a_12947_71576# a_38358_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11305 VDD VDD a_39362_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11306 VSS VDD a_35742_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11307 vcm_commonmode a_16362_10496# a_22386_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11308 a_9431_60214# a_6417_62215# a_9359_60214# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11309 a_31330_12870# a_12877_16911# a_31822_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1131 a_27195_32375# a_26985_31605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11310 a_2307_31965# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11311 a_38450_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11312 a_7467_61751# a_8039_61493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11313 a_20378_61190# a_16746_61192# a_20286_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11314 vcm_commonmode a_16362_60186# a_47486_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11315 a_6646_54135# a_5254_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X11316 vcm_commonmode a_16362_19532# a_47486_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11317 a_28902_28335# a_13643_28327# a_28733_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11318 a_27314_7850# VDD a_27806_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11319 a_24698_55166# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1132 VDD a_11803_55311# a_16746_61192# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X11320 a_1933_5059# a_1761_2767# a_1861_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11321 a_8219_54447# a_7210_55081# a_8082_54599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11322 a_24698_13874# a_12877_16911# a_24302_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11323 vcm_commonmode VSS a_31422_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11324 a_1945_16911# a_1908_17141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11325 a_33734_7850# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11326 a_49798_63198# a_15439_49525# a_49402_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11327 a_25306_68218# a_12727_67753# a_25798_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11328 a_36746_66210# a_12983_63151# a_36350_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11329 a_2319_59317# a_2124_59459# a_2629_59709# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X1133 VSS a_12727_15529# a_42770_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11330 a_33430_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11331 a_24394_60186# a_16746_60188# a_24302_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11332 a_24394_19532# a_16746_19530# a_24302_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11333 VDD a_10515_23975# a_34342_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11334 VDD a_12727_58255# a_28318_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11335 vcm_commonmode a_16362_16520# a_21382_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11336 a_12381_43957# a_37799_43777# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X11337 VDD a_11964_71855# a_12139_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11338 VDD a_1775_60663# a_1775_60439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X11339 VDD a_8896_65015# a_8453_64757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1134 a_11985_69455# a_11943_69367# a_10747_68565# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X11340 a_42715_29423# a_41597_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X11341 VSS VDD a_41766_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11342 VSS a_7676_61493# a_7622_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11343 VDD a_5336_54965# a_5274_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11344 VSS a_2111_38279# a_2052_38377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X11345 a_16928_36391# a_15959_36415# a_16832_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11346 a_29322_67214# a_12983_63151# a_29814_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11347 VDD a_35493_43421# a_35099_43447# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11348 VSS a_4298_58951# a_8133_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X11349 a_30326_62194# a_12355_15055# a_30818_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1135 a_10403_48285# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11350 a_35438_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11351 a_2104_52271# a_1987_52484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11352 a_11599_65693# a_10975_65327# a_11491_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X11353 VDD a_15074_50871# a_14681_50247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X11354 a_38358_63198# a_16362_63198# a_38450_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11355 a_20682_7850# VDD a_20286_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11356 VSS a_25493_29967# a_26612_29473# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X11357 a_35039_51335# a_29361_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11358 a_23790_57496# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11359 VDD a_2672_15113# a_2847_15039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1136 VDD a_12947_71576# a_33338_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11360 a_29718_22910# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11361 vcm_commonmode a_16362_68218# a_37446_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11362 a_37446_7484# VDD a_37354_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11363 VSS a_7439_64213# a_7387_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11364 VSS a_1925_22583# a_1738_22325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11365 a_11711_12559# a_10753_12559# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11366 a_40049_27497# a_18979_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11367 a_4061_40079# a_3305_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X11368 VSS a_2292_43291# a_5313_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11369 a_31726_71230# a_12947_71576# a_31330_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1137 a_25306_17890# a_12899_10927# a_25798_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11370 VDD a_4482_57863# a_33515_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11371 VDD a_22062_31287# a_21273_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11372 VSS a_12877_16911# a_23694_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11373 VDD a_16043_38825# a_16556_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X11374 VSS a_10506_29967# a_14939_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11375 a_6327_34863# a_5691_36727# a_5964_35015# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11376 vcm_commonmode a_16362_9492# a_18370_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11377 a_31280_36165# a_30311_35877# a_31243_35831# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X11378 a_2215_69135# a_1591_69141# a_2107_69513# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11379 VDD a_1643_56597# a_1591_56623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1138 VSS a_12947_23413# a_25702_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11380 a_13743_35836# a_18811_34789# a_19684_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11381 VSS a_12355_15055# a_48794_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11382 a_3421_57167# a_3295_62083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11383 a_12723_14191# a_11067_63143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11384 VSS a_28883_52031# a_28817_52105# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X11385 a_44474_57174# a_16746_57176# a_44382_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11386 a_45782_18894# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11387 a_8373_26409# a_3607_34639# a_8289_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11388 a_2319_59317# a_2163_59585# a_2464_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X11389 a_40233_31605# a_8491_41383# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1139 a_25447_34743# a_12713_36483# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X11390 a_27406_67214# a_16746_67216# a_27314_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11391 a_32584_50639# a_29361_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X11392 VSS a_17039_51157# a_16997_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11393 a_33830_22512# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11394 a_14289_29687# a_13239_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11395 a_26310_22910# a_16362_22544# a_26402_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11396 a_22386_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11397 VDD a_12355_65103# a_36350_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11398 a_7571_20291# a_7377_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X11399 a_8126_46287# a_7368_46403# a_7563_46261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 VSS a_2223_28617# a_2981_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X1140 a_33430_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11400 a_30418_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11401 a_16746_18526# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11402 a_9135_29423# a_7841_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X11403 a_33741_32463# a_29927_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11404 a_7203_24527# a_4571_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.1275e+11p pd=3.87e+06u as=0p ps=0u w=650000u l=150000u
X11405 a_18674_61190# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11406 a_17366_59182# a_16746_59184# a_17274_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11407 VDD a_15439_49525# a_49402_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11408 a_6559_72512# a_6327_72917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X11409 a_20286_71230# a_16362_71230# a_20378_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1141 a_31787_36919# a_32181_36893# a_31847_36893# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11410 a_25702_62194# a_12981_62313# a_25306_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11411 a_31422_29423# a_22843_29415# a_31127_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11412 a_24541_47741# a_24497_47349# a_24375_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11413 a_2012_9839# a_1867_10927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X11414 a_12591_31029# a_8461_32937# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11415 VSS a_12895_13967# a_22690_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11416 a_11812_30511# a_11183_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X11417 a_8364_44655# a_7295_44647# a_8143_44982# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11418 a_37354_72234# VDD a_37846_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11419 VSS a_4771_56597# a_1823_66941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1142 vcm_commonmode a_16362_8488# a_20378_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11420 a_41862_70548# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11421 a_34342_14878# a_16362_14512# a_34434_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11422 VDD a_3143_22364# a_4139_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11423 a_31648_43781# a_30679_43493# a_31552_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11424 a_11311_74005# a_11136_74031# a_11490_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11425 a_37846_60508# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11426 a_45478_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11427 vcm_commonmode VSS a_18370_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11428 VDD a_2672_49929# a_2847_49855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11429 a_24302_70226# a_16362_70226# a_24394_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1143 a_16362_71230# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11430 a_3026_36861# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11431 a_23694_14878# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11432 a_7799_46831# a_6835_46823# a_7436_46983# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11433 VSS a_1950_59887# a_3983_68591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11434 a_1853_27247# a_1683_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11435 VDD a_4685_37583# a_8332_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11436 VSS a_4035_54965# a_1823_58773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11437 a_27806_71552# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11438 a_35742_67214# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11439 VSS a_12473_37429# a_27415_36341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1144 vcm_commonmode a_16362_60186# a_42466_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11440 VDD a_12985_19087# a_42374_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11441 VDD a_11067_67279# a_27314_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11442 a_42770_68218# a_12901_66959# a_42374_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11443 a_26631_35877# a_25484_37253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X11444 a_4653_60797# a_4274_60431# a_4581_60797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11445 a_27314_61190# a_16362_61190# a_27406_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11446 a_48794_66210# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11447 VSS a_7901_13077# a_7797_13885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X11448 vcm_commonmode a_16362_21540# a_37446_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11449 a_46390_23914# a_12947_23413# a_46882_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1145 a_46882_59504# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11450 a_46390_19898# a_16362_19532# a_46482_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11451 VDD a_10055_58791# a_17274_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11452 a_1757_9839# a_1591_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11453 VDD a_5993_32687# a_7067_30663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11454 a_24556_49551# a_23830_49525# a_7479_54439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X11455 VDD a_15968_36061# a_15069_35805# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X11456 VSS a_27869_50095# a_29364_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11457 a_35438_72234# VDD a_35346_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11458 a_45782_59182# a_12727_58255# a_45386_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11459 VSS a_12947_56817# a_42770_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1146 a_18674_18894# a_12899_10927# a_18278_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11460 a_39854_18496# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11461 a_36350_15882# a_12727_13353# a_36842_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11462 a_28410_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11463 a_39758_24918# VSS a_39362_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11464 VDD a_12727_13353# a_43378_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11465 a_40858_13476# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11466 a_28714_69222# a_12516_7093# a_28318_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11467 VSS a_10975_66407# a_25702_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11468 a_6980_49917# a_6863_49722# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11469 a_37512_50755# a_36821_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1147 vcm_commonmode a_16362_19532# a_42466_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11470 a_14524_48437# a_11067_13095# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=0p ps=0u w=650000u l=150000u
X11471 a_44474_10496# a_16746_10494# a_44382_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11472 VSS a_2411_18517# a_6141_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11473 a_76365_39738# a_76461_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11474 a_37951_42089# a_38345_42044# a_38011_42035# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11475 VSS a_7436_46983# a_7387_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11476 VDD a_2411_18517# a_11296_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11477 a_27406_20536# a_16746_20534# a_27314_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11478 a_30418_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11479 a_40366_9858# a_16362_9492# a_40458_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1148 a_23309_31849# a_5915_35943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X11480 VSS a_13576_40413# a_12677_40157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X11481 VSS a_4119_70741# a_4065_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11482 a_44382_67214# a_16362_67214# a_44474_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11483 VSS VSS a_46786_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11484 a_30722_72234# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11485 VDD a_32327_40191# a_32187_40513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11486 a_41443_41855# a_38011_42035# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X11487 VSS a_12355_65103# a_29718_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11488 a_8630_48463# a_7553_48469# a_8468_48841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11489 a_34834_69544# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1149 vcm_commonmode a_16362_70226# a_25398_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11490 a_17366_12504# a_16746_12502# a_17274_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11491 VDD a_12899_11471# a_29322_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11492 a_27406_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11493 a_16746_63200# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11494 a_34342_59182# a_16362_59182# a_34434_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11495 a_47886_68540# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11496 a_26402_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11497 a_22536_41831# a_21663_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11498 a_6094_67825# a_3143_66972# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11499 a_16746_10494# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X115 a_7005_55223# a_7210_55081# a_7168_55107# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1150 a_30418_8488# a_16746_8486# a_30326_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11500 a_14859_37737# a_14919_37683# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11501 a_17274_69222# a_16362_69222# a_17366_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11502 VSS a_12257_56623# a_19678_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11503 a_18539_47617# a_4191_33449# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11504 VDD config_2_in[0] a_1591_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11505 a_39771_31375# a_35815_31751# a_13643_28327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X11506 a_21479_36965# a_20713_36929# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X11507 a_21382_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11508 a_11599_61341# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11509 a_23694_55166# VSS a_23298_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1151 a_32612_51727# a_33360_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.8668e+12p pd=1.774e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X11510 a_7992_17277# a_7649_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11511 a_5601_11471# a_5199_11791# a_5437_11791# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X11512 a_12901_66959# a_11067_67279# a_12901_67279# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11513 a_35346_65206# a_12355_65103# a_35838_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11514 a_5225_52271# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11515 a_38499_42943# a_36432_42919# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X11516 VDD a_12901_66959# a_24302_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11517 a_48398_64202# a_11067_13095# a_48890_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11518 VDD a_6066_28309# a_6809_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11519 VSS a_6066_28309# a_6559_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1152 a_34391_48682# a_34221_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11520 a_24698_63198# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11521 VSS a_10391_67477# a_10325_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11522 vcm_commonmode a_16362_58178# a_20378_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11523 vcm_commonmode a_16362_71230# a_34434_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11524 a_4941_35727# a_1915_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11525 a_35742_20902# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11526 VSS a_12947_23413# a_38754_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11527 vcm_commonmode a_16362_57174# a_33430_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11528 a_9184_49159# a_9392_48981# a_9326_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X11529 a_42770_21906# a_12985_7663# a_42374_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1153 VDD a_12901_66665# a_37354_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11530 VSS a_19596_40743# a_19559_41001# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11531 a_22084_49007# a_21003_49007# a_21737_49249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11532 a_38358_56170# a_12947_56817# a_38850_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11533 VDD a_15009_47919# a_15617_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X11534 VDD a_10515_22671# a_45386_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11535 a_9794_51549# a_9707_51325# a_9390_51435# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X11536 VSS a_7467_57863# a_6880_58773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X11537 a_22294_22910# a_10515_23975# a_22786_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11538 VSS a_29927_29199# a_36264_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11539 VDD a_12591_31029# a_12120_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1154 a_29322_16886# a_12899_11471# a_29814_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11540 VDD a_12727_67753# a_28318_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11541 a_25798_64524# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11542 a_40343_37737# a_40737_37692# a_40403_37683# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11543 a_2215_51549# a_1923_54591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11544 VDD VDD a_47394_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11545 VSS VDD a_43774_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11546 VDD a_2235_30503# a_25321_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11547 a_32730_13874# a_12877_16911# a_32334_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11548 ctopn a_3339_43023# ctopn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u M=2
X11549 a_28410_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1155 VDD a_11617_18785# a_11507_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X11550 a_36746_9858# a_12985_19087# a_36350_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11551 a_3026_26159# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11552 a_10492_60809# a_9411_60437# a_10145_60405# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11553 a_45782_12870# a_10055_58791# a_45386_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11554 a_8325_18517# a_6816_19355# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11555 a_28714_22910# a_11067_21583# a_28318_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11556 a_6095_44807# a_7815_45503# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11557 a_5239_48767# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11558 VSS a_1586_51335# a_11711_50645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11559 VSS a_12516_7093# a_37750_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1156 a_44778_63198# a_15439_49525# a_44382_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11560 a_30326_70226# a_12516_7093# a_30818_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11561 a_24698_9858# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11562 VSS a_26417_40193# a_26919_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X11563 VSS a_1586_51335# a_1683_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11564 a_26310_60186# a_12727_58255# a_26802_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11565 a_12231_55509# a_12056_55535# a_12410_55535# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11566 a_35438_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11567 a_8782_65015# a_11771_68021# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=0p ps=0u w=650000u l=150000u
X11568 a_32401_46831# a_22843_29415# a_28756_55394# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11569 vcm_commonmode a_16362_15516# a_42466_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1157 a_30326_11866# a_10055_58791# a_30818_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11570 a_4095_29423# a_1915_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X11571 a_19774_55488# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11572 a_6914_14735# a_4629_13647# a_6611_14967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11573 a_29322_12870# a_12877_16911# a_29814_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11574 VSS a_13357_32143# a_26157_31605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11575 a_30127_38053# a_29361_38017# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X11576 VDD a_29545_40193# a_29804_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11577 a_9863_51420# a_9707_51325# a_10008_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X11578 a_42466_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11579 a_45386_7850# VSS a_45478_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1158 VDD a_37939_43455# a_37799_43777# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11580 a_44778_18894# a_12899_10927# a_44382_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11581 a_3605_13647# a_3023_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11582 a_10969_71631# a_2451_72373# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11583 a_13909_35395# a_18627_35327# a_19500_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11584 a_18370_61190# a_16746_61192# a_18278_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11585 VSS a_7039_65469# a_7000_65595# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11586 a_31898_30761# a_30790_30663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=9.65e+11p pd=7.93e+06u as=0p ps=0u w=1e+06u l=150000u
X11587 VSS a_12727_67753# a_31726_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11588 a_4433_26703# a_4151_28879# a_4351_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11589 a_10097_62973# a_10053_62581# a_9931_62985# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1159 a_20286_68218# a_12727_67753# a_20778_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11590 VSS a_12985_16367# a_19678_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11591 a_9221_15279# a_2004_42453# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11592 a_42374_19898# a_11067_67279# a_42866_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11593 vcm_commonmode VSS a_29414_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11594 a_10747_16950# a_5535_18012# a_10288_17143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11595 vcm_commonmode a_16362_62194# a_41462_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11596 VSS a_2847_36799# a_2781_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X11597 a_46482_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11598 VSS a_12877_14441# a_45782_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11599 a_4893_33821# a_1915_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X116 a_7377_18012# a_12139_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X1160 inn_analog a_3339_43023# ctopn VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7645e+12p ps=2.191e+07u w=1.9e+06u l=220000u M=4
X11600 a_24302_63198# a_12981_62313# a_24794_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11601 a_6829_15055# a_5399_13255# a_6611_14967# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11602 vcm_commonmode a_16362_16520# a_19374_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11603 a_31726_56170# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11604 a_28318_18894# a_12895_13967# a_28810_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11605 VDD VDD a_36350_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11606 VDD a_12947_8725# a_19282_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11607 a_5915_35943# a_15681_27497# a_21490_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X11608 a_23390_14512# a_16746_14510# a_23298_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11609 vcm_commonmode a_16362_11500# a_20378_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1161 VDD a_12727_58255# a_23298_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11610 a_26694_29473# a_2787_30503# a_26612_29473# VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X11611 a_2011_34837# a_4903_29975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11612 a_32826_16488# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11613 a_31330_8854# a_12985_19087# a_31822_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11614 a_3016_60949# a_4864_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11615 a_7939_27497# a_3301_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X11616 VDD a_2686_70223# a_7755_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.99e+12p ps=2.398e+07u w=1e+06u l=150000u M=4
X11617 a_2928_22583# a_2315_24540# a_3070_22717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11618 VDD a_33656_43439# a_33762_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11619 a_36442_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1162 VDD a_5013_20473# a_5043_20214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11620 VDD a_12947_71576# a_49402_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11621 a_8739_28879# a_8206_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11622 a_8001_40125# a_7373_40847# a_7929_40125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11623 a_25388_43781# a_24515_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11624 a_14131_44135# a_3339_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11625 vcm_commonmode a_16362_10496# a_33430_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11626 a_19374_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11627 a_2007_39978# a_2052_38377# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X11628 VDD a_13835_41001# a_13980_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11629 a_49494_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1163 VSS a_12877_14441# a_19678_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11630 VDD a_18695_47349# a_18626_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11631 a_23553_31171# a_15548_30761# a_23481_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11632 a_34342_22910# a_16362_22544# a_34434_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11633 a_3828_15823# a_3391_15797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11634 VDD a_4903_31849# a_10045_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11635 a_48490_66210# a_16746_66212# a_48398_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11636 VSS a_13984_43781# a_13947_43447# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11637 VDD a_12447_29199# a_40139_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X11638 a_23298_69222# a_12901_66959# a_23790_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11639 a_47394_21906# a_16362_21540# a_47486_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1164 vcm_commonmode a_16362_61190# a_28410_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11640 a_34738_67214# a_12727_67753# a_34342_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11641 vcm_commonmode a_16362_63198# a_18370_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11642 VDD a_1643_72917# a_1591_72943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11643 a_2163_64381# a_1586_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11644 a_2325_44897# a_2107_44655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X11645 a_15439_49525# a_15575_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11646 VDD a_11521_66567# a_11613_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X11647 a_8753_19319# a_5535_18012# a_8916_19203# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11648 VSS a_16265_39868# a_15957_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11649 a_7808_48829# a_7557_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1165 VSS a_35959_30485# a_22015_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u M=2
X11650 a_8325_18517# a_6816_19355# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11651 VSS a_12899_10927# a_43774_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11652 a_4788_45565# a_4758_45369# a_4308_45431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11653 a_28195_35327# a_27429_35301# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X11654 a_22399_32143# a_22148_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X11655 a_5823_44905# a_5173_44655# a_5905_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11656 a_24394_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11657 a_6649_25615# a_5211_24759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11658 VSS a_2011_34837# a_1969_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X11659 VSS a_3203_17620# a_1895_18756# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1166 VSS a_2479_50899# a_1923_54591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X11660 VSS a_2319_57948# a_2250_58077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11661 a_10761_29745# a_8485_29673# a_10689_29745# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11662 a_30943_38695# a_1761_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X11663 a_20682_17890# a_12899_11471# a_20286_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11664 a_44778_13874# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11665 a_24768_27247# a_9529_28335# a_24683_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X11666 a_2041_61519# a_1954_61677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11667 a_9526_61751# a_9431_60214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11668 a_6649_37289# a_4685_37583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11669 a_27710_23914# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1167 a_10055_58791# a_7000_43541# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X11670 a_4035_11989# a_3327_9308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11671 a_17366_8488# a_16746_8486# a_17274_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11672 VSS a_11067_21583# a_31726_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11673 a_28410_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11674 a_39454_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11675 VSS a_2007_39978# a_1778_42631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X11676 VSS a_34943_51335# a_34411_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11677 a_36350_66210# a_16362_66210# a_36442_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11678 VDD a_5612_58229# a_5550_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11679 a_37195_47919# a_16863_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1168 a_7467_61751# a_8039_61493# a_7812_61839# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X11680 VDD a_13692_34191# a_13798_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11681 a_9366_14735# a_8289_14741# a_9204_15113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X11682 vcm_commonmode a_16362_68218# a_48490_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11683 a_16746_59184# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X11684 VSS a_35683_50613# a_35495_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11685 a_17280_48695# a_17488_48731# a_17422_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X11686 a_17670_15882# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11687 a_49402_9858# a_16362_9492# a_49494_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11688 a_12082_25077# a_9751_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11689 VSS a_12727_15529# a_21686_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1169 a_8762_36815# a_7749_37903# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11690 a_2107_26159# a_1591_26159# a_2012_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X11691 a_24638_49871# a_23774_49551# a_7479_54439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X11692 a_4948_63695# a_4734_63695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X11693 a_4458_45565# a_2927_39733# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11694 a_28814_50345# a_4351_67279# a_28730_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11695 VSS a_12981_62313# a_46786_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11696 a_43774_60186# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11697 a_42466_58178# a_16746_58180# a_42374_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11698 a_43774_19898# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11699 a_76971_38925# a_76346_40594# VSS VDD sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=4.74e+06u as=0p ps=0u w=500000u l=500000u M=2
X117 a_39362_7850# VDD a_39854_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1170 a_75794_38962# a_75628_38962# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X11700 a_43624_30287# a_18979_30287# a_43321_29941# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11701 VSS a_10975_66407# a_33734_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11702 a_26706_70226# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11703 a_25398_68218# a_16746_68220# a_25306_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11704 VSS a_32795_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X11705 a_26319_36341# a_12641_36596# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11706 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11707 a_16746_71232# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11708 VDD a_10975_66407# a_34342_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11709 VSS a_2511_42479# a_2292_43291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X1171 a_32426_18528# a_16746_18526# a_32334_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11710 VSS a_1923_54591# a_4549_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11711 VSS a_35739_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X11712 a_44874_22512# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11713 a_38067_47349# a_29927_29199# a_38213_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11714 a_34434_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11715 a_23694_63198# a_15439_49525# a_23298_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11716 VSS a_12727_58255# a_20682_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11717 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11718 VDD a_26319_37429# a_16152_37601# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11719 VSS a_11067_67279# a_20682_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1172 a_1920_59861# a_2099_59861# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11720 VDD a_1923_54591# a_10008_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11721 VDD a_19127_43439# a_19233_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11722 a_11661_18543# a_11617_18785# a_11495_18543# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11723 VSS a_2847_26133# a_2781_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11724 VDD a_12899_11471# a_37354_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11725 a_34834_14480# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11726 a_31330_71230# a_16362_71230# a_31422_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11727 a_34738_20902# a_11067_67279# a_34342_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11728 a_17766_24520# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11729 a_8682_42301# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1173 a_5607_44343# a_4443_46607# a_5781_44449# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11730 a_48398_72234# VDD a_48890_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11731 VDD a_11067_21583# a_21290_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11732 a_18045_41281# a_17983_41855# a_18856_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11733 VSS a_7387_64239# a_7758_65693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11734 a_48890_21508# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11735 a_6106_35190# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X11736 a_25091_37782# a_24413_39087# a_25019_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11737 a_48490_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11738 a_45386_14878# a_16362_14512# a_45478_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11739 a_19967_41781# a_52778_39936# a_53570_39250# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=0p ps=0u w=800000u l=150000u
X1174 VDD a_4351_67279# a_8675_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X11740 a_6980_49917# a_6863_49722# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11741 a_3749_73853# a_3705_73461# a_3583_73865# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X11742 a_3355_25071# a_3104_25321# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X11743 a_38850_13476# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11744 a_35346_10862# a_12985_16367# a_35838_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11745 VDD a_3759_39991# a_3663_39991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11746 VDD a_12985_16367# a_42374_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11747 a_27710_64202# a_12355_65103# a_27314_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11748 VDD a_12901_66959# a_32334_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11749 a_18278_20902# a_12985_7663# a_18770_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1175 a_24302_67214# a_12983_63151# a_24794_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11750 a_18278_16886# a_16362_16520# a_18370_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11751 a_11151_14428# a_10956_14459# a_11461_14191# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X11752 a_25798_72556# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11753 a_3107_53359# a_2177_53359# a_2744_53511# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X11754 VDD a_12985_7663# a_25306_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11755 a_22386_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11756 a_49402_13874# a_16362_13508# a_49494_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11757 a_28410_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11758 a_25306_62194# a_16362_62194# a_25398_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11759 a_46786_67214# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1176 a_40773_30511# a_12447_29199# a_40691_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11760 a_37446_17524# a_16746_17522# a_37354_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11761 a_17670_56170# a_12257_56623# a_17274_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11762 VDD a_1803_19087# a_1945_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11763 vcm_commonmode a_16362_67214# a_24394_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11764 VDD a_3247_20495# a_7153_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X11765 vcm_commonmode a_16362_21540# a_48490_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11766 a_33830_64524# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11767 a_36746_59182# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11768 VDD a_10055_58791# a_28318_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11769 a_2215_23439# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1177 a_2107_36873# a_1757_36501# a_2012_36861# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11770 VSS a_12257_56623# a_40762_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11771 a_26402_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11772 a_46882_63520# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11773 a_10705_68841# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X11774 vcm_commonmode a_16362_13508# a_38450_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11775 a_11048_29423# a_6459_30511# a_10825_29688# VSS sky130_fd_pr__nfet_01v8 ad=1.323e+11p pd=1.47e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11776 a_42466_11500# a_16746_11498# a_42374_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11777 VSS a_14049_40693# a_13983_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11778 VSS a_6269_43567# a_6661_42255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11779 VSS a_1761_25071# a_32695_43455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1178 a_35742_65206# a_10975_66407# a_35346_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11780 a_31422_56170# a_16746_56172# a_31330_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11781 a_32730_17890# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11782 VDD a_12895_13967# a_41370_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11783 a_25398_21540# a_16746_21538# a_25306_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11784 VSS a_4676_47607# a_4491_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11785 a_34342_60186# a_12727_58255# a_34834_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11786 a_38754_8854# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11787 a_42374_68218# a_16362_68218# a_42466_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11788 VDD a_75445_39738# a_75258_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11789 VDD a_34759_31029# a_36001_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1179 a_33727_44265# a_32795_44031# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X11790 VDD a_11311_74005# a_11298_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11791 VDD a_15439_49525# a_23298_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11792 a_6676_69455# a_5924_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11793 VDD a_29072_38567# a_28976_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X11794 VSS a_32970_31145# a_40323_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X11795 a_45878_69544# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11796 a_11780_69679# a_10699_69679# a_11433_69921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11797 VSS a_10515_22671# a_17670_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11798 a_24302_71230# a_12901_66665# a_24794_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11799 a_45386_59182# a_16362_59182# a_45478_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X118 VDD a_4891_47388# a_22921_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X1180 a_40491_27247# a_40218_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11800 a_8636_63669# a_7155_55509# a_9028_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X11801 a_28318_69222# a_16362_69222# a_28410_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11802 a_25091_37455# a_24837_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11803 VDD a_12981_62313# a_27314_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11804 a_32426_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11805 a_46390_65206# a_12355_65103# a_46882_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11806 a_19410_43439# a_19233_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X11807 a_9184_13255# a_7841_12167# a_9326_13103# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X11808 a_41862_8456# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11809 a_13143_29575# a_13241_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X1181 a_4036_51157# a_4215_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11810 a_12965_27791# a_12631_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X11811 a_22386_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11812 a_49402_58178# a_16362_58178# a_49494_58178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11813 VSS a_19596_34215# a_19559_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11814 VSS VSS a_36746_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11815 vcm_commonmode a_16362_58178# a_31422_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11816 vcm_commonmode a_16362_71230# a_45478_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11817 VSS a_2872_44111# a_19113_51005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11818 a_22690_66210# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11819 a_36350_57174# a_12257_56623# a_36842_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1182 a_48794_64202# a_12355_65103# a_48398_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11820 a_40858_55488# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11821 a_49402_17890# a_12899_10927# a_49894_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11822 VSS a_12947_23413# a_49798_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11823 a_46786_20902# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11824 a_20286_23914# a_12947_23413# a_20778_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11825 a_20286_19898# a_16362_19532# a_20378_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11826 a_9989_46831# a_9821_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X11827 VDD a_12947_8725# a_27314_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11828 VSS a_12985_19087# a_23694_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11829 vcm_commonmode a_16362_20536# a_24394_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1183 VDD a_2451_72373# a_2882_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11830 a_7624_68021# a_7155_55509# a_8016_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X11831 VDD a_29361_38017# a_29620_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11832 a_33338_22910# a_10515_23975# a_33830_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11833 a_26402_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11834 a_23298_55166# VSS a_23390_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11835 VSS a_12727_13353# a_39758_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11836 a_12793_35862# a_12621_36091# a_12579_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X11837 a_36746_12870# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11838 a_22386_71230# a_16746_71232# a_22294_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11839 vcm_commonmode a_16362_70226# a_49494_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1184 vcm_commonmode a_16362_14512# a_33430_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11840 a_2295_17429# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X11841 a_43774_13874# a_12877_16911# a_43378_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11842 VSS a_12985_16367# a_40762_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11843 VDD a_3693_68047# a_5060_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11844 a_3510_70223# a_3280_70501# a_2824_70197# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11845 VDD a_15095_41781# a_15009_40193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11846 a_26802_17492# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11847 a_23298_14878# a_12877_14441# a_23790_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11848 a_26706_23914# a_10515_23975# a_26310_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11849 a_27219_44011# a_12357_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1185 VDD a_12985_7663# a_46390_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11850 a_24302_18894# a_16362_18528# a_24394_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11851 a_10870_31599# a_8273_42479# a_10784_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11852 VDD a_12877_14441# a_30326_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11853 a_7170_21263# a_5535_18012# a_7086_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.8e+11p pd=2.76e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11854 VSS a_9307_30663# a_11048_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11855 a_44382_68218# a_12727_67753# a_44874_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11856 vcm_commonmode a_16362_62194# a_39454_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11857 a_21101_31055# a_5915_35943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11858 a_43470_60186# a_16746_60188# a_43378_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11859 a_8268_35381# a_4685_37583# a_8397_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X1186 a_2007_65002# a_2099_64757# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X11860 VDD a_12727_58255# a_47394_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11861 vcm_commonmode a_16362_16520# a_40458_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11862 a_43470_19532# a_16746_19530# a_43378_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11863 a_36116_50959# a_35676_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11864 a_22026_27247# a_17222_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X11865 a_26402_70226# a_16746_70228# a_26310_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11866 VDD a_4809_18785# a_4699_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11867 VDD a_11855_51959# a_11759_51959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11868 a_29718_56170# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11869 a_27314_13874# a_12727_15529# a_27806_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1187 a_26610_49257# a_6831_63303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X11870 VDD config_1_in[2] a_1591_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11871 a_40458_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11872 a_16556_39429# a_15683_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11873 a_31822_11468# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11874 VDD a_5964_67655# a_5167_68060# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11875 a_25306_8854# a_16362_8488# a_25398_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11876 a_21782_68540# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11877 a_20286_7850# VDD a_20778_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11878 a_16362_62194# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X11879 a_5039_42167# a_5098_41641# a_5962_41391# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X1188 a_12381_43957# a_37799_43777# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11880 a_5105_47673# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11881 a_17766_58500# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11882 VSS a_13975_44527# a_14081_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11883 a_5987_16733# a_5363_16367# a_5879_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11884 VSS a_10055_58791# a_17670_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11885 a_29414_61190# a_16746_61192# a_29322_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11886 VDD VSS a_39362_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11887 vcm_commonmode a_16362_17524# a_26402_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11888 a_30818_7452# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11889 a_18627_35327# a_15011_34717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X1189 a_24698_22910# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11890 VDD a_21233_40956# a_20839_41001# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11891 a_30418_15516# a_16746_15514# a_30326_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11892 VDD a_39468_37479# a_39372_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X11893 result_out[4] a_1644_58773# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X11894 a_2742_42997# a_2592_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.184e+11p pd=2.2e+06u as=0p ps=0u w=840000u l=150000u
X11895 a_7107_65871# a_6927_65871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11896 a_17803_36649# a_18197_36604# a_17863_36595# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X11897 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X11898 a_22294_64202# a_11067_13095# a_22786_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11899 a_9865_68047# a_10010_68021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X119 VSS a_15253_37692# a_14945_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X1190 a_9135_27239# a_41334_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X11900 a_24800_41953# a_24331_40767# a_25204_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11901 VSS a_2794_62697# a_2589_62839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11902 VSS a_9624_65301# a_10301_66237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11903 a_34434_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11904 VDD a_2969_41909# a_2859_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11905 a_22436_51005# a_10503_52828# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11906 a_8836_74953# a_7755_74581# a_8489_74549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11907 vcm_commonmode a_16362_11500# a_31422_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11908 a_14005_50959# a_12993_50345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11909 VSS a_23901_35516# a_23593_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1191 a_49494_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11910 a_34738_70226# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11911 a_33430_68218# a_16746_68220# a_33338_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11912 a_47486_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11913 VDD a_7159_22583# a_7111_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X11914 a_30818_19500# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11915 a_13795_37782# a_13613_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11916 VSS a_4001_56377# a_3935_56445# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11917 a_7479_17607# a_7407_18038# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11918 a_9651_49929# a_9135_49557# a_9556_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X11919 a_4065_25321# a_2315_24540# a_3983_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1192 a_46390_62194# a_16362_62194# a_46482_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11920 VSS a_29175_28335# a_41599_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X11921 a_46482_67214# a_16746_67216# a_46390_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11922 VDD a_12546_22351# a_34342_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11923 vcm_commonmode a_16362_64202# a_43470_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11924 VSS a_27245_41829# a_27747_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11925 a_9913_67503# a_9869_67745# a_9747_67503# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11926 a_45386_22910# a_16362_22544# a_45478_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11927 a_23498_28585# a_14926_31849# a_23385_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X11928 a_1642_18231# a_1738_17973# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11929 VDD a_11053_62607# a_11909_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1193 a_7376_59343# a_6737_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X11930 VSS a_27429_35301# a_28115_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X11931 a_37750_61190# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11932 a_4161_30761# a_3325_29967# a_4065_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X11933 a_36442_59182# a_16746_59184# a_36350_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11934 a_77002_40202# a_77098_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11935 VDD a_10515_63143# a_14655_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11936 a_4032_49159# a_4240_48981# a_4174_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11937 VSS a_12895_13967# a_41766_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11938 a_19374_69222# a_16746_69224# a_19282_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11939 a_6531_38377# a_5631_38127# a_6459_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1194 a_17554_30663# a_17358_31069# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X11940 a_4960_40847# a_4259_40847# a_4792_41167# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u M=2
X11941 a_27710_72234# VDD a_27314_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11942 a_20378_64202# a_16746_64204# a_20286_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11943 a_18278_24918# VSS a_18370_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11944 a_22386_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11945 a_15397_39631# a_15131_39997# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11946 a_3801_13647# a_1929_10651# a_3677_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X11947 VSS a_4893_33821# a_4999_33781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X11948 a_30816_41605# a_29943_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11949 vcm_commonmode VSS a_37446_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1195 a_14679_31288# a_10506_29967# a_14949_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=1e+12p pd=6e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X11950 a_34763_47349# a_34906_47491# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11951 a_7755_70223# a_7289_70767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X11952 a_42770_14878# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11953 a_5087_23145# a_5211_24759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11954 a_12579_35862# a_12621_36091# a_12579_36189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11955 a_25702_24918# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11956 a_33830_72556# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11957 a_31726_17890# a_12899_11471# a_31330_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11958 a_11877_50645# a_11711_50645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X11959 a_4081_37289# a_1689_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1196 a_5695_74031# a_5345_74031# a_5600_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X11960 a_39758_58178# a_12901_58799# a_39362_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11961 VDD a_12985_19087# a_36350_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11962 VDD a_12981_59343# a_33338_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11963 a_46882_71552# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11964 a_17554_30663# a_14926_31849# a_18061_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X11965 a_6818_50959# a_5135_50069# a_6559_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X11966 VSS a_12727_58255# a_18674_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11967 VDD a_22063_47594# a_19788_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X11968 VSS a_11067_67279# a_18674_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11969 VDD a_9751_25071# a_11413_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1197 a_4985_31849# a_4702_32143# a_4903_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11970 VSS a_35463_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X11971 a_32795_41855# a_32029_41829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X11972 VDD a_2292_17179# a_8076_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11973 a_8029_11587# a_3327_9308# a_7938_11587# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X11974 a_24302_9858# a_12546_22351# a_24794_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X11975 a_2781_36873# a_1591_36501# a_2672_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X11976 VDD a_5599_74549# a_5475_74895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X11977 a_29322_71230# a_16362_71230# a_29414_71230# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X11978 VDD a_12231_60949# a_12218_61341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11979 a_1586_18695# a_10883_18007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1198 a_38754_56170# a_12257_56623# a_38358_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X11980 a_2163_63293# a_1586_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11981 a_10382_58487# a_10478_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11982 a_28714_15882# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11983 VSS a_6098_73095# a_7725_72765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11984 a_18731_38825# a_17799_38591# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11985 VSS a_8080_47607# a_6727_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11986 VSS a_2411_19605# a_2369_23805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X11987 VSS a_12727_15529# a_32730_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11988 VDD a_12947_71576# a_23298_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11989 VSS a_7210_55081# a_9278_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1199 a_40383_29575# a_12447_29199# a_40557_29451# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11990 VDD a_27797_29423# a_28089_31157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11991 VDD a_12355_15055# a_19282_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X11992 a_12161_31849# a_11143_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u
X11993 a_28423_52245# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X11994 a_9218_25321# a_9260_25045# a_9218_25071# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X11995 a_23390_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11996 a_47790_69222# a_12516_7093# a_47394_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X11997 VSS a_10975_66407# a_44778_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11998 a_33430_21540# a_16746_21538# a_33338_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X11999 vcm_commonmode a_16362_60186# a_32426_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_76346_38962# a_76180_38962# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X120 a_5546_12675# a_1929_12131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X1200 VDD config_2_in[8] a_1591_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12000 vcm_commonmode a_16362_19532# a_32426_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12001 a_42866_23516# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12002 a_42466_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12003 a_4458_45315# a_2927_39733# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12004 VDD a_3016_60949# a_4357_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12005 a_5315_68413# a_5167_68060# a_4952_68279# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12006 a_5964_35015# a_5691_36727# a_6106_35190# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X12007 VDD a_10145_60405# a_10035_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12008 a_46482_20536# a_16746_20534# a_46390_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12009 VDD a_12901_66665# a_27314_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1201 a_31822_56492# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12010 a_17274_11866# a_16362_11500# a_17366_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12011 a_45478_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12012 VSS a_22132_40865# a_22411_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12013 VDD a_12899_10927# a_35346_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12014 a_5087_29423# a_2011_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X12015 a_27421_42923# a_27271_37455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12016 a_21686_66210# a_12983_63151# a_21290_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12017 a_9782_71311# a_9024_71427# a_9219_71285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12018 VSS a_12355_65103# a_48794_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12019 VDD a_4298_58951# a_7019_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X1202 a_2847_12863# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12020 VDD a_12899_11471# a_48398_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12021 a_36442_12504# a_16746_12502# a_36350_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12022 a_7221_43541# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12023 a_45878_14480# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12024 a_43378_15882# a_16362_15516# a_43470_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12025 a_46482_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12026 VDD a_11943_63125# a_11851_64391# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12027 VDD a_12757_9295# a_12815_7663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12028 a_19374_22544# a_16746_22542# a_19282_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12029 a_34016_31849# a_33798_31145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1203 a_2899_28111# a_2473_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X12030 a_12727_58255# a_10055_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X12031 VSS a_12257_56623# a_38754_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12032 a_76648_39738# a_76744_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12033 a_42770_55166# VSS a_42374_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12034 a_18674_64202# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12035 a_8183_17289# a_7737_16917# a_8087_17289# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12036 VSS a_30762_49641# a_30557_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12037 a_20925_40743# a_21233_40956# a_19245_39747# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X12038 a_25702_65206# a_10975_66407# a_25306_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12039 VDD a_3484_61493# a_2944_63400# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1204 a_49798_72234# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X12040 a_49894_13476# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12041 a_46390_10862# a_12985_16367# a_46882_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12042 a_28817_52105# a_27627_51733# a_28708_52105# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X12043 a_20378_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12044 VDD a_12901_66959# a_43378_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12045 a_23298_63198# a_16362_63198# a_23390_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12046 a_35438_18528# a_16746_18526# a_35346_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12047 a_23845_29245# a_23195_29967# a_23739_29245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.596e+11p ps=1.6e+06u w=420000u l=150000u
X12048 VSS a_25321_29673# a_26112_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12049 VDD a_12901_58799# a_39362_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1205 vcm_commonmode a_16362_67214# a_45478_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12050 a_17643_48829# a_7050_53333# a_17280_48695# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12051 vcm_commonmode a_16362_68218# a_22386_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12052 a_39758_11866# a_12985_16367# a_39362_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12053 a_28714_56170# a_12257_56623# a_28318_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12054 a_24331_38591# a_23565_38565# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X12055 VDD a_12877_16911# a_26310_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12056 a_30912_39429# a_29943_39141# a_30816_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12057 VSS a_30035_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12058 VSS VDD a_37750_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12059 VDD a_12727_67753# a_47394_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1206 VDD a_12877_16911# a_36350_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12060 a_44874_64524# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12061 a_41370_61190# a_12981_59343# a_41862_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12062 a_5599_74549# a_6435_74005# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12063 vcm_commonmode a_16362_14512# a_36442_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12064 vcm_commonmode a_16362_59182# a_25398_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12065 a_29322_7850# VDD a_29814_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12066 a_30722_18894# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12067 a_23172_31573# a_23626_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X12068 a_34834_56492# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12069 VDD a_4578_40455# a_4529_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1207 a_8071_13255# a_1929_10651# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12070 a_18674_9858# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12071 a_5905_57961# a_4891_47388# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12072 a_9217_26703# a_4495_35925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X12073 a_47790_22910# a_11067_21583# a_47394_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12074 a_6927_39215# a_6473_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12075 VDD a_2840_66103# a_35069_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12076 a_17766_66532# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12077 a_30561_50959# a_26397_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12078 a_1761_27791# a_1591_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12079 a_2926_52637# a_1849_52271# a_2764_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1208 VDD a_10515_23975# a_19282_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12080 VDD a_12355_65103# a_21290_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12081 a_31753_47919# a_31186_48169# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12082 a_45386_60186# a_12727_58255# a_45878_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12083 a_9031_54135# a_9240_53877# a_9198_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X12084 VSS a_11179_9981# a_11140_10107# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12085 VDD a_14831_50095# a_30479_48576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X12086 VSS a_12659_54965# a_12987_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12087 a_17274_56170# a_16362_56170# a_17366_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12088 a_3935_56445# a_3005_56079# a_3572_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12089 VDD a_3307_18259# a_2411_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X1209 VDD a_10055_58791# a_49402_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12090 vcm_commonmode a_16362_58178# a_29414_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12091 a_40132_27247# a_29175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12092 a_5239_48767# a_5064_48841# a_5418_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12093 a_38850_55488# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12094 VSS a_28717_42917# a_29119_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12095 a_4429_14191# a_4075_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12096 a_22294_72234# VDD a_22786_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12097 VSS a_27652_38237# a_26753_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X12098 a_33734_70226# a_12901_66665# a_33338_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12099 VDD VDD a_40366_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X121 a_37446_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1210 a_4758_45369# a_5239_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X12100 a_12599_37782# a_12417_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12101 a_18278_62194# a_12355_15055# a_18770_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12102 a_7221_43541# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12103 a_22786_60508# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12104 a_30418_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12105 vcm_commonmode a_16362_17524# a_34434_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12106 a_4440_32259# a_2011_34837# a_4345_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=0p ps=0u w=420000u l=150000u
X12107 a_2553_47741# a_2509_47349# a_2387_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12108 VSS a_3301_26703# a_7755_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12109 a_3413_10389# a_3247_10389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1211 a_47486_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12110 VSS a_12985_16367# a_38754_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12111 a_13461_48579# a_5039_42167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12112 a_24849_51183# a_24683_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12113 a_3905_60797# a_3870_60563# a_3667_60405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12114 a_33727_42089# a_32795_41855# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12115 a_36746_61190# a_12355_15055# a_36350_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12116 a_22690_7850# VDD a_22294_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12117 a_2216_16885# a_2040_17289# a_2360_17277# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12118 VSS a_5671_21495# a_5547_21379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12119 a_13557_37999# a_13291_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1212 vcm_commonmode a_16362_59182# a_35438_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12120 a_75445_40202# a_75541_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12121 vcm_commonmode VSS a_43470_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12122 a_19678_71230# a_12947_71576# a_19282_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12123 a_3611_25731# a_3578_25625# a_3529_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12124 a_20682_67214# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12125 a_39454_7484# VDD a_39362_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12126 VDD a_12381_35836# a_12793_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12127 a_16746_13506# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X12128 VSS a_29391_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12129 a_6095_54697# a_6236_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1213 VSS a_12546_22351# a_48794_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12130 a_47394_18894# a_12895_13967# a_47886_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12131 VSS VSS a_47790_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12132 a_33734_66210# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12133 vcm_commonmode a_16362_21540# a_22386_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12134 a_31330_23914# a_12947_23413# a_31822_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12135 a_31330_19898# a_16362_19532# a_31422_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12136 VDD a_2672_26159# a_2847_26133# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12137 a_38450_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12138 a_17394_32275# a_17672_32259# a_17628_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12139 VSS a_12899_11471# a_37750_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1214 VSS a_12355_15055# a_43774_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12140 a_34267_31599# a_34016_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12141 a_20378_72234# VDD a_20286_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12142 a_41766_14878# a_12727_15529# a_41370_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12143 a_5600_10927# a_5483_11140# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12144 a_35438_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12145 a_8575_74853# a_10147_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X12146 VDD a_5024_67885# a_9775_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12147 a_2244_18231# config_1_in[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12148 a_5915_30511# a_6039_30663# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12149 a_30722_59182# a_12727_58255# a_30326_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1215 a_40762_18894# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12150 a_21290_15882# a_12727_13353# a_21782_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12151 a_24794_18496# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12152 a_24698_24918# VSS a_24302_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12153 VSS a_32227_48169# a_33669_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12154 VDD a_9484_11989# a_10259_10703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12155 a_42374_69222# a_12901_66959# a_42866_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12156 a_28410_15516# a_16746_15514# a_28318_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12157 vcm_commonmode a_16362_12504# a_25398_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12158 vcm_commonmode a_16362_63198# a_37446_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12159 a_2125_68053# a_1959_68053# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1216 vcm_commonmode a_16362_69222# a_18370_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12160 a_24394_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12161 a_38358_59182# a_12901_58799# a_38850_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12162 VSS a_34699_38771# a_34639_38825# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12163 a_2163_59585# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12164 a_27710_57174# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12165 VSS VSS a_31726_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12166 a_6096_28335# a_6066_28309# a_5906_28585# VSS sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=2.86e+11p ps=2.18e+06u w=650000u l=150000u
X12167 a_15259_46805# a_7000_43541# a_15457_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X12168 a_17869_28585# a_13390_29575# a_17869_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12169 a_43470_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1217 VSS VDD a_26706_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12170 vcm_commonmode a_16362_11500# a_29414_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12171 a_39454_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12172 a_28810_19500# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12173 a_5337_24643# a_4333_22895# a_5265_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12174 a_32826_68540# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12175 VDD a_11053_69135# a_11803_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X12176 a_27406_62194# a_16746_62196# a_27314_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12177 a_11482_16733# a_10405_16367# a_11320_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12178 VDD a_26495_38517# a_26319_38517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X12179 VSS a_75475_40594# a_76180_40594# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1218 a_22386_67214# a_16746_67216# a_22294_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12180 a_20286_65206# a_12355_65103# a_20778_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12181 a_41766_71230# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12182 a_40458_69222# a_16746_69224# a_40366_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12183 VSS a_30565_30199# a_17712_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12184 VDD a_3215_68351# a_3202_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12185 a_2847_45503# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12186 a_33338_64202# a_11067_13095# a_33830_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12187 a_25198_47741# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12188 VDD a_33155_40191# a_33015_40513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12189 VDD a_1923_54591# a_5592_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1219 VSS a_12677_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12190 VDD a_33839_28309# a_35616_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X12191 a_14369_27497# a_9529_28335# a_14287_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.15e+11p pd=2.83e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12192 VSS config_2_in[15] a_1591_52815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12193 a_18370_64202# a_16746_64204# a_18278_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12194 VSS a_9529_28335# a_22577_29111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12195 VDD a_26345_40871# a_19919_38695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X12196 VDD a_4951_44330# a_4839_43780# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12197 a_20682_20902# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12198 VSS a_12947_23413# a_23694_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12199 a_45478_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X122 a_11304_18543# a_10961_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X1220 VDD a_19596_34215# a_19500_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X12200 VDD a_8453_64757# a_5595_63125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12201 a_23298_56170# a_12947_56817# a_23790_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12202 VSS a_14471_28585# a_16101_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12203 a_6263_15645# a_5639_15279# a_6155_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12204 VDD a_10515_22671# a_30326_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12205 VSS a_12447_29199# a_29416_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12206 a_15788_28335# a_15315_27791# a_15697_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12207 a_45782_70226# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12208 a_28357_52271# a_27167_52271# a_28248_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X12209 a_44474_68218# a_16746_68220# a_44382_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1221 a_30722_70226# a_12901_66665# a_30326_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12210 vcm_commonmode a_16362_65206# a_41462_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12211 a_7175_53135# a_2840_53511# a_6985_52815# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X12212 a_43378_23914# a_16362_23548# a_43470_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12213 a_8367_74953# a_7921_74581# a_8271_74953# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X12214 a_1757_51183# a_1591_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12215 a_35742_62194# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12216 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12217 a_19697_29423# a_18829_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X12218 a_30722_12870# a_10055_58791# a_30326_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12219 a_42770_63198# a_15439_49525# a_42374_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1222 a_5363_30503# a_20881_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12220 a_18674_72234# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12221 a_27314_55166# VSS a_27806_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12222 VSS a_25263_29981# a_26020_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12223 VSS a_1761_35407# a_32143_35281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12224 VSS a_10717_17209# a_10651_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12225 a_5803_48285# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X12226 VDD a_3123_53047# a_2559_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X12227 VSS a_12516_7093# a_22690_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12228 a_48794_61190# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12229 a_47486_59182# a_16746_59184# a_47394_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1223 VDD a_76365_39738# a_76178_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12230 a_42374_9858# a_16362_9492# a_42466_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12231 a_4968_60405# a_5421_60137# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12232 a_20378_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12233 VDD a_39836_38567# a_39449_39868# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X12234 a_31725_31627# a_31659_31751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12235 a_36842_24520# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12236 VDD a_10680_54171# a_8199_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X12237 VDD a_11067_21583# a_40366_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12238 VDD a_12983_63151# a_39362_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12239 a_43085_30761# a_33641_29967# a_43003_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1224 a_4259_40847# a_4314_40821# a_4259_41167# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X12240 a_15775_40229# a_15009_40193# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X12241 a_27710_10862# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12242 a_23592_52271# a_4891_47388# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=0p ps=0u w=650000u l=150000u M=2
X12243 a_21663_41855# a_20715_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X12244 VDD a_19333_48463# a_19991_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12245 VSS a_7078_36103# a_7019_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.6975e+11p ps=2.13e+06u w=650000u l=150000u
X12246 a_40133_48463# a_18703_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12247 VDD a_11433_69921# a_11323_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12248 a_39454_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12249 a_7171_49929# a_6725_49557# a_7075_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1225 a_21290_22910# a_16362_22544# a_21382_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12250 VDD a_5320_18231# a_5271_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12251 VSS a_12981_59343# a_25702_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12252 a_28410_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12253 VDD a_1586_66567# a_1591_66415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12254 VSS a_2419_55687# a_2419_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12255 a_41351_39141# a_40403_37683# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X12256 a_11495_71855# a_11049_71855# a_11399_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12257 a_3484_61493# a_2959_47113# a_3704_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12258 a_37354_20902# a_12985_7663# a_37846_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12259 a_44874_72556# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1226 a_8132_53511# a_15285_52245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X12260 a_37354_16886# a_16362_16520# a_37446_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12261 a_33741_32463# a_19807_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12262 a_41462_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12263 VDD a_12981_59343# a_44382_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12264 a_31096_38341# a_30127_38053# a_31000_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12265 a_44382_62194# a_16362_62194# a_44474_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12266 VDD a_1761_52815# a_12191_37999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12267 VDD a_19478_51959# a_19435_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12268 a_2787_30503# a_13390_29575# a_14061_29199# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X12269 a_27314_72234# VSS a_27406_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1227 VDD a_2744_53511# a_2007_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12270 VSS a_12727_58255# a_29718_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12271 a_3876_61519# a_2787_62063# a_3621_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X12272 VSS a_11067_67279# a_29718_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12273 a_25398_55166# VDD a_25306_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12274 a_26706_16886# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12275 a_8566_39215# a_8127_39465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X12276 a_11339_24233# a_7571_29199# a_11121_23957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12277 a_31422_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12278 a_10257_56377# a_5682_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12279 a_16707_42359# a_15775_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1228 VDD a_15439_49525# a_44382_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12280 a_42718_27497# a_41334_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12281 VSS a_12877_14441# a_30722_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12282 a_40458_22544# a_16746_22542# a_40366_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12283 a_15599_28585# a_14273_27791# a_15793_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12284 VDD a_10515_23975# a_17274_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12285 a_39740_38567# a_38867_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12286 VDD VDD a_21290_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12287 VDD a_10055_58791# a_47394_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12288 VSS a_30091_35253# a_29177_34753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12289 a_5800_71855# a_4719_71855# a_5453_72097# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1229 vcm_commonmode a_16362_58178# a_39454_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12290 a_17274_64202# a_16362_64202# a_17366_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12291 a_38754_69222# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12292 a_35382_51157# a_35061_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12293 VSS a_13357_32143# a_26985_31605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12294 VDD a_18844_43439# a_18950_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12295 a_2215_18909# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12296 a_21382_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12297 VSS a_12983_63151# a_42770_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12298 a_2589_55535# a_2419_55535# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12299 a_20734_47158# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X123 a_10391_49855# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1230 a_20682_62194# a_12981_62313# a_20286_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12300 VDD a_2417_52513# a_2307_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12301 VSS a_31659_31751# a_37557_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12302 VSS a_28881_52271# a_37520_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12303 a_77664_39480# a_75475_40594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12304 a_38754_9858# a_12985_19087# a_38358_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12305 a_44474_21540# a_16746_21538# a_44382_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12306 a_18278_70226# a_12516_7093# a_18770_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12307 a_3149_68425# a_1959_68053# a_3040_68425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12308 a_18370_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12309 a_76346_40594# a_76180_40594# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X1231 VSS a_1586_9991# a_1591_16917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12310 a_32334_21906# a_16362_21540# a_32426_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12311 VDD a_15439_49525# a_42374_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12312 a_28318_11866# a_16362_11500# a_28410_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12313 a_34434_13508# a_16746_13506# a_34342_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12314 VDD a_12899_10927# a_46390_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12315 a_17366_23548# a_16746_23546# a_17274_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12316 VSS a_5547_31599# a_5915_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12317 VSS a_19780_38341# a_19743_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12318 VDD a_1586_36727# a_1591_36501# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12319 a_7464_39215# a_6927_39215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X1232 a_20713_40193# a_21387_39679# a_22260_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12320 a_47486_12504# a_16746_12502# a_47394_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12321 VSS a_23192_27791# a_27745_27275# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12322 a_35615_30199# a_35815_31751# a_35765_30287# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X12323 VSS a_24194_35823# a_24703_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12324 VSS a_10515_22671# a_36746_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12325 a_18661_28363# a_9529_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12326 a_29805_48829# a_17682_50095# a_29733_48829# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12327 VSS a_12727_67753# a_19678_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12328 a_16746_21538# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X12329 a_39362_61190# a_12981_59343# a_39854_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1233 VSS a_22062_31287# a_21273_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12330 a_47394_69222# a_16362_69222# a_47486_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12331 VSS a_12257_56623# a_49798_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12332 a_47394_7850# VSS a_47486_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12333 VDD a_23685_29111# a_24991_28129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12334 VDD a_12516_7093# a_41370_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12335 a_35838_8456# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12336 VDD a_2283_32362# a_1987_31812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12337 a_7289_70767# a_5877_70197# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X12338 a_41462_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12339 VSS a_13349_37973# a_13381_38365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1234 VSS a_3112_19319# a_3063_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12340 a_3859_10761# a_3413_10389# a_3763_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12341 a_24394_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12342 a_21290_66210# a_16362_66210# a_21382_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12343 a_26706_57174# a_10515_22671# a_26310_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12344 a_3663_39991# a_3759_39991# a_4061_40079# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12345 VSS a_7803_55509# a_8638_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12346 vcm_commonmode a_16362_68218# a_33430_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12347 VSS a_5043_19306# a_4379_18756# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12348 a_28816_28335# a_23192_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12349 a_13015_43493# a_12249_43457# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X1235 VSS a_12899_10927# a_30722_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12350 a_3137_28111# a_2315_24540# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12351 a_38358_67214# a_12983_63151# a_38850_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12352 VSS a_12985_19087# a_17670_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12353 a_33338_8854# a_12985_19087# a_33830_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12354 a_9011_74879# a_8836_74953# a_9190_74941# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12355 a_42866_65528# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12356 VDD a_4443_46607# a_5607_44343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12357 VSS a_20267_30503# a_42985_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12358 VSS a_9735_63669# a_9860_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12359 a_42374_55166# VSS a_42466_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1236 VSS a_2411_26133# a_2461_33597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12360 a_12189_46805# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12361 VSS a_25019_47679# a_24953_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X12362 VSS a_12981_62313# a_31726_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12363 a_32730_24918# a_12899_3855# a_32334_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12364 a_41462_71230# a_16746_71232# a_41370_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12365 a_28410_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12366 VDD a_1915_51946# a_1867_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12367 a_38754_22910# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12368 a_45782_23914# a_10515_23975# a_45386_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12369 a_42374_14878# a_12877_14441# a_42866_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1237 a_2840_66103# a_34895_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12370 VSS a_12985_7663# a_42770_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12371 VDD a_19675_49525# a_14985_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12372 a_6365_62063# a_2840_53511# a_5497_63303# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12373 a_4157_14191# a_3019_13621# a_4075_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12374 VDD a_4685_37583# a_6531_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12375 VDD a_1586_69367# a_1959_68053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12376 a_1887_12342# a_1929_12131# a_1887_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12377 a_1863_42729# a_2004_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12378 a_45878_56492# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12379 VDD a_2163_59585# a_2124_59459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1238 a_8652_17289# a_7737_16917# a_8305_16885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X12380 a_25306_24918# VSS a_25798_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12381 a_37761_44759# a_37857_44501# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12382 a_12907_56399# a_39503_43957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12383 a_2215_10205# a_1591_9839# a_2107_9839# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X12384 a_35742_15882# a_12877_14441# a_35346_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12385 a_8491_27023# a_12815_4399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12386 a_12357_37999# a_12191_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12387 a_29913_43457# a_29483_42943# a_30356_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12388 a_28318_56170# a_16362_56170# a_28410_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12389 VDD a_12899_11471# a_22294_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1239 a_22843_29415# a_37527_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X12390 a_35228_47375# a_22015_28111# a_34763_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12391 VDD a_12947_8725# a_20286_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12392 a_49894_55488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12393 a_29322_23914# a_12947_23413# a_29814_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12394 a_2834_14735# a_1757_14741# a_2672_15113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12395 a_29322_19898# a_16362_19532# a_29414_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12396 a_33338_72234# VDD a_33830_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12397 a_44778_70226# a_12901_66665# a_44382_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12398 a_36842_58500# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12399 VDD a_6467_55527# a_7171_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X124 a_18770_66532# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1240 a_27793_51733# a_27627_51733# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12400 a_30326_14878# a_16362_14512# a_30418_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12401 a_18370_72234# VDD a_18278_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12402 VDD a_7519_59575# a_7794_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12403 VSS a_10055_58791# a_36746_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12404 a_48490_61190# a_16746_61192# a_48398_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12405 a_32121_40741# a_32795_39679# a_33727_39913# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12406 vcm_commonmode a_16362_17524# a_45478_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12407 a_19282_15882# a_12727_13353# a_19774_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12408 VSS a_11067_21583# a_19678_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12409 a_34738_62194# a_12981_62313# a_34342_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1241 VSS a_6816_19355# a_7757_21379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X12410 VSS a_12985_16367# a_49798_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12411 a_13053_30511# a_12340_29967# a_12950_30511# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X12412 a_39113_32204# a_37557_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12413 a_23790_13476# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12414 a_10103_11079# a_9484_11989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12415 a_20286_10862# a_12985_16367# a_20778_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12416 VDD VSS a_26310_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12417 a_19374_8488# a_16746_8486# a_19282_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12418 VSS a_3357_22649# a_3291_22717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12419 a_6453_71855# a_5975_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1242 a_39055_39913# a_39449_39868# a_13909_39747# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X12420 a_18045_39105# a_17799_38591# a_18731_38825# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12421 VDD a_6791_70455# a_6598_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X12422 a_38454_43983# a_38277_43983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12423 a_31726_67214# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12424 a_20655_41271# a_21049_41245# a_20715_41245# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X12425 VDD a_2672_19631# a_2847_19605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12426 a_22386_17524# a_16746_17522# a_22294_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12427 VDD a_2847_30271# a_2834_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12428 vcm_commonmode a_16362_16520# a_49494_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12429 a_2300_61879# a_1823_72381# a_2228_61879# VSS sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1243 a_45386_71230# a_12901_66665# a_45878_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12430 a_26706_10862# a_12546_22351# a_26310_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12431 vcm_commonmode a_16362_21540# a_33430_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12432 a_22757_28585# a_2235_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12433 a_21686_59182# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12434 a_49494_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12435 a_9413_26703# a_6773_27805# a_9289_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X12436 a_32887_40767# a_32121_40741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X12437 a_2215_45021# a_1591_44655# a_2107_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X12438 a_22015_51840# a_19478_51959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X12439 a_4461_53113# a_3668_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1244 a_20975_37455# a_20827_37737# a_20612_37607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12440 a_31822_63520# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12441 a_26402_16520# a_16746_16518# a_26310_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12442 vcm_commonmode a_16362_13508# a_23390_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12443 VDD a_11067_67279# a_36350_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12444 VDD a_12202_54599# a_12631_52928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X12445 a_39454_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12446 a_36350_61190# a_16362_61190# a_36442_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12447 a_10515_22671# a_15617_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X12448 vcm_commonmode a_16362_63198# a_48490_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12449 VSS a_10964_25615# a_14711_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X1245 a_40458_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12450 a_2882_73309# a_2124_73211# a_2319_73180# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12451 a_12513_26409# a_7571_26151# a_12441_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12452 a_37888_34191# a_37711_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12453 a_25702_58178# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12454 VSS a_8753_19319# a_8104_18517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12455 a_39758_71230# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12456 a_38450_69222# a_16746_69224# a_38358_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12457 vcm_commonmode a_16362_66210# a_35438_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12458 VSS a_33080_37149# a_32181_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X12459 a_2834_49551# a_1757_49557# a_2672_49929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1246 VSS a_20747_27765# a_20685_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.3585e+12p ps=1.328e+07u w=650000u l=150000u M=4
X12460 VSS a_11999_67477# a_11957_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12461 a_37354_24918# VSS a_37446_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12462 a_5600_74031# a_5483_74244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12463 a_41462_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12464 VSS a_26397_51183# a_33045_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12465 a_37446_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12466 VSS a_26661_34428# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12467 VDD a_12967_50943# a_12954_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12468 a_19028_35823# a_18851_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12469 a_17889_44007# a_18197_44220# a_17863_44211# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1247 VDD a_4528_26159# a_7473_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12470 VDD a_5190_59575# a_14008_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12471 a_30818_69544# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12472 VSS a_12981_59343# a_33734_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12473 a_25398_63198# a_16746_63200# a_25306_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12474 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12475 VSS a_3751_72373# a_3697_72719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12476 vcm_commonmode a_16362_65206# a_39454_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12477 a_30326_59182# a_16362_59182# a_30418_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12478 a_12624_63151# a_11067_63143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12479 a_35581_31599# a_11067_46823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1248 a_26319_42869# a_26495_42869# a_26447_42895# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X12480 a_44778_24918# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12481 a_32494_48463# a_28108_48463# a_32402_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X12482 VDD a_25300_38567# a_25204_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12483 VDD a_3981_10357# a_3871_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12484 VDD a_23631_50069# a_23535_50247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12485 a_5297_52271# a_4918_52637# a_5225_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12486 VSS a_23911_35823# a_24017_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12487 a_35765_30287# a_33641_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12488 a_17366_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12489 a_6069_30761# a_6243_30662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1249 a_17670_60186# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12490 a_31330_65206# a_12355_65103# a_31822_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12491 a_18278_9858# a_12546_22351# a_18770_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12492 a_33430_55166# VDD a_33338_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12493 a_34738_16886# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12494 VSS a_41289_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12495 a_21012_30761# a_20946_30669# a_20904_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12496 a_12663_35431# a_32187_36161# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12497 a_9353_72399# a_9075_72737# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X12498 a_16362_65206# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X12499 VSS a_6243_30662# a_7295_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X125 a_49894_7452# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1250 a_16362_58178# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X12500 a_12318_18543# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12501 a_47790_15882# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12502 VSS VSS a_21686_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12503 a_18370_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12504 vcm_commonmode a_16362_71230# a_30418_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12505 a_29414_64202# a_16746_64204# a_29322_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12506 a_21290_57174# a_12257_56623# a_21782_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12507 VSS a_6816_19355# a_8256_20969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12508 VSS a_17799_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12509 a_32795_38053# a_31096_38341# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X1251 a_45386_8854# a_12985_19087# a_45878_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12510 VDD a_12947_71576# a_42374_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12511 a_31726_20902# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12512 VDD a_12355_15055# a_38358_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12513 a_1644_63669# a_1823_63677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12514 a_39272_31573# a_8491_41383# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12515 VSS a_4339_64521# a_9652_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12516 a_1954_61677# a_4307_67477# a_4253_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12517 VDD a_13510_44759# a_13515_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12518 a_19374_56170# a_16746_56172# a_19282_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12519 VSS a_5254_67503# a_8060_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1252 a_17670_19898# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12520 a_20685_28335# a_15661_29199# a_20972_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X12521 VSS a_12727_13353# a_24698_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12522 a_27710_18894# a_12899_10927# a_27314_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12523 VDD a_2041_61519# a_2141_61635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12524 a_21686_12870# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12525 VSS a_3667_60405# a_1823_62589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12526 a_8903_42301# a_8273_42479# a_8540_42167# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12527 VDD a_19596_42919# a_19500_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12528 a_46786_62194# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12529 VDD a_26495_37429# a_26319_37429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1253 VDD a_12981_62313# a_48398_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12530 a_17475_51157# a_17300_51183# a_17654_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12531 VSS a_12473_41781# a_12417_42134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12532 a_16753_49007# a_16587_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12533 a_10680_52245# a_33360_51701# a_32972_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12534 VSS config_2_in[6] a_1591_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12535 a_12473_41781# a_30715_41835# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X12536 VDD a_1923_54591# a_4771_56597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12537 a_40762_66210# a_12983_63151# a_40366_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12538 vcm_commonmode a_16362_62194# a_24394_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12539 a_11053_62607# a_10575_62911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1254 a_2689_65103# a_1768_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12540 a_25306_58178# a_10515_22671# a_25798_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12541 VSS a_12877_14441# a_28714_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12542 a_25702_11866# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12543 a_3672_58371# a_3618_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12544 a_38450_22544# a_16746_22542# a_38358_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12545 a_7623_13621# a_7797_13885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=5.72e+06u as=0p ps=0u w=1e+06u l=150000u
X12546 a_47886_24520# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12547 a_12047_57685# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12548 a_37446_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12549 a_32920_34191# a_32743_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1255 VSS a_1923_54591# a_1881_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12550 a_38380_30287# a_15607_46805# a_38077_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X12551 a_37750_64202# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12552 a_3677_13647# a_2283_15797# a_3605_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12553 a_35346_21906# a_11067_21583# a_35838_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12554 VSS a_1923_59583# a_10097_62973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12555 a_35346_17890# a_16362_17524# a_35438_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12556 VDD a_12727_15529# a_41370_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12557 a_12713_41923# a_15683_40767# a_16556_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12558 a_4620_55541# a_4433_55581# a_4533_55799# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X12559 VDD VSS a_24302_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1256 a_2080_56989# a_1643_56597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X12560 a_42374_63198# a_16362_63198# a_42466_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12561 a_48398_20902# a_12985_7663# a_48890_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12562 a_48398_16886# a_16362_16520# a_48490_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12563 a_1915_51946# a_2007_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12564 a_43870_8456# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12565 a_17670_67214# a_12727_67753# a_17274_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12566 a_20592_46983# a_12869_2741# a_20734_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X12567 a_47790_56170# a_12257_56623# a_47394_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12568 a_22535_28879# a_13357_32143# a_22441_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X12569 a_12039_69367# a_11803_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1257 VDD a_36116_44765# a_36336_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X12570 a_38358_12870# a_12877_16911# a_38850_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12571 a_5695_10927# a_5179_10927# a_5600_10927# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X12572 VDD a_12877_16911# a_45386_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12573 a_42866_10464# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12574 a_22448_39429# a_21479_39141# a_22352_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12575 a_10023_60809# a_9577_60437# a_9927_60809# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12576 VDD a_10515_23975# a_28318_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12577 a_25798_20504# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12578 VSS a_17311_46833# a_17257_46859# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12579 VSS a_12727_67753# a_40762_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1258 a_37534_51701# a_35568_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X12580 a_25398_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12581 a_28318_64202# a_16362_64202# a_28410_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12582 a_5595_33205# a_15911_31784# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12583 a_31004_40743# a_30035_40767# a_30967_41001# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12584 a_32426_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12585 vcm_commonmode a_16362_59182# a_44474_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12586 a_12410_60975# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12587 vcm_commonmode VSS a_38450_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12588 vcm_commonmode a_16362_69222# a_27406_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12589 VDD a_12877_14441# a_18278_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1259 a_29414_57174# a_16746_57176# a_29322_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12590 a_22762_27791# a_21012_30761# a_22649_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X12591 a_31422_67214# a_16746_67216# a_31330_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12592 a_13837_39860# a_13867_38870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12593 a_19258_47375# a_18539_47617# a_18695_47349# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X12594 a_36842_66532# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12595 a_2417_31841# a_2199_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12596 VSS a_1929_12131# a_7493_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12597 a_2325_69109# a_2107_69513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X12598 a_30326_22910# a_16362_22544# a_30418_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12599 VDD a_12355_65103# a_40366_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X126 a_45782_7850# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1260 a_1586_66567# a_4075_63151# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12600 a_11245_74031# a_10055_74031# a_11136_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X12601 a_29414_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12602 a_26310_12870# a_16362_12504# a_26402_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12603 VDD a_1586_21959# a_1591_29973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12604 VSS a_15775_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12605 a_2325_36469# a_2107_36873# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X12606 a_22690_61190# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12607 a_21382_59182# a_16746_59184# a_21290_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12608 VSS a_35463_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12609 a_19282_66210# a_16362_66210# a_19374_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1261 a_39758_8854# a_12947_8725# a_39362_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12610 VSS a_19028_35823# a_19134_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12611 a_45478_13508# a_16746_13506# a_45386_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12612 a_25312_37455# a_24413_39087# a_25091_37782# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X12613 a_19774_11468# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12614 VDD VDD a_34342_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12615 VDD a_5428_63669# a_5366_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X12616 VDD a_30855_41809# a_30715_41835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12617 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12618 VSS a_9989_46831# a_12263_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12619 a_30530_51183# a_28968_50871# a_30720_51183# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X1262 VDD a_13484_39325# a_26353_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12620 a_37354_62194# a_12355_15055# a_37846_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12621 a_2417_33205# a_2199_33609# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X12622 a_13692_44527# a_13515_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12623 VSS a_10515_22671# a_47790_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12624 a_16707_41271# a_15775_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12625 a_41862_60508# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12626 a_27314_8854# a_16362_8488# a_27406_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12627 a_22294_7850# VDD a_22786_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12628 VDD a_8197_31599# a_15290_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12629 a_26447_37455# a_13097_37455# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1263 a_31726_13874# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12630 a_6769_14013# a_4429_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12631 VDD a_12907_27023# a_39396_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12632 vcm_commonmode VSS a_22386_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12633 a_16666_7850# VDD a_16270_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12634 a_32826_7452# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12635 a_12139_71829# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12636 VDD a_25019_47679# a_25006_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X12637 a_32507_50959# a_2959_47113# a_32370_50871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12638 a_7073_51433# a_5909_51433# a_7001_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X12639 VDD a_10975_66407# a_17274_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1264 a_4842_45467# a_3987_19623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X12640 a_8273_42479# a_7815_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12641 a_24698_58178# a_12901_58799# a_24302_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12642 a_38754_71230# a_12947_71576# a_38358_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12643 a_31822_71552# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12644 a_27806_61512# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12645 a_17670_20902# a_11067_67279# a_17274_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12646 VSS a_4685_37583# a_6653_36611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X12647 a_4491_49334# a_4240_48981# a_4032_49159# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X12648 a_10501_55535# a_10075_55862# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12649 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1265 a_7580_61751# a_5682_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X12650 VSS a_12139_18517# a_12073_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12651 a_36746_23914# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12652 VSS a_25269_27791# a_27250_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X12653 a_2319_73180# a_2124_73211# a_2629_72943# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X12654 a_43870_18496# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12655 a_43774_24918# VSS a_43378_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12656 a_40366_15882# a_12727_13353# a_40858_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12657 VSS a_11067_21583# a_40762_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12658 VSS a_7775_10625# a_7736_10499# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12659 a_37446_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1266 a_18770_22512# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12660 VSS a_12355_65103# a_12899_11471# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12661 a_5749_18297# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12662 a_18445_46805# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12663 vcm_commonmode a_16362_12504# a_44474_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12664 VSS a_2872_44111# a_27945_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12665 a_42188_37149# a_41351_39141# a_42283_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12666 a_40276_28335# a_38436_29941# a_40176_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X12667 VSS a_12412_32143# a_14298_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X12668 a_2401_41941# a_2235_41941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12669 vcm_commonmode a_16362_22544# a_27406_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1267 a_32426_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12670 a_33734_16886# a_12727_13353# a_33338_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12671 a_9125_24527# a_9263_24501# a_9209_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12672 a_31422_20536# a_16746_20534# a_31330_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12673 a_26310_57174# a_16362_57174# a_26402_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12674 a_30418_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12675 VSS a_2411_19605# a_11661_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12676 a_26219_31171# a_25263_29981# a_26147_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12677 a_46786_15882# a_12877_14441# a_46390_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12678 VDD a_12899_10927# a_20286_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12679 VDD a_7571_26151# a_11865_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1268 a_22786_71552# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12680 a_29718_67214# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12681 a_8289_26409# a_4571_26677# a_8205_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12682 a_12786_30761# a_12999_29423# a_13053_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u w=650000u l=150000u
X12683 VDD a_9063_71553# a_9024_71427# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12684 a_21382_12504# a_16746_12502# a_21290_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12685 a_33430_63198# a_16746_63200# a_33338_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12686 a_30818_14480# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12687 a_2473_40821# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12688 VSS a_10288_53047# a_9507_53877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12689 a_34834_59504# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1269 a_49402_70226# a_12516_7093# a_49894_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12690 a_15039_38909# a_14859_38909# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12691 a_31422_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12692 a_38076_31573# a_35815_31751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12693 vcm_commonmode VSS a_30418_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12694 a_46482_62194# a_16746_62196# a_46390_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12695 a_19678_59182# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12696 VDD a_25015_48437# a_24773_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12697 a_47886_58500# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12698 vcm_commonmode a_16362_18528# a_43470_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12699 a_39673_28111# a_37699_27221# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X127 VSS a_12901_58799# a_25702_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1270 VSS a_5497_63303# a_5445_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X12700 a_36579_38007# a_35647_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12701 a_19678_17890# a_12899_11471# a_19282_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12702 VSS a_12257_56623# a_23694_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12703 a_17274_16886# a_12899_11471# a_17766_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12704 a_3330_70223# a_2960_70565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12705 VSS a_4127_63669# a_2927_68565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12706 a_6066_28309# a_2317_28892# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X12707 VSS a_5631_38127# a_5504_37815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X12708 a_29414_72234# VDD a_29322_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12709 VSS a_10055_58791# a_47790_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1271 VDD a_11067_67279# a_22294_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12710 a_10075_55862# a_8132_53511# a_10075_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12711 a_2319_63388# a_2163_63293# a_2464_63517# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X12712 a_8215_31055# a_7460_31055# a_8297_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X12713 a_11491_65327# a_10975_65327# a_11396_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X12714 VSS a_5254_67503# a_7479_57175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12715 a_31330_10862# a_12985_16367# a_31822_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12716 VDD a_12985_19087# a_38358_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12717 a_2104_33597# a_1987_33402# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12718 a_7113_24233# a_7059_24135# a_6989_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X12719 VDD a_30375_51335# a_19576_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1272 a_25388_35077# a_12713_36483# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X12720 VDD a_3031_47679# a_2959_47113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X12721 VDD a_12901_58799# a_24302_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12722 a_20378_18528# a_16746_18526# a_20286_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12723 a_32856_48463# a_32319_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12724 VSS a_5465_14967# a_5052_14709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X12725 a_24698_11866# a_12985_16367# a_24302_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12726 VDD a_6619_47607# a_5963_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X12727 a_38067_47349# a_27535_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12728 a_9135_25321# a_9260_25045# a_9218_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12729 a_42374_56170# a_12947_56817# a_42866_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1273 a_27710_8854# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12730 a_28810_69544# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12731 a_25306_66210# a_10975_66407# a_25798_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12732 a_8827_29967# a_3339_32463# a_8733_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X12733 VDD a_5453_72097# a_5343_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12734 a_36746_64202# a_12355_65103# a_36350_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12735 a_6435_47893# a_6260_47919# a_6614_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12736 VSS a_12249_43457# a_12283_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X12737 a_6515_67477# a_2952_66139# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X12738 a_12165_55535# a_10975_55535# a_12056_55535# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X12739 a_8958_65961# a_10747_68565# a_10705_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1274 a_29913_43457# a_29483_42943# a_30415_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X12740 VDD a_12985_7663# a_34342_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12741 a_18811_36965# a_15305_38543# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X12742 vcm_commonmode a_16362_14512# a_21382_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12743 VSS a_4461_48981# a_4395_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12744 a_35061_51727# a_34895_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12745 VSS a_12970_34191# a_13515_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12746 a_37446_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12747 a_36350_9858# a_16362_9492# a_36442_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12748 a_37750_72234# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12749 a_14293_37455# a_13867_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1275 a_38327_44759# a_34222_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12750 VSS a_12516_7093# a_41766_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12751 VSS a_12231_60949# a_12165_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12752 a_29322_65206# a_12355_65103# a_29814_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12753 a_9497_10383# a_9219_11471# a_9414_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12754 VSS a_17682_50095# a_25317_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12755 a_30326_60186# a_12727_58255# a_30818_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12756 a_30967_41001# a_30035_40767# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12757 a_49494_69222# a_16746_69224# a_49402_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12758 vcm_commonmode a_16362_66210# a_46482_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12759 a_35438_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1276 VSS a_22995_30663# a_22151_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12760 VSS a_12381_35836# a_12800_36189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12761 a_5443_62063# a_4758_45369# a_5274_62313# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X12762 a_75475_38962# a_75199_38962# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12763 VSS a_4951_44330# a_4839_43780# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12764 a_9405_56623# a_3295_62083# a_9187_56597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X12765 VSS a_4762_35484# a_4941_35727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12766 a_19282_57174# a_12257_56623# a_19774_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12767 a_23790_55488# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12768 a_29718_20902# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12769 a_4499_45743# a_4149_45743# a_4404_45743# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1277 VDD a_19502_51157# a_6559_59879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12770 VSS a_12981_59343# a_44778_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12771 VSS a_10275_21495# a_9263_24501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X12772 a_40458_56170# a_16746_56172# a_40366_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12773 a_41766_17890# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12774 a_7803_11703# a_8167_11561# a_8102_11587# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X12775 VSS a_12901_66665# a_27710_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12776 a_10995_14333# a_1586_18695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12777 a_6733_69135# a_5924_69135# a_4307_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12778 VDD a_12899_3855# a_32334_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12779 a_4057_13647# a_3677_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X1278 VSS a_27247_43047# a_24893_37429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12780 a_19678_12870# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12781 a_25398_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12782 VSS a_12985_16367# a_23694_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12783 a_12473_42869# a_32187_40513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X12784 VSS a_6271_72943# a_6927_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12785 VDD a_1916_33927# a_1867_32839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12786 VDD a_26397_51183# a_32311_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12787 a_24937_39306# a_1761_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12788 a_21686_61190# a_12355_15055# a_21290_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12789 VSS a_12727_58255# a_48794_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1279 a_22294_61190# a_16362_61190# a_22386_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12790 a_44474_55166# VDD a_44382_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12791 a_45782_16886# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12792 VSS a_11067_67279# a_48794_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12793 VDD a_2376_23047# a_2007_21237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12794 VDD a_18539_47617# a_18500_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12795 a_27406_65206# a_16746_65208# a_27314_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12796 a_43378_10862# a_16362_10496# a_43470_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12797 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X12798 a_19203_39958# a_15189_39889# a_19131_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X12799 VSS a_4891_47388# a_27009_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X128 a_24987_36649# a_24055_36415# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X1280 a_8747_14735# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X12800 VDD a_3983_10927# a_1689_10396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X12801 a_33830_20504# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12802 VDD VDD a_40366_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12803 a_33430_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12804 a_32334_18894# a_12895_13967# a_32826_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12805 VSS a_12899_3855# a_32730_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12806 a_29414_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12807 a_26310_20902# a_16362_20536# a_26402_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12808 VSS a_34297_35516# a_33989_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12809 VDD a_12981_62313# a_36350_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1281 VSS a_12901_66959# a_46786_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12810 a_16746_16518# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X12811 a_21382_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12812 a_7829_74281# a_6224_73095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12813 VSS VDD a_39758_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12814 a_11902_27247# a_8935_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X12815 a_17366_57174# a_16746_57176# a_17274_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12816 a_18674_18894# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12817 VDD a_12355_15055# a_49402_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12818 a_23390_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12819 a_1644_65845# a_1823_65853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1282 a_43774_66210# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12820 a_25702_60186# a_12981_59343# a_25306_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12821 a_25702_19898# a_12895_13967# a_25306_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12822 VSS a_12899_11471# a_22690_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12823 a_11756_12381# a_11542_12381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12824 a_20378_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12825 VSS a_5039_42167# a_4989_42255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12826 VDD a_3452_70537# a_3510_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12827 a_1761_2767# a_1591_2767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12828 a_49798_7850# VDD a_49402_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12829 a_37354_70226# a_12516_7093# a_37846_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1283 a_2143_15271# a_5147_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X12830 a_18947_51017# a_18501_50645# a_18851_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12831 a_19446_51183# a_4758_45369# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X12832 a_34342_12870# a_16362_12504# a_34434_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12833 a_4499_45743# a_3983_45743# a_4404_45743# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X12834 a_17983_41855# a_16744_41605# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X12835 VSS a_12901_66959# a_34738_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12836 VSS a_2289_35113# a_3342_34639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12837 a_2672_36873# a_1757_36501# a_2325_36469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12838 vcm_commonmode a_16362_63198# a_22386_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12839 a_47394_11866# a_16362_11500# a_47486_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1284 a_41370_23914# a_12947_23413# a_41862_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12840 a_23298_59182# a_12901_58799# a_23790_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12841 VDD a_11067_46823# a_14365_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12842 VSS a_35382_51157# a_34943_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12843 a_36520_36165# a_35647_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X12844 a_36442_23548# a_16746_23546# a_36350_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12845 a_35438_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12846 VSS a_2713_35925# a_2647_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12847 a_8005_53333# a_4339_64521# a_8258_53359# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X12848 a_2107_15113# a_1591_14741# a_2012_15101# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X12849 a_49494_22544# a_16746_22542# a_49402_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1285 a_41370_19898# a_16362_19532# a_41462_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12850 VSS a_12727_67753# a_38754_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12851 a_35742_65206# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12852 VDD VDD a_42374_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12853 a_35838_17492# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12854 VSS a_30412_34337# a_29513_34428# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X12855 VSS a_41167_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12856 a_24394_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12857 a_9543_65327# a_5024_67885# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12858 a_48794_64202# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12859 a_46390_21906# a_11067_21583# a_46882_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1286 a_11067_63143# a_14634_47349# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X12860 VSS a_1586_18695# a_8123_14741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12861 a_46390_17890# a_16362_17524# a_46482_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12862 a_2399_47375# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12863 VDD a_12546_22351# a_17274_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12864 a_8228_38377# a_3949_41935# a_8129_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12865 a_32730_58178# a_12901_58799# a_32334_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12866 a_11599_55901# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12867 a_35438_70226# a_16746_70228# a_35346_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12868 VSS a_2686_70223# a_4345_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12869 a_15970_38870# a_12663_39783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1287 VSS a_1761_37039# a_31131_35281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12870 a_38754_56170# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12871 a_43470_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12872 a_40366_66210# a_16362_66210# a_40458_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12873 a_45782_57174# a_10515_22671# a_45386_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12874 a_39854_16488# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12875 a_36350_13874# a_12727_15529# a_36842_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12876 a_40858_11468# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12877 a_28714_67214# a_12727_67753# a_28318_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12878 a_7293_45173# a_7075_45577# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12879 VSS a_11067_13095# a_25702_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1288 a_32311_48169# a_31753_47919# a_32227_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.95e+11p pd=5.19e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12880 VDD a_37706_44135# a_37711_43983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12881 vcm_commonmode a_16362_9492# a_46482_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12882 a_26310_65206# a_16362_65206# a_26402_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12883 a_11054_59343# a_11019_59575# a_10751_59575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12884 a_30418_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12885 a_18674_59182# a_12727_58255# a_18278_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12886 VDD a_5271_17999# a_5363_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X12887 a_40366_7850# VSS a_40458_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12888 a_1849_31599# a_1683_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12889 a_13867_37782# a_13097_37455# a_13795_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X1289 VDD a_9305_53511# a_7764_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X12890 a_17798_32143# a_17672_32259# a_17394_32275# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X12891 a_28708_52105# a_27793_51733# a_28361_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X12892 a_30722_70226# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12893 a_2781_15529# a_2143_15271# a_1895_14906# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X12894 a_2847_38975# a_2672_39049# a_3026_39037# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12895 a_11602_25071# a_11163_25321# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X12896 a_34834_67536# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12897 VSS a_1923_73087# a_9913_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12898 VDD a_12877_14441# a_29322_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12899 a_17366_10496# a_16746_10494# a_17274_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X129 VDD a_12355_65103# a_22294_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1290 a_48490_23548# a_16746_23546# a_48398_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12900 a_19580_49159# a_19788_48981# a_19722_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X12901 a_8038_18870# a_6816_19355# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12902 a_44382_24918# VSS a_44874_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12903 a_13123_38231# a_32831_35307# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X12904 VSS a_2283_32362# a_1987_31812# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X12905 a_34342_57174# a_16362_57174# a_34434_57174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X12906 a_47886_66532# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12907 a_20682_62194# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12908 a_26402_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12909 a_4233_30761# a_2216_28309# a_4161_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1291 vcm_commonmode a_16362_20536# a_45478_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X12910 VDD a_15011_34717# a_15037_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X12911 a_17274_67214# a_16362_67214# a_17366_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12912 VSS VSS a_19678_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12913 a_47394_56170# a_16362_56170# a_47486_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12914 VSS a_7749_55535# a_8128_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X12915 VSS a_10515_23975# a_34738_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12916 a_33734_61190# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12917 a_32426_59182# a_16746_59184# a_32334_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12918 a_12591_31029# a_12935_31287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12919 VSS a_2467_53034# a_1987_52484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1292 a_39029_29673# a_33641_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X12920 a_12680_53511# a_4351_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X12921 a_2315_24540# a_2847_23743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X12922 VDD a_12257_56623# a_41370_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12923 a_14079_41046# a_12801_38517# a_13620_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12924 a_21782_24520# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12925 VSS a_18811_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X12926 VDD a_12983_63151# a_24302_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12927 a_48398_62194# a_12355_15055# a_48890_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12928 a_2672_36873# a_1591_36501# a_2325_36469# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X12929 VDD a_34391_48682# a_31768_55394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1293 a_26802_70548# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12930 a_22448_38341# a_21479_38053# a_22352_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X12931 a_24394_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12932 a_9443_23145# a_8933_22583# a_9223_22895# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X12933 a_25300_39655# a_24331_39679# a_25263_39913# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12934 a_1757_40303# a_1591_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12935 a_21051_47158# a_7571_29199# a_20592_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12936 a_6559_63401# a_4119_70741# a_6641_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X12937 VSS a_11067_21583# a_38754_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12938 a_32951_27247# a_30788_28487# a_32779_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X12939 vcm_commonmode VSS a_33430_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1294 a_47486_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12940 VSS a_30565_30199# a_42709_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12941 a_25484_37253# a_24515_36965# a_25447_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X12942 a_2952_46805# a_4123_37013# a_4081_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12943 a_31422_9492# a_16746_9490# a_31330_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12944 VDD VSS a_45386_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12945 a_36746_72234# VDD a_36350_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12946 a_22294_20902# a_12985_7663# a_22786_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12947 a_13097_37455# a_12671_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X12948 a_2464_59343# a_2250_59343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12949 a_22294_16886# a_16362_16520# a_22386_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1295 a_19282_14878# a_16362_14512# a_19374_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X12950 VDD a_12901_58799# a_32334_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12951 VSS a_4351_67279# a_8675_68047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X12952 VDD a_10975_66407# a_28318_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12953 a_25798_62516# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12954 VDD a_12587_51335# a_11855_51959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12955 a_49798_71230# a_12947_71576# a_49402_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12956 a_32730_11866# a_12985_16367# a_32334_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12957 VDD a_29887_32375# a_18151_52263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X12958 VSS a_4719_33239# a_4191_33449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X12959 a_14373_50095# a_6646_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X1296 VDD a_10472_26159# a_11522_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X12960 a_3697_35523# a_2011_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12961 a_75162_39738# a_75258_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X12962 VDD a_2840_66103# a_7933_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12963 a_2467_53034# a_2559_52789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X12964 a_28410_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12965 a_41462_17524# a_16746_17522# a_41370_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12966 VDD a_19780_41605# a_19684_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X12967 a_15970_38543# a_12663_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X12968 a_45782_10862# a_12546_22351# a_45386_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X12969 VDD a_10515_22671# a_18278_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1297 VSS a_4985_61021# a_5091_60981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X12970 a_8305_16885# a_8087_17289# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X12971 VDD a_4227_73791# a_4214_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12972 a_19591_50943# a_19416_51017# a_19770_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X12973 a_7637_53877# a_6559_59663# a_7794_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X12974 a_28810_14480# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12975 a_28714_20902# a_11067_67279# a_28318_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12976 a_32125_29673# a_32038_29575# a_25971_52263# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X12977 VDD a_8583_33551# a_32743_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12978 a_40762_59182# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12979 a_4220_68021# a_3693_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1298 a_40762_59182# a_12727_58255# a_40366_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12980 a_23694_69222# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12981 VDD a_1586_45431# a_3983_45743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12982 VSS config_1_in[4] a_1591_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X12983 a_10037_73487# a_8003_72917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12984 a_3026_12925# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12985 vcm_commonmode a_16362_13508# a_42466_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12986 a_1761_40847# a_1591_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X12987 a_18674_12870# a_10055_58791# a_18278_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12988 a_8581_18319# a_8539_18231# a_8111_18825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X12989 a_13867_37455# a_13613_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1299 VDD a_12947_8725# a_32334_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X12990 a_1757_18543# a_1591_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X12991 a_5803_48285# a_5179_47919# a_5695_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12992 a_41334_29575# a_41232_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X12993 a_27422_29789# a_5363_30503# a_26694_29473# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12994 vcm_commonmode a_16362_23548# a_25398_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12995 a_27195_32375# a_26985_31605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X12996 a_38358_71230# a_16362_71230# a_38450_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12997 a_29322_10862# a_12985_16367# a_29814_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X12998 a_44778_58178# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12999 a_11120_69679# a_8958_65961# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u M=1397
X130 a_3301_27791# a_2899_28111# a_3137_28111# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X1300 VDD a_3339_30503# a_15661_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.6e+11p ps=7.72e+06u w=1e+06u l=150000u
X13000 a_4287_65540# a_4167_64783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X13001 a_44778_16886# a_12727_13353# a_44382_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13002 a_8038_18543# a_6816_19355# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13003 a_27710_68218# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13004 a_44382_9858# a_16362_9492# a_44474_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13005 a_18370_18528# a_16746_18526# a_18278_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13006 VDD a_12899_10927# a_31330_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13007 a_9526_61751# a_9431_60214# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13008 VSS a_14076_35077# a_14039_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13009 a_32426_12504# a_16746_12502# a_32334_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1301 VDD a_5254_67503# a_7479_57175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13010 VSS a_4248_29967# a_8117_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13011 a_44474_63198# a_16746_63200# a_44382_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13012 vcm_commonmode a_16362_60186# a_41462_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13013 vcm_commonmode a_16362_19532# a_41462_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13014 a_45878_59504# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13015 a_8041_15279# a_7987_15431# a_7959_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13016 VSS a_10515_22671# a_21686_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13017 a_2319_56860# a_2163_56765# a_2464_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X13018 VSS a_5239_48767# a_4891_47388# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X13019 a_11771_23671# a_7841_22895# a_11945_23777# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1302 a_34834_18496# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13020 a_24302_61190# a_12981_59343# a_24794_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13021 a_33430_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13022 VDD a_29513_34428# a_29119_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13023 a_32334_69222# a_16362_69222# a_32426_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13024 vcm_commonmode a_16362_14512# a_19374_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13025 VDD a_12901_66665# a_36350_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13026 a_28318_16886# a_12899_11471# a_28810_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13027 a_7100_72105# a_6913_72399# a_7009_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13028 a_10767_20495# a_8933_22583# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X13029 a_9290_54991# a_6515_62037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1303 a_34738_24918# a_12899_3311# a_34342_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13030 a_20433_29967# a_7862_34025# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13031 a_36442_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13032 a_19374_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13033 VSS a_9513_65301# a_10317_67191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13034 VDD a_17039_51157# a_19675_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13035 a_15812_31029# a_16101_31029# a_16035_31375# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X13036 a_34342_20902# a_16362_20536# a_34434_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13037 a_39176_44527# a_38999_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13038 a_48490_64202# a_16746_64204# a_48398_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13039 a_40366_57174# a_12257_56623# a_40858_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1304 a_23390_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13040 a_10935_11989# a_11138_12267# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13041 VDD a_4812_13879# a_5169_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13042 a_23298_67214# a_12983_63151# a_23790_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13043 VDD a_2928_67191# a_2559_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13044 a_34738_65206# a_10975_66407# a_34342_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13045 VDD a_32121_44545# a_33668_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X13046 a_22411_39095# a_21479_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X13047 a_12263_26409# a_7571_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X13048 a_1945_43023# a_1593_42479# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13049 a_38450_56170# a_16746_56172# a_38358_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1305 VSS a_24331_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13050 a_39758_17890# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13051 VDD a_19217_51701# a_12755_53030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13052 VSS a_12727_13353# a_43774_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13053 a_40762_12870# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13054 VSS a_9367_29397# a_12244_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13055 a_23694_22910# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13056 a_9289_26703# a_3607_34639# a_9217_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13057 a_30722_23914# a_10515_23975# a_30326_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13058 a_5707_59887# a_5653_60039# a_5611_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13059 a_30818_56492# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1306 a_17497_29423# a_2235_30503# a_17415_29423# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13060 a_48794_72234# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13061 a_44382_58178# a_10515_22671# a_44874_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13062 a_20682_15882# a_12877_14441# a_20286_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13063 VSS a_22632_41831# a_22595_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13064 a_44778_11866# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13065 VSS a_8575_74853# a_10833_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13066 a_18105_32509# a_2099_59861# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13067 VSS a_32365_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13068 a_6607_39991# a_4314_40821# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13069 VSS a_2944_64488# a_2882_64605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X1307 a_23694_69222# a_12516_7093# a_23298_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13070 a_27710_21906# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13071 a_22259_48981# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13072 a_29483_42943# a_28717_42917# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X13073 a_28248_52271# a_27333_52271# a_27901_52513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13074 VSS a_12355_15055# a_42770_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13075 a_39454_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13076 VDD a_5913_11169# a_5803_11293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13077 a_21712_43781# a_20743_43493# a_21675_43447# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13078 VDD a_39244_41953# a_38345_42044# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X13079 VSS VDD a_25702_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1308 VSS a_10975_66407# a_20682_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13080 a_16746_57176# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X13081 a_26267_34473# a_26661_34428# a_13484_39325# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X13082 a_21782_58500# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13083 a_17670_13874# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13084 a_30764_7638# a_26523_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X13085 a_49402_7850# VSS a_49494_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13086 a_11298_74397# a_10221_74031# a_11136_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13087 VDD a_9260_25045# a_9209_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13088 VSS a_10055_58791# a_21686_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13089 a_18370_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1309 VSS a_20612_37607# a_13837_38772# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13090 vcm_commonmode a_16362_17524# a_30418_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13091 VDD VSS a_43378_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13092 a_37846_8456# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13093 vcm_commonmode a_16362_58178# a_38450_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13094 VSS a_11067_13095# a_33734_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13095 VDD a_34699_37683# a_34725_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13096 VDD a_11053_62607# a_11763_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13097 a_2376_23047# a_2317_28892# a_2518_23222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X13098 a_12981_62313# a_12712_62313# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13099 a_34342_65206# a_16362_65206# a_34434_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X131 a_26137_29423# a_26063_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1310 a_11251_59879# a_14365_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u M=2
X13100 a_8015_21807# a_7571_22057# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X13101 VDD a_10515_23975# a_47394_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13102 a_4595_48841# a_4149_48469# a_4499_48841# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X13103 a_44874_20504# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13104 a_44474_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13105 a_17889_36391# a_18197_36604# a_17863_36595# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X13106 a_1846_64491# a_2124_64507# a_2080_64605# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13107 VSS a_12985_19087# a_19678_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13108 VSS a_12981_62313# a_19678_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13109 a_14634_47349# a_11067_46823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1311 a_11521_66567# a_12047_57685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13110 a_4219_34551# a_2473_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X13111 a_47394_64202# a_16362_64202# a_47486_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13112 a_1586_66567# a_4075_63151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13113 a_12157_64015# a_11053_62607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13114 a_27183_36965# a_25300_38567# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X13115 a_10699_25731# a_9955_20969# a_10603_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13116 a_6713_37903# a_3305_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.7125e+11p pd=4.05e+06u as=0p ps=0u w=650000u l=150000u
X13117 a_30035_40767# a_29269_40741# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X13118 a_29718_8854# a_12947_8725# a_29322_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13119 a_35932_41953# a_35647_41317# a_36520_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1312 a_47790_65206# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13120 VDD a_12877_14441# a_37354_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13121 a_34834_12472# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13122 a_29863_39913# a_28931_39679# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X13123 VSS a_9083_13879# a_10339_14735# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13124 a_17766_22512# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13125 VSS a_2847_9813# a_2781_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X13126 VSS a_5363_30503# a_20821_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13127 a_3885_35523# a_3697_35523# a_3803_35523# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13128 VDD a_34062_47607# a_33868_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13129 a_10008_51549# a_9794_51549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1313 a_38450_15516# a_16746_15514# a_38358_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13130 a_48398_70226# a_12516_7093# a_48890_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13131 VDD a_11067_67279# a_21290_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13132 a_48490_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13133 a_45386_12870# a_16362_12504# a_45478_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13134 a_5331_18517# a_5156_18543# a_5510_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13135 a_24746_31849# a_24667_31055# a_25013_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.9825e+11p pd=1.91e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X13136 a_24394_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13137 a_21290_61190# a_16362_61190# a_21382_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13138 VSS a_12901_66959# a_45782_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13139 VDD a_14076_35077# a_13980_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1314 a_47886_17492# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13140 a_19596_42919# a_18627_42943# a_19559_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13141 vcm_commonmode a_16362_63198# a_33430_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13142 a_34434_24552# VDD a_34342_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13143 VSS a_2847_12863# a_2781_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X13144 VDD a_1586_69367# a_2971_73493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13145 a_24698_71230# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13146 a_23390_69222# a_16746_69224# a_23298_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13147 a_11713_66415# a_11659_66567# a_11617_66415# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X13148 vcm_commonmode a_16362_66210# a_20378_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13149 a_38850_11468# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1315 vcm_commonmode a_16362_12504# a_35438_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13150 VDD a_20359_29199# a_32509_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X13151 a_10562_62607# a_9485_62613# a_10400_62985# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13152 a_47486_23548# a_16746_23546# a_47394_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13153 a_22294_24918# VSS a_22386_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13154 VDD a_12983_63151# a_32334_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13155 VDD a_20612_37607# a_13837_38772# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13156 a_25798_70548# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13157 VSS a_1586_66567# a_1591_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13158 VSS a_5190_59575# a_5179_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X13159 a_18278_14878# a_16362_14512# a_18370_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1316 a_45386_18894# a_16362_18528# a_45478_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13160 VDD a_12947_8725# a_22294_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13161 a_16270_7850# VDD a_16762_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13162 a_41167_42943# a_37551_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X13163 a_29915_49007# a_14831_50095# a_29055_49525# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X13164 a_22386_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13165 VSS a_32029_41829# a_33543_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13166 a_15557_52245# a_15892_51843# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13167 a_28410_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13168 a_25306_60186# a_16362_60186# a_25398_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13169 a_7086_21263# a_3339_43023# a_7002_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 vcm_commonmode a_16362_22544# a_18370_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13170 VSS a_12727_67753# a_49798_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13171 a_46786_65206# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13172 vcm_commonmode a_16362_8488# a_35438_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13173 a_37446_15516# a_16746_15514# a_37354_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13174 VDD a_1591_72943# a_2083_74913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13175 a_12985_25615# a_12394_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13176 vcm_commonmode a_16362_65206# a_24394_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13177 VSS a_2319_59317# a_2250_59343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X13178 VSS a_35568_49525# a_36116_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13179 a_5877_54421# a_5531_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1318 a_15009_47919# a_14655_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13180 a_3594_15955# a_3911_16065# a_3869_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X13181 a_45478_8488# a_16746_8486# a_45386_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13182 a_36746_57174# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13183 a_33830_62516# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13184 a_11759_51959# a_5190_59575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13185 a_5023_72068# a_7100_72105# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X13186 VDD a_12546_22351# a_28318_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13187 a_2834_26525# a_1757_26159# a_2672_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13188 VDD a_13528_36055# a_12641_36596# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13189 a_43774_58178# a_12901_58799# a_43378_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1319 a_22386_20536# a_16746_20534# a_22294_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13190 VSS VSS a_40762_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13191 a_9670_24527# a_9043_24527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13192 VDD a_12999_29423# a_12786_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13193 a_28883_52031# a_28708_52105# a_29062_52093# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13194 a_26706_68218# a_12901_66959# a_26310_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13195 a_46882_61512# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13196 a_12671_43222# a_12713_43011# a_12671_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13197 vcm_commonmode a_16362_11500# a_38450_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13198 VSS a_8105_21263# a_7841_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13199 vcm_commonmode a_16362_56170# a_27406_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X132 a_12907_27023# a_40599_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X1320 a_37750_57174# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13200 a_37846_19500# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13201 a_5964_35015# a_4811_34855# a_6106_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13202 a_32730_15882# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13203 a_20286_8854# a_16362_8488# a_20378_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13204 a_6750_19126# a_3247_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X13205 a_4149_65327# a_3983_65327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13206 a_41441_28335# a_29175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13207 a_2369_9839# a_2325_10081# a_2203_9839# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13208 VDD a_16928_44007# a_16832_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13209 a_19774_63520# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1321 VSS a_7755_54999# a_7210_55081# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X13210 a_29718_59182# a_12727_58255# a_29322_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13211 VDD a_12355_15055# a_23298_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13212 a_25873_51183# a_24683_51183# a_25764_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13213 a_30418_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13214 VDD a_8575_74853# a_9364_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13215 a_32396_49007# a_14831_50095# a_32135_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X13216 a_16997_51183# a_16953_51425# a_16831_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X13217 a_7557_49007# a_7387_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X13218 a_45878_67536# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13219 a_38210_30199# a_12447_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1322 a_15775_42405# a_14919_43421# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X13220 VSS a_2419_48783# a_11753_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13221 a_32134_49159# a_27869_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X13222 a_2899_27023# a_2315_24540# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13223 VDD a_7067_30663# a_7019_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13224 VSS a_32823_29397# a_40276_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13225 a_15683_39141# a_13097_39631# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X13226 a_45386_57174# a_16362_57174# a_45478_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13227 a_1765_5059# a_1681_5175# a_1683_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13228 a_31726_62194# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13229 a_13669_35253# a_33015_36161# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X1323 VSS VSS a_41766_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13230 a_34337_29967# a_30788_28487# a_32038_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X13231 a_28318_67214# a_16362_67214# a_28410_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13232 VDD a_12981_59343# a_27314_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13233 a_17222_27247# a_16865_27511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X13234 VSS a_10515_23975# a_45782_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13235 VSS a_7203_10383# a_9219_11471# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X13236 a_32232_30511# a_31659_31751# a_31741_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13237 VDD a_41842_27221# a_43085_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13238 VSS a_75199_40594# a_75628_40594# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13239 a_23390_22544# a_16746_22542# a_23298_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1324 a_7862_34025# a_6662_34025# a_7526_33775# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X13240 a_18278_59182# a_16362_59182# a_18370_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13241 a_32826_24520# a_12899_3855# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13242 VSS a_8079_43732# a_6863_42692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13243 a_22386_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13244 a_38754_17890# a_12899_11471# a_38358_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13245 a_5959_13621# a_5755_14709# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13246 a_7436_46983# a_7644_46805# a_7578_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13247 VDD a_9613_48981# a_9643_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13248 a_48490_72234# VDD a_48398_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13249 a_22690_64202# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1325 VSS a_23830_49525# a_24638_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13250 a_36350_55166# VSS a_36842_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13251 a_4717_48437# a_4499_48841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X13252 a_9301_67503# a_9135_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13253 a_49402_15882# a_12727_13353# a_49894_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13254 a_20286_21906# a_11067_21583# a_20778_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13255 VSS a_11067_21583# a_49798_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13256 a_20286_17890# a_16362_17524# a_20378_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13257 a_5880_41641# a_4960_40847# a_5039_42167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13258 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X13259 a_9405_31599# a_8117_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1326 a_47486_70226# a_16746_70228# a_47394_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13260 vcm_commonmode a_16362_61190# a_35438_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13261 a_33338_20902# a_12985_7663# a_33830_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13262 a_33338_16886# a_16362_16520# a_33430_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13263 VSS a_8273_42479# a_9253_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13264 a_14081_37782# a_13909_37571# a_13867_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X13265 a_2417_52513# a_2199_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X13266 vcm_commonmode a_16362_71230# a_18370_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13267 VDD a_12901_58799# a_43378_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13268 VSS a_12727_15529# a_39758_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13269 a_36746_10862# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1327 a_11763_21237# a_9955_21807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=5.72e+06u as=0p ps=0u w=1e+06u l=150000u
X13270 a_43774_11866# a_12985_16367# a_43378_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13271 a_35319_34191# a_35142_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13272 VSS a_7563_46261# a_7494_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X13273 a_3026_19631# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13274 a_26802_15484# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13275 a_26706_21906# a_12985_7663# a_26310_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13276 a_23298_12870# a_12877_16911# a_23790_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13277 a_26319_41781# a_26495_41781# a_26447_41807# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X13278 VDD a_12877_16911# a_30326_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13279 VDD a_10515_22671# a_29322_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1328 a_15288_50639# a_7050_53333# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X13280 a_44382_66210# a_10975_66407# a_44874_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13281 vcm_commonmode a_16362_60186# a_39454_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13282 a_3137_27023# a_2315_24540# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13283 vcm_commonmode a_16362_19532# a_39454_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13284 a_2847_49855# a_2672_49929# a_3026_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13285 vcm_commonmode a_16362_14512# a_40458_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13286 a_8289_14741# a_8123_14741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13287 a_30567_49257# a_30534_49393# a_30485_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13288 a_19943_49007# a_14985_51701# a_19580_49159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13289 VDD a_5547_36495# a_5455_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1329 a_27710_68218# a_12901_66959# a_27314_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13290 a_12993_50095# a_6646_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X13291 a_11542_12381# a_11455_12157# a_11138_12267# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X13292 vcm_commonmode VSS a_23390_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13293 a_29718_12870# a_10055_58791# a_29322_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13294 a_36350_72234# VSS a_36442_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13295 a_12218_61341# a_11141_60975# a_12056_60975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13296 a_27314_11866# a_10055_58791# a_27806_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13297 a_40458_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13298 a_17274_68218# a_12727_67753# a_17766_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13299 a_16746_65208# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X133 a_7479_54439# a_23774_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X1330 VSS a_12355_65103# a_24698_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13300 a_21782_66532# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13301 a_16362_60186# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13302 a_16362_19532# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13303 VSS a_11747_28639# a_11710_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13304 a_7155_55509# a_7479_67075# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13305 a_9278_57487# a_8491_57487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13306 VDD a_11067_21583# a_39362_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13307 vcm_commonmode a_16362_15516# a_26402_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13308 a_29414_18528# a_16746_18526# a_29322_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13309 a_2700_43023# a_1757_43029# a_2592_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1331 VDD a_6782_58951# a_6739_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X13310 VSS a_27183_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13311 a_30418_13508# a_16746_13506# a_30326_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13312 a_10317_13647# a_9963_13760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13313 VSS VDD a_33734_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13314 a_4563_32900# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13315 result_out[7] a_1644_63669# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X13316 VSS a_29847_48734# a_29805_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13317 a_22294_62194# a_12355_15055# a_22786_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13318 VSS a_12901_66665# a_46786_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13319 VSS a_10515_22671# a_32730_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1332 a_9021_71677# a_8459_71285# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13320 a_42466_66210# a_16746_66212# a_42374_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13321 VSS a_5993_32687# a_6651_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13322 a_36328_49525# a_34145_49007# a_36720_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X13323 VSS a_4497_29673# a_5087_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13324 a_41370_21906# a_16362_21540# a_41462_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13325 a_44474_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13326 VSS a_24423_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13327 a_3019_13621# a_2847_15039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13328 a_26310_19898# a_11067_67279# a_26802_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13329 a_47486_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1333 VDD a_12899_11471# a_24302_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13330 a_12621_44099# a_21479_44581# a_22411_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X13331 a_40762_61190# a_12355_15055# a_40366_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13332 a_28810_56492# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13333 a_3529_25731# a_3325_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13334 a_30052_32117# a_30203_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X13335 a_23694_71230# a_12947_71576# a_23298_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13336 VDD a_12343_42333# a_12369_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X13337 a_46482_65206# a_16746_65208# a_46390_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13338 a_25355_40183# a_24423_40229# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13339 a_7387_69929# a_2689_65103# a_7637_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1334 vcm_commonmode a_16362_11500# a_39454_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13340 a_4001_56377# a_3668_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13341 a_45386_20902# a_16362_20536# a_45478_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13342 a_48490_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13343 a_32795_29967# a_32544_30083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13344 a_39391_47919# a_20635_29415# a_39222_48169# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X13345 VDD a_7939_30503# a_25759_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13346 VDD a_3031_47679# a_3018_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13347 a_36442_57174# a_16746_57176# a_36350_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13348 a_2163_57853# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13349 VDD a_12231_55509# a_12218_55901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1335 a_48398_13874# a_12727_15529# a_48890_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13350 a_37750_18894# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13351 VSS a_12899_11471# a_41766_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13352 VSS a_18105_40157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13353 a_19374_67214# a_16746_67216# a_19282_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13354 a_26112_30663# a_7862_34025# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13355 a_27710_70226# a_12901_66665# a_27314_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13356 a_49494_56170# a_16746_56172# a_49402_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13357 a_21686_23914# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13358 a_18278_22910# a_16362_22544# a_18370_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13359 VDD a_3417_31599# a_4233_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1336 a_6180_69929# a_6598_69653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13360 a_22386_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13361 a_27890_32459# a_5363_30503# a_27808_32459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13362 VDD a_31551_31751# a_30155_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X13363 a_17670_62194# a_12981_62313# a_17274_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13364 a_42374_59182# a_12901_58799# a_42866_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13365 VSS a_41351_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13366 a_10667_60735# a_10492_60809# a_10846_60797# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13367 a_2339_38129# a_2847_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13368 VSS a_12899_10927# a_27710_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13369 a_33830_70548# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1337 a_22386_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13370 a_22890_27247# a_17222_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13371 a_31726_15882# a_12877_14441# a_31330_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13372 VDD a_1761_32143# a_31959_34751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X13373 VSS a_12981_62313# a_40762_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13374 VDD a_1824_61127# a_1775_60663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X13375 a_2557_54447# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13376 a_37446_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13377 VDD VDD a_36350_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13378 a_7841_12167# a_53260_40156# a_53410_40254# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=0p ps=0u w=800000u l=150000u
X13379 a_8496_53359# a_7479_54439# a_8005_53333# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X1338 a_3123_53047# a_1952_60431# a_3297_53153# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13380 a_6373_15521# a_6155_15279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13381 a_43470_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13382 a_30720_49667# a_26397_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13383 VSS a_12473_36341# a_26495_36341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13384 a_3325_49551# a_2847_49855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13385 a_29322_8854# a_16362_8488# a_29414_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13386 a_24302_7850# VDD a_24794_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13387 VDD a_2325_36469# a_2215_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13388 a_31422_62194# a_16746_62196# a_31330_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13389 a_32826_58500# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1339 VDD a_2163_56765# a_2124_56891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13390 a_28714_13874# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13391 a_2325_44897# a_2107_44655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X13392 VSS a_10055_58791# a_32730_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13393 a_29414_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13394 a_2107_19631# a_1591_19631# a_2012_19631# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13395 a_18674_7850# VDD a_18278_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13396 a_19774_71552# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13397 a_30722_7850# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13398 a_4429_50095# a_3325_49551# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13399 a_19282_61190# a_16362_61190# a_19374_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X134 VSS a_1923_59583# a_2369_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1340 a_38850_19500# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13400 a_12353_20969# a_7377_18012# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13401 a_11599_65693# a_1950_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13402 a_2250_59343# a_2163_59585# a_1846_59475# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X13403 a_38378_30511# a_33694_30761# a_38292_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13404 a_47790_67214# a_12727_67753# a_47394_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13405 VDD a_5913_74273# a_5803_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13406 VSS a_11067_13095# a_44778_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13407 a_38358_23914# a_12947_23413# a_38850_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13408 a_38358_19898# a_16362_19532# a_38450_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13409 a_10221_74031# a_10055_74031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1341 a_42866_68540# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13410 a_11981_57487# a_11521_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13411 a_42866_21508# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13412 a_42466_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13413 a_30609_49159# a_30479_48576# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13414 a_4238_55123# a_4516_55107# a_4472_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13415 a_45386_65206# a_16362_65206# a_45478_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13416 a_27393_47919# a_26917_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X13417 VDD a_1586_9991# a_3247_10389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13418 VSS a_18413_47919# a_19258_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13419 a_37750_59182# a_12727_58255# a_37354_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1342 a_37446_62194# a_16746_62196# a_37354_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13420 VSS a_12947_56817# a_34738_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13421 VDD a_14926_31849# a_17507_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13422 VSS a_28648_50101# a_26662_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X13423 VDD a_12727_13353# a_35346_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13424 a_3885_28995# a_2011_34837# a_3789_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13425 VSS a_10975_66407# a_17670_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13426 a_6824_58799# a_6782_58951# a_6521_58773# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X13427 VSS a_2944_63400# a_2882_63517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X13428 a_7749_42479# a_6559_42479# a_7640_42479# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X13429 a_12323_51017# a_11877_50645# a_12227_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1343 VSS a_4811_34855# a_23727_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X13430 a_21686_64202# a_12355_65103# a_21290_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13431 VSS a_2847_19605# a_2781_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13432 a_16753_49007# a_16587_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13433 a_36442_10496# a_16746_10494# a_36350_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13434 VDD a_12877_14441# a_48398_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13435 a_45878_12472# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13436 a_2215_69135# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13437 a_43378_13874# a_16362_13508# a_43470_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13438 a_19374_20536# a_16746_20534# a_19282_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13439 a_22386_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1344 a_42283_39095# a_42188_37149# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X13440 a_23731_28023# a_2235_30503# a_23905_28129# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13441 VSS VSS a_38754_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13442 VSS config_2_in[0] a_1591_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13443 a_14737_47919# a_7000_43541# a_14655_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13444 a_34434_7484# VDD a_34342_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13445 a_22690_72234# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13446 VDD a_5682_69367# a_10289_55862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X13447 a_7839_21379# a_3339_43023# a_7757_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13448 a_17628_32143# a_17191_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13449 VDD a_11311_74005# a_8003_72917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1345 a_4771_42167# a_4446_40553# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X13450 VSS a_5877_70197# a_10615_72399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13451 a_45478_24552# VDD a_45386_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13452 VDD a_18487_28487# a_18126_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X13453 a_49402_66210# a_16362_66210# a_49494_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13454 a_5906_28335# a_5073_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X13455 a_19374_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13456 vcm_commonmode a_16362_66210# a_31422_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13457 a_8827_17215# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13458 a_7189_35015# a_4495_35925# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13459 a_49894_11468# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1346 a_29943_41317# a_28980_41831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X13460 a_20378_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13461 a_39854_68540# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13462 VDD a_20635_29415# a_41159_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X13463 a_28048_52093# a_6467_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13464 VSS a_27337_38565# a_27379_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13465 a_33338_24918# VSS a_33430_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13466 VDD a_12983_63151# a_43378_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13467 a_40858_63520# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13468 VSS a_40921_41245# a_40613_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13469 VDD a_14859_51183# a_15261_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1347 VDD a_2689_65103# a_4811_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13470 a_10595_30511# a_6459_30511# a_10506_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X13471 a_3107_46831# a_2959_47113# a_2744_46983# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X13472 a_10259_10703# a_9642_10357# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13473 a_35438_16520# a_16746_16518# a_35346_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13474 a_7000_43541# a_8384_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13475 a_3173_46805# a_2656_45895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X13476 VDD a_7571_29199# a_18579_27399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13477 vcm_commonmode VSS a_32426_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13478 VDD a_26523_29199# a_34337_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13479 a_43470_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1348 a_13867_35606# a_13909_35395# a_13867_35279# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13480 a_2859_41935# a_2235_41941# a_2751_42313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13481 a_11569_57711# a_11525_57953# a_11403_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X13482 a_2834_19997# a_1757_19631# a_2672_19631# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13483 VDD a_32367_28309# a_36797_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X13484 a_26402_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13485 a_25398_9492# a_16746_9490# a_25306_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13486 a_11136_74031# a_10221_74031# a_10789_74273# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13487 VDD a_12985_16367# a_26310_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13488 VSS a_14625_30761# a_15812_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13489 a_6608_19319# a_4792_20443# a_6750_19126# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X1349 a_8123_56399# a_10687_52553# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13490 a_22562_28023# a_22441_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X13491 VDD a_10975_66407# a_47394_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13492 a_44874_62516# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13493 VSS a_12473_42869# a_24931_42657# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13494 a_17869_28335# a_15799_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13495 a_26778_29473# a_27016_29587# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X13496 a_5367_34435# a_2216_28309# a_5271_34435# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13497 VDD a_1642_22583# a_1591_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13498 a_30816_35077# a_29943_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13499 a_29718_62194# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X135 VSS a_7815_49855# a_7749_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X1350 VSS a_12947_56817# a_27710_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13500 vcm_commonmode a_16362_57174# a_25398_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13501 a_33727_36649# a_32795_36415# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13502 a_30105_32463# a_30052_32117# a_29887_32375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13503 VDD a_18662_43671# a_18667_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13504 a_30722_16886# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13505 VDD a_10515_22671# a_37354_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13506 a_7903_48841# a_7387_48469# a_7808_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X13507 a_47790_20902# a_11067_67279# a_47394_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13508 a_17766_64524# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13509 VDD a_12981_62313# a_21290_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1351 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X13510 a_42770_69222# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13511 a_17475_51157# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13512 a_37750_12870# a_10055_58791# a_37354_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13513 VSS a_21948_34973# a_22411_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13514 vcm_commonmode a_16362_23548# a_44474_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13515 a_9951_68367# a_9914_68279# a_8772_63927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13516 a_13643_28327# a_32823_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X13517 VSS a_13565_44135# a_13510_44759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13518 a_22294_70226# a_12516_7093# a_22786_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13519 a_43378_58178# a_16362_58178# a_43470_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1352 vcm_commonmode a_16362_8488# a_29414_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13520 a_11155_30663# a_10761_29745# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13521 a_13716_43047# a_33015_40513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X13522 a_41878_31375# a_28757_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X13523 a_7171_62313# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13524 a_18278_60186# a_12727_58255# a_18770_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13525 a_38358_9858# a_16362_9492# a_38450_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13526 a_26310_68218# a_16362_68218# a_26402_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13527 VSS a_33486_34191# a_34859_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13528 a_49984_39288# a_49750_39288# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.394e+11p pd=2.82e+06u as=0p ps=0u w=420000u l=150000u M=2
X13529 vcm_commonmode a_16362_15516# a_34434_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1353 VDD a_12355_15055# a_12727_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X13530 a_43378_17890# a_12899_10927# a_43870_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13531 a_12323_20904# a_7377_18012# a_12709_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X13532 a_32334_11866# a_16362_11500# a_32426_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13533 a_29416_31171# a_8491_41383# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13534 a_17943_30761# a_17651_30485# a_7295_44647# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=0p ps=0u w=1e+06u l=150000u
X13535 VDD a_9613_13077# a_9643_13430# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13536 a_2781_12937# a_1591_12565# a_2672_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13537 a_28980_41831# a_28011_41855# a_28884_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13538 VSS a_7072_56053# a_6072_56872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X13539 a_3509_58487# a_3714_58345# a_3672_58371# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1354 a_40458_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13540 a_21382_23548# a_16746_23546# a_21290_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13541 VSS a_5682_69367# a_10296_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13542 a_77285_40202# a_77381_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13543 a_20378_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13544 a_34434_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13545 a_36746_18894# a_12899_10927# a_36350_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13546 a_33668_44007# a_32795_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13547 VDD a_27560_34337# a_26661_34428# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X13548 a_15103_49525# a_15439_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13549 vcm_commonmode a_16362_70226# a_43470_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1355 a_16362_11500# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X13550 a_2685_59933# a_1954_61677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13551 VDD a_13669_37429# a_14081_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13552 VSS a_12727_67753# a_23694_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13553 a_20682_65206# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13554 a_49798_59182# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13555 VDD a_3987_19623# a_6993_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13556 a_49798_17890# a_12899_11471# a_49402_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13557 a_42188_37149# a_41351_39141# a_42224_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13558 VSS a_2775_46025# a_32582_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13559 a_20778_17492# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1356 VDD a_12727_13353# a_28318_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13560 VDD a_9314_69367# a_10699_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13561 a_47394_16886# a_12899_11471# a_47886_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13562 VDD a_11430_26159# a_13335_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13563 VSS a_41842_27221# a_42887_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13564 a_34342_19898# a_11067_67279# a_34834_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13565 a_33734_64202# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13566 a_10317_30287# a_8273_42479# a_9963_29967# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X13567 a_36735_49257# a_35568_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13568 a_4692_55541# a_1823_58773# a_4620_55541# VSS sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X13569 VDD a_3016_60949# a_3621_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1357 a_10045_21379# a_6559_22671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13570 a_22351_47893# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13571 a_31330_21906# a_11067_21583# a_31822_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13572 a_31330_17890# a_16362_17524# a_31422_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13573 a_38450_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13574 VDD a_12727_58255# a_41370_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13575 vcm_commonmode VSS a_16362_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13576 VSS a_12877_14441# a_37750_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13577 a_19128_48829# a_18413_47919# a_18907_48502# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X13578 a_20378_70226# a_16746_70228# a_20286_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13579 vcm_commonmode a_16362_61190# a_46482_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1358 a_25798_13476# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13580 VSS a_12901_58799# a_26706_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13581 a_23694_56170# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13582 a_30722_57174# a_10515_22671# a_30326_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13583 a_24794_16488# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13584 a_21290_13874# a_12727_15529# a_21782_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13585 a_10035_60431# a_9411_60437# a_9927_60809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13586 VDD a_30412_42589# a_29513_42333# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X13587 a_42374_67214# a_12983_63151# a_42866_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13588 a_28410_13508# a_16746_13506# a_28318_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13589 vcm_commonmode a_16362_10496# a_25398_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1359 a_13809_48463# a_13461_48579# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X13590 VSS a_4215_51157# a_26155_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13591 VDD a_2952_66139# a_7479_67075# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13592 a_23390_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13593 VSS a_38345_42044# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13594 a_10665_58487# a_6417_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13595 a_27710_55166# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13596 VSS a_9367_29397# a_9355_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13597 a_46786_9858# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13598 a_42770_22910# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13599 a_39362_21906# a_16362_21540# a_39454_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X136 VDD a_1586_66567# a_10975_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1360 a_4259_41167# a_3949_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X13600 VDD a_1887_34863# a_2289_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13601 a_37919_28111# a_36904_28879# a_37747_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X13602 VSS a_2592_43023# a_3162_43023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13603 a_28318_68218# a_12727_67753# a_28810_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13604 a_39758_66210# a_12983_63151# a_39362_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13605 a_18844_43439# a_18667_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13606 a_11403_57711# a_10957_57711# a_11307_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13607 a_32826_66532# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13608 a_27406_60186# a_16746_60188# a_27314_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13609 a_2704_16911# a_1757_16917# a_2596_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1361 a_16707_44535# a_15775_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X13610 a_27406_19532# a_16746_19530# a_27314_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13611 VSS a_1586_9991# a_1591_14741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13612 a_5190_59575# a_14985_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X13613 a_32334_56170# a_16362_56170# a_32426_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13614 a_16362_21540# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X13615 VSS a_10472_26159# a_12300_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X13616 a_37557_32463# a_27535_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13617 VSS a_32121_42369# a_33727_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13618 VSS a_2865_58799# a_2882_59343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X13619 a_41059_32143# a_31659_31751# a_41141_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X1362 a_7352_35113# a_4495_35925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13620 VDD a_3023_16341# a_2899_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X13621 a_37427_47893# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X13622 a_49402_57174# a_12257_56623# a_49894_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13623 vcm_commonmode a_16362_69222# a_36442_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13624 a_12056_55535# a_11141_55535# a_11709_55777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13625 VSS VDD a_44778_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13626 a_40458_67214# a_16746_67216# a_40366_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13627 a_33338_62194# a_12355_15055# a_33830_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13628 a_12818_52521# a_12202_54599# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13629 VSS a_32318_48695# a_32319_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1363 VDD a_3112_9527# a_3063_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13630 a_33734_9858# a_12985_19087# a_33338_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13631 a_2080_54813# a_1643_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13632 a_19678_23914# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13633 VSS a_13669_37429# a_14088_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13634 a_49798_12870# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13635 VSS a_11067_21583# a_23694_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13636 a_39272_31573# a_8491_41383# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13637 VSS a_9424_60949# a_9370_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13638 VSS a_1925_18231# a_1738_17973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13639 a_4343_60405# a_4187_60673# a_4488_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X1364 VSS a_41211_28023# a_39727_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13640 a_26802_57496# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13641 a_12174_12381# a_11416_12283# a_11611_12252# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13642 VDD VSS a_30326_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13643 a_21686_72234# VDD a_21290_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13644 a_11513_53609# a_6095_44807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X13645 a_26508_40969# a_24561_41583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13646 a_37423_51335# a_37512_50755# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13647 a_2886_53686# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X13648 a_7009_56873# a_1823_66941# a_6927_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13649 a_7060_61225# a_5024_67885# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1365 VDD a_2787_32679# a_8461_32937# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X13650 VSS a_12546_22351# a_31726_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13651 a_34482_29941# a_37503_31393# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X13652 a_24991_28129# a_23195_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13653 VSS a_12877_16911# a_26706_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13654 VSS a_12981_62313# a_38754_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13655 a_35742_60186# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13656 a_34434_58178# a_16746_58180# a_34342_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13657 a_35742_19898# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13658 a_30722_10862# a_12546_22351# a_30326_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13659 vcm_commonmode a_16362_9492# a_48490_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1366 a_46882_67536# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13660 VDD a_4461_48981# a_4491_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13661 a_16707_36919# a_15775_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13662 a_18674_70226# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13663 a_17366_68218# a_16746_68220# a_17274_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13664 a_2620_43389# a_2040_43401# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13665 VDD a_1923_73087# a_2464_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13666 a_5225_58621# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13667 a_42374_7850# VSS a_42466_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13668 a_47486_57174# a_16746_57176# a_47394_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13669 a_48794_18894# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1367 a_43378_64202# a_11067_13095# a_43870_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13670 VSS a_30412_42589# a_35099_43447# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X13671 VDD a_6835_46823# a_26341_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13672 VDD a_26523_28111# a_35601_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X13673 VSS a_1923_73087# a_2369_69501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13674 a_12565_9633# a_11067_67279# a_12479_9633# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13675 a_9075_72737# a_7707_70741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13676 a_36842_22512# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13677 VSS a_28931_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X13678 a_40858_71552# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13679 VDD a_11067_67279# a_40366_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1368 a_29414_10496# a_16746_10494# a_29322_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13680 VSS a_19096_44129# a_18197_44220# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X13681 VDD a_12355_65103# a_39362_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13682 a_43470_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13683 a_40366_61190# a_16362_61190# a_40458_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13684 a_2319_56860# a_2124_56891# a_2629_56623# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X13685 VSS a_3143_66972# a_5484_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X13686 a_4717_65569# a_4499_65327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X13687 a_28714_62194# a_12981_62313# a_28318_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13688 a_28410_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13689 a_23298_71230# a_16362_71230# a_23390_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1369 a_16362_8488# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X13690 a_5274_54991# a_4555_55233# a_4711_54965# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X13691 VSS a_12895_13967# a_25702_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13692 a_2635_55329# a_1591_54447# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13693 a_7075_45577# a_6559_45205# a_6980_45565# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13694 a_44874_70548# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13695 a_37354_14878# a_16362_14512# a_37446_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13696 VSS a_7571_29199# a_11711_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13697 a_16955_52047# a_38067_47349# a_37839_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X13698 a_41462_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13699 a_5405_25615# a_5309_25853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X137 a_41370_67214# a_12983_63151# a_41862_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1370 VSS a_16244_34973# a_16707_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13700 VDD a_33080_37149# a_33668_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X13701 a_41766_69222# a_12516_7093# a_41370_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13702 a_44382_60186# a_16362_60186# a_44474_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13703 VDD a_3541_9593# a_3571_9334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13704 VDD a_12473_41781# a_12417_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13705 a_27314_70226# a_16362_70226# a_27406_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13706 a_30818_59504# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13707 a_26706_14878# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13708 VSS a_13047_29575# a_12999_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13709 vcm_commonmode a_16362_22544# a_36442_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1371 VDD a_1644_62037# result_out[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X13710 a_8129_29967# a_4495_35925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13711 a_2847_66389# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13712 VSS a_5535_18012# a_11564_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X13713 a_17766_72556# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13714 a_40458_20536# a_16746_20534# a_40366_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13715 VDD a_12985_7663# a_17274_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13716 VDD a_12901_66665# a_21290_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13717 VDD a_12546_22351# a_47394_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13718 VSS a_8583_33551# a_19439_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X13719 a_17274_62194# a_16362_62194# a_17366_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1372 a_1757_23445# a_1591_23445# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13720 a_38754_67214# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13721 a_10575_62911# a_10400_62985# a_10754_62973# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13722 a_21382_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13723 a_45782_68218# a_12901_66959# a_45386_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13724 VSS a_12355_65103# a_42770_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13725 VDD a_12757_8207# a_12815_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13726 VSS a_10073_23439# a_11390_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X13727 a_40458_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13728 a_12713_20495# a_5535_18012# a_12166_21501# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13729 VSS a_11947_68279# a_11771_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1373 a_4974_56875# a_5291_56765# a_5249_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X13730 vcm_commonmode a_16362_66210# a_29414_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13731 a_2886_53359# a_2840_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13732 a_18370_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13733 a_38850_63520# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13734 a_48794_59182# a_12727_58255# a_48398_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13735 VSS a_12947_56817# a_45782_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13736 a_2107_45577# a_1757_45205# a_2012_45565# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X13737 a_16992_50959# a_13445_50639# a_16902_50639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X13738 VDD a_12355_15055# a_42374_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13739 VDD a_75445_40202# a_75258_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1374 VSS a_12947_23413# a_33734_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13740 VDD a_12727_13353# a_46390_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13741 a_34434_11500# a_16746_11498# a_34342_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13742 VSS a_7313_53047# a_7271_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X13743 a_23390_56170# a_16746_56172# a_23298_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13744 a_24698_17890# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13745 VDD a_12895_13967# a_33338_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13746 a_17366_21540# a_16746_21538# a_17274_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13747 VDD a_2847_21781# a_2834_22173# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13748 VSS a_5363_30503# a_27387_32373# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13749 a_47486_10496# a_16746_10494# a_47394_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1375 a_32730_62194# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13750 a_4514_58387# a_4792_58371# a_4748_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13751 a_34342_68218# a_16362_68218# a_34434_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13752 a_8544_15101# a_8361_15529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13753 a_9931_69513# a_9485_69141# a_9835_69513# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X13754 a_7407_18365# a_7153_18038# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13755 VDD a_12899_10927# a_19282_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13756 a_47394_67214# a_16362_67214# a_47486_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13757 VSS VSS a_49798_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13758 VDD config_2_in[14] a_1591_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13759 a_33486_34191# a_33309_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1376 VSS a_35932_37601# a_36579_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13760 a_33734_72234# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13761 a_37846_69544# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13762 a_13620_40871# a_12801_38517# a_13762_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13763 VDD a_12727_67753# a_41370_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13764 VDD a_20535_51727# a_22015_51840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13765 VSS a_15607_46805# a_30975_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13766 a_17394_32275# a_17711_32385# a_17669_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X13767 a_9707_51325# a_1586_51335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13768 VDD a_1923_59583# a_4488_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13769 a_37354_59182# a_16362_59182# a_37446_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1377 a_29322_67214# a_16362_67214# a_29414_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13770 VSS a_77568_39738# a_77381_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13771 a_41462_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13772 a_24394_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13773 a_26706_55166# VSS a_26310_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13774 a_41766_22910# a_11067_21583# a_41370_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13775 a_22632_42919# a_21663_42943# a_22536_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13776 a_38358_65206# a_12355_65103# a_38850_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13777 a_27710_63198# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13778 vcm_commonmode a_16362_58178# a_23390_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13779 vcm_commonmode a_16362_71230# a_37446_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1378 VDD VDD a_21290_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13780 a_2283_15797# a_3166_16911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13781 VDD a_32365_37692# a_31971_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13782 a_38754_20902# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13783 VDD a_1823_63677# a_5541_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X13784 a_3697_72719# a_2686_70223# a_2747_72007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13785 a_25204_39655# a_24331_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X13786 a_42374_12870# a_12877_16911# a_42866_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13787 a_45782_21906# a_12985_7663# a_45386_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13788 a_5411_68086# a_5160_68315# a_4952_68279# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13789 VDD a_12703_38517# a_12341_41281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1379 a_3883_24643# a_2317_28892# a_3801_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13790 a_8379_74575# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X13791 VDD a_10515_22671# a_48398_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13792 a_25306_22910# a_10515_23975# a_25798_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13793 a_20685_28335# a_15661_29199# a_21140_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13794 a_18370_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13795 a_15548_30761# a_14361_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X13796 VSS a_7815_19319# a_7756_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13797 a_5913_48161# a_5695_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X13798 a_32334_64202# a_16362_64202# a_32426_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X13799 a_35742_13874# a_12877_16911# a_35346_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X138 a_27406_13508# a_16746_13506# a_27314_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1380 VDD a_28757_27247# a_30748_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3e+11p ps=5.26e+06u w=1e+06u l=150000u M=2
X13800 a_6553_16367# a_5363_16367# a_6444_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13801 a_2847_30271# a_2672_30345# a_3026_30333# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13802 a_8259_18543# a_8111_18825# a_7896_18695# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X13803 vcm_commonmode VSS a_42466_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13804 a_18770_17492# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13805 a_18674_23914# a_10515_23975# a_18278_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13806 a_4952_68279# a_5160_68315# a_5094_68413# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13807 VDD a_12877_14441# a_22294_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13808 a_48794_12870# a_10055_58791# a_48398_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13809 a_25321_29423# a_9529_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1381 a_5550_58255# a_4831_58497# a_4987_58229# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X13810 a_38076_31573# a_35815_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13811 VDD a_12725_44527# a_27983_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13812 a_29322_21906# a_11067_21583# a_29814_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13813 a_28733_28585# a_23928_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13814 a_33338_70226# a_12516_7093# a_33830_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13815 a_29322_17890# a_16362_17524# a_29414_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13816 a_8256_20969# a_7377_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13817 a_41370_18894# a_12895_13967# a_41862_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13818 a_30326_12870# a_16362_12504# a_30418_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13819 VSS a_15828_38695# a_15193_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1382 VDD a_10515_22671# a_40366_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13820 a_27388_49007# a_26662_48981# a_26218_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X13821 VSS a_2292_17179# a_8349_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13822 a_18370_70226# a_16746_70228# a_18278_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13823 a_2657_60949# a_2497_61519# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13824 VSS a_12901_66959# a_30722_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13825 vcm_commonmode a_16362_15516# a_45478_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13826 a_48490_18528# a_16746_18526# a_48398_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13827 a_19282_13874# a_12727_15529# a_19774_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13828 a_34738_60186# a_12981_59343# a_34342_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13829 a_23790_11468# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1383 VSS a_10515_23975# a_46786_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13830 a_34738_19898# a_12895_13967# a_34342_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X13831 a_14421_49007# a_13809_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X13832 a_32426_23548# a_16746_23546# a_32334_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13833 VSS a_5023_13255# a_4995_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13834 VDD a_28980_41831# a_28884_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X13835 a_4181_50345# a_4127_50069# a_3983_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X13836 a_16843_51549# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X13837 a_45478_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13838 VSS a_1923_54591# a_4549_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X13839 VDD a_16928_36391# a_16832_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1384 a_26860_41605# a_25987_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X13840 VSS a_10964_25615# a_13527_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X13841 VDD a_2944_64488# a_2882_64605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X13842 vcm_commonmode a_16362_17524# a_18370_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13843 a_37527_29397# a_38378_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13844 a_35036_34191# a_34859_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13845 VDD a_4191_33449# a_16587_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13846 VDD a_3751_72373# a_6835_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X13847 a_8453_64757# a_8782_65015# a_8740_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13848 a_31726_65206# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13849 a_22386_15516# a_16746_15514# a_22294_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1385 a_19774_69544# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13850 VSS a_5259_39367# a_3759_39991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13851 vcm_commonmode a_16362_14512# a_49494_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13852 a_40457_27765# a_40086_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13853 a_1915_21482# a_2007_21237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X13854 a_28405_52093# a_28361_51701# a_28239_52105# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X13855 a_45386_19898# a_11067_67279# a_45878_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13856 a_39854_8456# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13857 a_35742_8854# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13858 a_21686_57174# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13859 a_7561_36815# a_7001_36495# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1386 VDD a_12727_67753# a_23298_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13860 a_49494_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13861 a_42770_71230# a_12947_71576# a_42374_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13862 VSS a_5136_34551# a_5079_35639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X13863 a_6271_72943# a_6224_73095# a_6182_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13864 a_27314_63198# a_12981_62313# a_27806_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13865 VDD a_10471_65002# a_8999_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13866 VDD VDD a_39362_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13867 a_31822_61512# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13868 VDD a_12947_8725# a_49402_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13869 VSS a_12985_19087# a_45782_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1387 a_20778_64524# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13870 a_26402_14512# a_16746_14510# a_26310_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13871 vcm_commonmode a_16362_11500# a_23390_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13872 VSS a_1586_51335# a_9411_60437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13873 a_35568_49525# a_2959_47113# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X13874 a_39454_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13875 a_22786_19500# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13876 a_14298_32143# a_14354_32117# a_14298_32463# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X13877 VSS a_30573_52271# a_30849_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13878 a_1761_25071# a_1591_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X13879 a_3049_14343# a_3019_13621# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1388 a_19282_59182# a_16362_59182# a_19374_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13880 a_38450_67214# a_16746_67216# a_38358_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13881 vcm_commonmode a_16362_64202# a_35438_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13882 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=5.1e+06u w=1.89e+07u
X13883 a_40762_23914# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13884 VDD a_13620_43047# a_12889_40977# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X13885 a_37354_22910# a_16362_22544# a_37446_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13886 a_7755_70223# a_2689_65103# a_8531_70543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X13887 VDD a_12231_65301# a_12218_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13888 a_11803_29967# a_8485_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X13889 a_41462_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1389 VSS a_7571_29199# a_20747_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X13890 a_7539_63695# a_6913_64239# a_7445_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X13891 a_3305_38671# a_2847_38975# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X13892 a_30375_51335# a_30947_51157# a_30720_51183# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X13893 a_26310_69222# a_12901_66959# a_26802_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13894 VSS a_2339_38129# a_5588_22467# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13895 a_41636_37601# a_41351_38053# a_42224_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13896 a_30818_67536# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13897 VSS a_12895_13967# a_33734_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13898 VSS a_12889_35537# a_12921_35279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13899 VSS a_32887_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X139 a_13173_29673# a_13390_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.55e+11p pd=5.31e+06u as=0p ps=0u w=1e+06u l=150000u
X1390 a_23390_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13900 a_9503_26151# a_41597_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X13901 a_17257_46859# a_4443_46607# a_17171_46859# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X13902 a_30326_57174# a_16362_57174# a_30418_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13903 a_7373_40847# a_7107_40847# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13904 VSS a_12899_10927# a_46786_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13905 a_2215_71311# a_1591_71317# a_2107_71689# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X13906 a_9872_20175# a_10275_21495# a_10311_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X13907 a_5529_11471# a_4812_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13908 a_4145_60797# a_3667_60405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X13909 a_7259_31375# a_5449_25071# a_7125_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1391 a_12447_29199# a_18162_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X13910 a_39223_32463# a_39113_32204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13911 VDD a_3295_54421# a_10791_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13912 VSS a_10515_23975# a_30722_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13913 a_27406_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13914 a_12263_26409# a_9955_20969# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13915 a_31543_51335# a_29361_51727# a_31669_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13916 a_18278_7850# VDD a_18770_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13917 a_34738_14878# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13918 VDD a_2007_65002# a_1895_66628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X13919 a_8206_28879# a_6649_25615# a_8123_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X1392 a_2199_52271# a_1683_52271# a_2104_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13920 a_2847_38975# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13921 a_2744_53511# a_2177_53359# a_2886_53686# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X13922 vcm_commonmode a_16362_8488# a_37446_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13923 a_17670_24918# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13924 a_23694_17890# a_12899_11471# a_23298_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13925 a_47790_13874# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13926 a_30722_8854# a_12947_8725# a_30326_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13927 a_23507_44265# a_23901_44220# a_23567_44211# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X13928 a_48490_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13929 a_38850_71552# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1393 a_11801_68047# a_11771_68021# a_8782_65015# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X13930 a_21290_55166# VSS a_21782_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13931 a_27155_40871# a_12725_44527# a_27329_40747# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13932 a_47486_8488# a_16746_8486# a_47394_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13933 VSS a_3305_38671# a_5631_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X13934 vcm_commonmode a_16362_61190# a_20378_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13935 a_6369_47919# a_5179_47919# a_6260_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X13936 a_14445_50095# a_9963_50959# a_14373_50095# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X13937 a_5963_20149# a_8256_20969# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13938 VSS a_11719_28023# a_11747_28639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13939 a_27710_16886# a_12727_13353# a_27314_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1394 VSS a_5211_24759# a_5449_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u M=4
X13940 VSS a_12727_15529# a_24698_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13941 a_21686_10862# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13942 a_4053_35523# a_2216_28309# a_3980_35523# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X13943 a_5723_27497# a_5085_23047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X13944 a_33688_46831# a_18979_30287# a_33385_46805# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X13945 a_1757_44655# a_1591_44655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X13946 VSS a_12981_62313# a_49798_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13947 VDD a_32167_29611# a_32125_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13948 VDD a_5831_39189# a_8357_44982# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X13949 a_46786_60186# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1395 a_40762_12870# a_10055_58791# a_40366_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13950 a_45478_58178# a_16746_58180# a_45386_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X13951 a_22294_8854# a_16362_8488# a_22386_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X13952 a_46786_19898# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13953 VSS a_6607_13879# a_6327_14343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13954 VSS a_10975_66407# a_36746_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13955 a_2882_59343# a_2163_59585# a_2319_59317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13956 a_37076_37253# a_36107_36965# a_36980_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X13957 a_32370_50871# a_29361_51727# a_32507_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13958 a_1644_58773# a_1823_58773# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13959 a_40762_64202# a_12355_65103# a_40366_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1396 a_23507_35561# a_23901_35516# a_23567_35507# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X13960 vcm_commonmode a_16362_60186# a_24394_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13961 vcm_commonmode a_16362_19532# a_24394_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13962 a_34834_23516# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13963 a_28810_59504# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13964 a_34434_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13965 a_9114_13763# a_9083_13879# a_9041_13763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13966 a_32426_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13967 VDD a_2216_42997# a_2126_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.89e+11p ps=1.74e+06u w=420000u l=150000u
X13968 VSS a_12757_9295# a_12815_7663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13969 a_38450_20536# a_16746_20534# a_38358_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1397 VDD a_3063_34319# a_3607_34639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X13970 VSS a_7833_66415# a_8491_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X13971 a_41462_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13972 a_47886_22512# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13973 VSS a_22063_47594# a_19788_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X13974 a_37446_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13975 a_21290_72234# VSS a_21382_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13976 a_26706_63198# a_15439_49525# a_26310_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13977 a_6653_36611# a_5631_38127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13978 a_29220_50639# a_27869_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13979 a_5023_72068# a_7100_72105# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1398 VSS a_1586_69367# a_1591_69141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13980 a_8219_54447# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13981 a_37846_14480# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13982 VDD a_36328_49525# a_35403_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X13983 a_38450_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X13984 a_35346_15882# a_16362_15516# a_35438_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13985 VDD a_10055_58791# a_41370_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13986 a_2873_31599# a_1683_31599# a_2764_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X13987 VSS a_40585_42369# a_42099_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X13988 VDD a_11067_21583# a_24302_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X13989 a_48398_14878# a_16362_14512# a_48490_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1399 a_4831_52413# a_1586_51335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13990 vcm_commonmode VSS a_26402_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13991 a_13335_27497# a_12349_25847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13992 a_7159_22583# a_7431_22441# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13993 VDD a_1586_40455# a_2235_41941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X13994 a_17670_65206# a_10975_66407# a_17274_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13995 VSS a_77568_40202# a_77381_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X13996 a_9209_24527# a_7203_24527# a_9125_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13997 a_38358_10862# a_12985_16367# a_38850_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13998 a_2007_10901# a_1887_10422# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X13999 VSS a_12473_42869# a_12892_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VSS a_2375_49172# a_1895_49722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X140 VSS a_3452_70537# a_3410_70589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1400 a_37354_55166# VSS a_37846_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14000 VSS a_12901_66665# a_31726_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14001 VDD a_12985_16367# a_45386_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14002 VDD a_12901_66959# a_35346_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14003 VDD a_3339_43023# a_3983_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14004 a_36746_68218# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14005 a_9123_55223# a_8453_51727# a_9290_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14006 VDD a_12985_7663# a_28318_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14007 VSS a_31280_40517# a_31243_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14008 a_1757_45205# a_1591_45205# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14009 a_46390_9858# a_12546_22351# a_46882_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1401 a_5959_13621# a_5755_14709# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14010 VSS a_6393_34837# a_6327_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14011 a_25398_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14012 a_36717_47375# a_36448_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X14013 a_1757_14741# a_1591_14741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X14014 a_28318_62194# a_16362_62194# a_28410_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14015 a_24331_34239# a_20715_34717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X14016 a_32426_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14017 VDD a_7803_55509# a_8162_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14018 vcm_commonmode a_16362_57174# a_44474_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14019 VSS a_8575_74853# a_8533_74941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1402 a_23694_22910# a_11067_21583# a_23298_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14020 VDD a_12877_16911# a_18278_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14021 vcm_commonmode a_16362_67214# a_27406_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14022 a_31422_65206# a_16746_65208# a_31330_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14023 a_31059_38007# a_30127_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14024 VSS a_9731_22895# a_13081_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14025 a_36842_64524# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14026 a_30326_20902# a_16362_20536# a_30418_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14027 a_4627_27613# a_3325_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14028 a_2781_40303# a_1591_40303# a_2672_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X14029 a_41370_69222# a_16362_69222# a_41462_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1403 VDD a_2672_9839# a_2847_9813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14030 VDD a_12981_62313# a_40366_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14031 a_29414_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14032 a_8297_31055# a_2787_32679# a_8215_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14033 VDD a_7815_42453# a_7802_42845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14034 VDD a_12381_43957# a_12325_44310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14035 a_12683_51329# a_13445_50639# a_14005_50959# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14036 vcm_commonmode a_16362_59182# a_17366_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14037 a_49894_63520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14038 VSS a_8295_47388# a_12899_3311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X14039 a_21382_57174# a_16746_57176# a_21290_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1404 a_7841_12167# a_53260_40156# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.604e+11p pd=2.92e+06u as=0p ps=0u w=420000u l=150000u
X14040 a_22690_18894# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14041 a_35076_51183# a_35039_51335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14042 VSS a_5831_39189# a_8364_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14043 a_45478_11500# a_16746_11498# a_45386_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14044 a_18307_27791# a_17774_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X14045 a_7187_37583# a_6559_37583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14046 VDD a_12895_13967# a_44382_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14047 a_4499_65327# a_4149_65327# a_4404_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X14048 a_2012_33927# a_4503_21523# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X14049 VDD a_12985_19087# a_33338_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1405 a_21290_60186# a_12727_58255# a_21782_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14050 a_34780_56398# a_34987_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X14051 a_37354_60186# a_12727_58255# a_37846_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14052 a_45386_68218# a_16362_68218# a_45478_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14053 VSS a_7019_35951# a_5490_41365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X14054 a_27425_47695# a_4891_47388# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14055 a_41697_27497# a_41842_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14056 VDD a_15439_49525# a_26310_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14057 a_5039_47741# a_4891_47388# a_4676_47607# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14058 a_24055_36415# a_22448_37253# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14059 a_3871_10383# a_3247_10389# a_3763_10761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1406 a_5421_60137# a_5333_59343# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X14060 VDD a_26465_48463# a_27929_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14061 VSS a_7865_46805# a_7799_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14062 a_30165_47695# a_26514_47375# a_29847_48734# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14063 a_18177_32509# a_17798_32143# a_18105_32509# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X14064 a_2369_36861# a_2325_36469# a_2203_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X14065 VSS a_9367_29397# a_11711_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X14066 VSS a_22989_48437# a_26225_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X14067 a_31822_9460# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14068 a_25764_51183# a_24849_51183# a_25417_51425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14069 a_6878_30287# a_6649_25615# a_6788_30287# VSS sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=0p ps=0u w=650000u l=150000u
X1407 a_16879_37999# a_16699_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14070 a_27263_40871# a_1761_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14071 a_27314_71230# a_12901_66665# a_27806_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14072 a_22386_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14073 a_48398_59182# a_16362_59182# a_48490_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14074 VDD a_13669_35253# a_13613_35606# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14075 VDD a_8373_26409# a_10055_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X14076 VSS a_12907_27023# a_13183_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14077 a_25317_49007# a_14831_50095# a_23631_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14078 a_8491_67279# a_5682_69367# a_7580_61751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X14079 vcm_commonmode VSS a_35438_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1408 a_48794_72234# VDD a_48398_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14080 a_20853_47375# a_20575_47713# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14081 a_25398_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14082 VDD a_2244_18231# a_2021_17973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14083 VDD a_6752_29941# a_8827_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14084 a_42770_56170# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14085 a_39362_18894# a_12895_13967# a_39854_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14086 a_36746_21906# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14087 VSS VSS a_39758_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14088 vcm_commonmode a_16362_71230# a_48490_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14089 a_4149_65327# a_3983_65327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1409 VSS a_4960_40847# a_5962_41391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X14090 a_5378_56989# a_5291_56765# a_4974_56875# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14091 a_43870_16488# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14092 a_40366_13874# a_12727_15529# a_40858_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14093 VSS a_12901_66959# a_28714_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14094 a_25702_66210# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14095 a_23298_23914# a_12947_23413# a_23790_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14096 a_23298_19898# a_16362_19532# a_23390_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14097 vcm_commonmode a_16362_10496# a_44474_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14098 a_17366_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14099 VDD a_38345_42044# a_37951_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X141 a_7289_70767# a_5877_70197# a_7651_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X1410 VDD a_10073_23439# a_10526_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X14100 vcm_commonmode a_16362_20536# a_27406_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14101 VSS a_38315_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X14102 a_33734_14878# a_12727_15529# a_33338_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14103 a_30326_65206# a_16362_65206# a_30418_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14104 a_42466_61190# a_16746_61192# a_42374_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14105 a_29414_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14106 a_26310_55166# VSS a_26402_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14107 a_5331_18517# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14108 a_3301_26703# a_2315_24540# a_3229_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14109 a_22690_59182# a_12727_58255# a_22294_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1411 vcm_commonmode a_16362_71230# a_19374_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14110 a_16666_24918# VSS a_16270_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14111 VDD a_5239_45717# a_4758_45369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X14112 a_41443_41855# a_38011_42035# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X14113 VDD a_35568_49525# a_37926_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14114 a_30565_30199# a_40691_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14115 a_25398_71230# a_16746_71232# a_25306_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14116 a_32311_48169# a_27869_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14117 VDD a_12727_13353# a_20286_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14118 a_46786_13874# a_12877_16911# a_46390_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14119 a_29718_65206# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1412 VDD a_9491_12297# a_10299_11703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14120 a_34342_69222# a_12901_66959# a_34834_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14121 vcm_commonmode a_16362_12504# a_17366_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14122 a_29814_17492# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14123 a_29718_23914# a_10515_23975# a_29322_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14124 a_34906_47491# a_34062_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14125 a_26310_14878# a_12877_14441# a_26802_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14126 a_21382_10496# a_16746_10494# a_21290_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14127 a_27314_18894# a_16362_18528# a_27406_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14128 a_30818_12472# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14129 a_39247_39095# a_38315_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1413 a_37750_10862# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14130 VSS a_1761_52815# a_26267_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14131 a_3327_9308# a_4503_10687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14132 a_47394_68218# a_12727_67753# a_47886_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14133 a_1929_12131# a_2847_12863# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14134 VSS a_9307_30663# a_9253_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14135 a_23763_49007# a_14831_50095# a_23669_49007# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X14136 a_7917_12265# a_7755_11471# a_7493_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14137 VSS a_29887_32375# a_18151_52263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14138 VDD a_13692_44527# a_13798_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14139 a_22632_41831# a_21663_41855# a_22536_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1414 VSS a_12591_31029# a_12120_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14140 a_19678_57174# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14141 a_46482_60186# a_16746_60188# a_46390_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14142 vcm_commonmode a_16362_16520# a_43470_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14143 a_46482_19532# a_16746_19530# a_46390_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14144 a_19678_15882# a_12877_14441# a_19282_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14145 VDD a_5211_24759# a_6743_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14146 VSS VSS a_23694_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14147 a_3339_30503# a_9529_28335# a_25462_27247# VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X14148 a_29414_70226# a_16746_70228# a_29322_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14149 a_38499_42943# a_36432_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X1415 VSS a_4903_23983# a_4571_26677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X14150 VDD a_4842_45467# a_5905_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14151 a_30418_24552# VDD a_30326_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14152 VDD VDD a_38358_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14153 VSS VDD a_34738_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14154 VDD a_3305_38671# a_7381_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14155 a_24794_68540# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14156 a_19374_62194# a_16746_62196# a_19282_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14157 VDD a_6792_43719# a_5715_44343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14158 a_10362_31171# a_4903_31849# a_10280_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14159 a_43623_27247# a_20635_29415# a_9503_26151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1416 a_34725_41831# a_35033_42044# a_34699_42035# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14160 a_9731_22895# a_9223_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14161 VDD a_8933_22583# a_10311_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X14162 a_20378_16520# a_16746_16518# a_20286_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14163 a_2840_53511# a_6743_54447# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14164 a_20351_49525# a_20195_49793# a_20496_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X14165 a_11399_18543# a_11049_18543# a_11304_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X14166 a_44778_7850# VDD a_44382_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14167 VSS a_10687_52553# a_8123_56399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X14168 a_10055_26409# a_6162_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14169 a_40762_72234# VDD a_40366_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1417 a_6007_23145# a_5085_23047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X14170 VDD a_4771_42167# a_2539_42106# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X14171 a_32730_7850# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14172 a_10200_47919# a_9392_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14173 a_28810_67536# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14174 VDD a_40737_37692# a_40343_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14175 a_25306_64202# a_11067_13095# a_25798_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14176 a_21627_49373# a_21003_49007# a_21519_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X14177 VDD a_7369_24233# a_10873_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X14178 VSS a_2411_18517# a_11017_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14179 VSS a_12546_22351# a_25702_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1418 VSS a_12967_50943# a_12901_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X14180 a_2781_15529# a_2926_15253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14181 a_36519_28879# a_28305_28879# a_36425_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X14182 a_37446_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14183 VSS a_1586_36727# a_1683_33237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14184 VDD a_10515_22671# a_22294_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14185 VSS a_10515_23975# a_28714_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14186 a_2369_26159# a_2325_26401# a_2203_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X14187 a_36350_7850# VSS a_36442_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14188 VDD a_1586_51335# a_3891_50645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14189 a_37750_70226# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1419 a_27710_21906# a_12985_7663# a_27314_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14190 a_36442_68218# a_16746_68220# a_36350_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14191 a_33668_36391# a_32795_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14192 a_35346_23914# a_16362_23548# a_35438_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14193 a_28870_51727# a_27793_51733# a_28708_52105# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14194 a_29038_50639# a_28968_50871# a_28789_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5e+11p pd=2.5e+06u as=3.85e+11p ps=2.77e+06u w=1e+06u l=150000u
X14195 a_49494_67214# a_16746_67216# a_49402_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14196 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14197 vcm_commonmode a_16362_64202# a_46482_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14198 a_48398_22910# a_16362_22544# a_48490_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14199 VDD a_24067_42583# a_23880_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X142 a_6913_72399# a_6559_72512# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1420 a_37839_47375# a_12907_27023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X14200 a_22690_12870# a_10055_58791# a_22294_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14201 a_20661_47713# a_4443_46607# a_20575_47713# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14202 a_19282_55166# VSS a_19774_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14203 a_36821_50095# a_34145_49007# a_36833_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X14204 a_7072_56053# a_7457_56053# a_7201_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X14205 VDD a_7803_55509# a_7107_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14206 a_39454_59182# a_16746_59184# a_39362_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14207 vcm_commonmode a_16362_56170# a_36442_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14208 VSS a_4685_37583# a_8656_34639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X14209 a_28817_28111# a_12907_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1421 a_22246_49373# a_21169_49007# a_22084_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14210 a_42374_71230# a_16362_71230# a_42466_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14211 a_47790_62194# a_12981_62313# a_47394_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14212 VSS a_12895_13967# a_44778_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14213 a_7721_69679# a_2686_70223# a_7637_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14214 a_41766_15882# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14215 a_20359_27791# a_15661_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14216 a_7637_53877# a_7803_55509# a_7890_54223# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X14217 a_36442_7484# VDD a_36350_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14218 VDD a_31964_30485# a_31898_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14219 a_36328_49525# a_36551_49007# a_36548_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1422 VSS a_12981_59343# a_35742_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14220 VSS a_1586_66567# a_9319_62613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14221 VDD a_11067_21583# a_32334_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14222 a_19678_10862# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14223 vcm_commonmode a_16362_9492# a_41462_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14224 a_25398_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14225 a_17216_28585# a_14471_28585# a_16961_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14226 a_22857_28111# a_17869_28585# a_22567_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14227 VSS a_12981_59343# a_17670_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14228 a_14073_28157# a_11602_25071# a_14001_28157# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14229 a_18063_31599# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1423 a_24302_12870# a_12877_16911# a_24794_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14230 a_11989_68367# a_11947_68279# a_8782_65015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14231 vcm_commonmode a_16362_9492# a_17366_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14232 a_21686_18894# a_12899_10927# a_21290_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14233 a_45782_14878# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14234 VDD a_2163_64381# a_2124_64507# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14235 VSS a_5964_35015# a_4123_37013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14236 a_36842_72556# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14237 a_28714_24918# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14238 a_32334_16886# a_12899_11471# a_32826_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14239 a_33430_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1424 a_2369_45565# a_2325_45173# a_2203_45577# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X14240 a_27406_9492# a_16746_9490# a_27314_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14241 VDD a_12901_66665# a_40366_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14242 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14243 VDD a_12981_59343# a_36350_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14244 a_49894_71552# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14245 a_12913_59049# a_11067_66191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X14246 a_16746_14510# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X14247 a_21382_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14248 a_24800_44129# a_24515_43493# a_25388_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14249 a_28881_52271# a_28423_52245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X1425 VDD a_1923_54591# a_4856_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X14250 a_20743_43493# a_19780_41605# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14251 a_19282_72234# VSS a_19374_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14252 VDD a_2223_28617# a_3957_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14253 a_17366_55166# VDD a_17274_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14254 a_18674_16886# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14255 a_49402_61190# a_16362_61190# a_49494_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14256 a_23390_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14257 VSS a_12877_14441# a_22690_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14258 vcm_commonmode a_16362_61190# a_31422_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14259 VDD a_12947_71576# a_26310_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1426 VSS a_11121_23957# a_11069_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14260 VSS a_12983_63151# a_34738_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14261 a_10660_16367# a_10543_16580# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14262 a_42709_29199# a_11067_46823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14263 a_33856_44869# a_32887_44581# a_33760_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14264 a_26402_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14265 VSS a_10975_66407# a_47790_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14266 a_8082_56775# a_7210_55081# a_8296_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=0p ps=0u w=1e+06u l=150000u
X14267 a_13287_29423# a_13239_29575# a_13180_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X14268 a_2672_40303# a_1591_40303# a_2325_40545# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X14269 a_36442_21540# a_16746_21538# a_36350_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1427 VDD a_13565_44135# a_13510_44759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14270 a_7377_60431# a_6417_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X14271 a_45878_23516# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14272 a_45478_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14273 a_75794_38962# a_75628_38962# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X14274 a_23669_49257# a_17682_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14275 a_7577_59343# a_7519_59575# a_7162_59575# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X14276 a_49494_20536# a_16746_20534# a_49402_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14277 a_24302_21906# a_16362_21540# a_24394_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14278 a_41766_56170# a_12257_56623# a_41370_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14279 a_35838_15484# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1428 VSS a_2939_52245# a_2873_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X14280 VDD a_12899_10927# a_38358_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14281 a_9865_14441# a_9275_15253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X14282 VSS a_23789_39100# a_23643_41569# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14283 VSS a_12757_8207# a_12815_6031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14284 a_2464_63517# a_2250_63517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14285 a_24698_66210# a_12983_63151# a_24302_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14286 a_3203_53686# a_2952_53333# a_2744_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14287 a_4165_22351# a_3325_18543# a_4083_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14288 a_17696_29967# a_2235_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X14289 a_39454_12504# a_16746_12502# a_39362_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1429 VSS a_25787_28327# a_33864_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.1125e+11p ps=1.95e+06u w=650000u l=150000u
X14290 VDD a_9215_58487# a_4674_57685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X14291 a_2107_9839# a_1591_9839# a_2012_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14292 VDD a_2742_42997# a_2700_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14293 a_6745_37289# a_3949_41935# a_6649_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14294 a_49494_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14295 VSS a_3391_15797# a_3023_16341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14296 a_46390_15882# a_16362_15516# a_46482_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14297 a_39362_69222# a_16362_69222# a_39454_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14298 a_43470_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14299 a_45782_55166# VSS a_45386_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X143 a_19282_62194# a_12355_15055# a_19774_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1430 a_35319_34191# a_35142_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14300 vcm_commonmode a_16362_69222# a_21382_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14301 a_36350_11866# a_10055_58791# a_36842_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14302 a_28714_65206# a_10975_66407# a_28318_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14303 VDD a_12516_7093# a_33338_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14304 a_10687_52553# a_33041_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X14305 a_27169_30083# a_25321_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14306 a_2203_26159# a_1757_26159# a_2107_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14307 VSS a_19889_27497# a_22890_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X14308 VSS a_5363_30503# a_24591_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.6875e+11p ps=4.35e+06u w=650000u l=150000u
X14309 VDD a_5791_43541# a_5778_43933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1431 VDD a_4311_58229# a_1823_65853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14310 a_5343_72221# a_4719_71855# a_5235_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14311 a_33430_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14312 a_26310_63198# a_16362_63198# a_26402_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14313 VDD a_12901_66959# a_46390_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14314 vcm_commonmode a_16362_58178# a_42466_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14315 a_16362_69222# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14316 a_18674_57174# a_10515_22671# a_18278_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14317 VDD a_7815_49855# a_7802_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14318 a_8117_30287# a_4495_35925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14319 a_8509_47673# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1432 a_46786_24918# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14320 a_15941_31375# a_14097_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14321 a_9318_32509# a_9355_32117# a_9135_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14322 vcm_commonmode a_16362_68218# a_25398_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14323 a_3066_62069# a_1591_63151# a_2985_62069# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X14324 a_34834_65528# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14325 VDD a_12877_16911# a_29322_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14326 a_1761_4399# a_1591_4399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X14327 a_7775_10625# a_1586_18695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X14328 a_44382_22910# a_10515_23975# a_44874_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14329 a_34342_55166# VSS a_34434_55166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1433 a_7741_64239# a_6515_62037# a_7439_64213# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6725e+11p ps=2.43e+06u w=650000u l=150000u
X14330 a_47886_64524# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14331 VDD a_31131_35281# a_30991_35307# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14332 a_42165_36367# a_41999_36367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X14333 VSS a_12981_62313# a_23694_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14334 a_20682_60186# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14335 a_20682_19898# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14336 VDD a_22132_44129# a_25204_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X14337 a_33430_71230# a_16746_71232# a_33338_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14338 a_5265_18543# a_4075_18543# a_5156_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X14339 VSS a_37706_44135# a_37711_43983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1434 a_17670_13874# a_12877_16911# a_17274_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14340 vcm_commonmode a_16362_59182# a_28410_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14341 a_37750_23914# a_10515_23975# a_37354_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14342 a_34342_14878# a_12877_14441# a_34834_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14343 VSS a_12985_7663# a_34738_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14344 a_32426_57174# a_16746_57176# a_32334_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14345 a_33734_18894# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14346 a_37846_56492# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14347 a_17274_24918# VSS a_17766_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14348 a_7910_38671# a_6372_38279# a_7838_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14349 a_48794_9858# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1435 a_35224_49871# a_28881_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.85e+11p pd=5.37e+06u as=0p ps=0u w=1e+06u l=150000u
X14350 a_21782_22512# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14351 a_23734_29941# a_7939_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14352 VDD a_12355_65103# a_24302_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14353 a_48398_60186# a_12727_58255# a_48890_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14354 a_6917_31055# a_6372_38279# a_6835_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14355 VSS a_13692_34191# a_13798_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14356 VSS a_17280_48695# a_17095_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14357 VSS a_29513_42333# a_29205_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14358 VSS a_3509_58487# a_2695_58951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14359 a_12806_13967# a_11067_63143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1436 vcm_commonmode VSS a_24394_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14360 a_11714_14557# a_10995_14333# a_11151_14428# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14361 VDD a_13909_39747# a_39141_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X14362 a_25306_72234# VDD a_25798_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14363 VSS a_3173_53333# a_3107_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14364 a_36746_70226# a_12901_66665# a_36350_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14365 a_21021_46805# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14366 VSS a_7749_55535# a_8496_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14367 a_22294_14878# a_16362_14512# a_22386_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14368 a_5594_36727# a_3305_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14369 a_7467_57863# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1437 VSS a_14425_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X14370 a_8937_18319# a_7377_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14371 a_25798_60508# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14372 VDD a_23901_44220# a_23507_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14373 a_30557_49783# a_30762_49641# a_30720_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14374 a_33730_47375# a_19807_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14375 a_3166_70589# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14376 vcm_commonmode a_16362_17524# a_37446_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14377 VDD a_27247_43047# a_24893_37429# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X14378 a_15315_27791# a_15064_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X14379 VDD a_10509_73193# a_10865_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1438 a_33668_38567# a_33764_38567# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X14380 a_41462_15516# a_16746_15514# a_41370_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14381 VDD a_24800_44129# a_23901_44220# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X14382 a_7335_18038# a_7153_18038# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14383 a_35742_9858# a_12985_19087# a_35346_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14384 vcm_commonmode a_16362_22544# a_21382_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14385 VDD a_18602_55312# a_18278_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14386 VSS a_15607_46805# a_40691_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14387 a_24423_40229# a_23415_41263# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14388 VDD a_11999_67477# a_11803_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14389 a_39758_61190# a_12355_15055# a_39362_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1439 a_2834_69135# a_1757_69141# a_2672_69513# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14390 a_28810_12472# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14391 a_10480_67075# a_10379_66389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14392 a_40762_57174# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14393 a_15489_50639# a_13445_50639# a_15074_50871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14394 vcm_commonmode VSS a_46482_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14395 VSS a_7461_27247# a_9307_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14396 a_2040_17289# a_1591_16917# a_1945_16911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X14397 a_2672_12937# a_1757_12565# a_2325_12533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14398 a_23694_67214# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14399 a_30722_68218# a_12901_66959# a_30326_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X144 a_26112_30663# a_14926_31849# a_26343_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1440 a_37354_72234# VSS a_37446_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14400 vcm_commonmode a_16362_11500# a_42466_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14401 VDD a_2235_30503# a_15941_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14402 a_18674_10862# a_12546_22351# a_18278_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14403 VDD a_3325_18543# a_4333_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14404 a_22351_47893# a_22176_47919# a_22530_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14405 a_41862_19500# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14406 vcm_commonmode a_16362_21540# a_25398_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14407 a_28410_24552# VDD a_28318_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14408 VSS a_2292_43291# a_5957_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14409 a_40458_62194# a_16746_62196# a_40366_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1441 VSS a_12727_58255# a_39758_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14410 VDD a_6619_16341# a_6606_16733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14411 VSS a_13357_32143# a_22148_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14412 a_44778_14878# a_12727_15529# a_44382_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14413 a_5515_60137# a_5653_60039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14414 a_23790_63520# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14415 a_3957_28995# a_2216_28309# a_3885_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14416 a_44382_7850# VSS a_44474_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14417 VSS a_12947_56817# a_30722_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14418 a_18370_16520# a_16746_16518# a_18278_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14419 a_27504_36165# a_26631_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X1442 VSS a_11067_67279# a_39758_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14420 VSS a_35493_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X14421 a_27806_18496# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14422 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14423 VDD a_12727_13353# a_31330_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14424 a_45386_69222# a_12901_66959# a_45878_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14425 vcm_commonmode a_16362_12504# a_28410_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14426 a_14273_27791# a_13919_27904# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14427 a_32426_10496# a_16746_10494# a_32334_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14428 VSS a_17763_35797# a_17585_37477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14429 a_17670_58178# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1443 a_42224_42693# a_41351_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X14430 a_5825_20495# a_3987_19623# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X14431 a_41351_42405# a_40585_42369# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14432 VSS a_1586_45431# a_6559_45205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14433 a_33430_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14434 a_32334_67214# a_16362_67214# a_32426_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14435 a_5906_28585# a_5449_25071# a_5906_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14436 a_2215_10205# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14437 a_30746_28335# a_28757_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14438 VDD a_12947_8725# a_18278_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14439 a_46482_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1444 a_35438_55166# VDD a_35346_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14440 a_22786_69544# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14441 VSS a_9314_69367# a_10699_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14442 a_17366_63198# a_16746_63200# a_17274_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14443 a_30326_8854# a_12985_19087# a_30818_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14444 a_13155_28111# a_11902_27497# a_12965_27791# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X14445 a_22294_59182# a_16362_59182# a_22386_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14446 a_35345_28879# a_28305_28879# a_35263_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14447 a_24698_8854# a_12947_8725# a_24302_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14448 a_42770_17890# a_12899_11471# a_42374_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14449 VSS a_30928_49007# a_36328_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1445 a_36746_16886# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14450 a_35069_51433# a_28881_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14451 VSS a_38315_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X14452 a_40366_55166# VSS a_40858_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14453 a_49798_23914# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14454 VDD a_7255_10357# a_7203_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14455 a_23298_65206# a_12355_65103# a_23790_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14456 a_7001_51433# a_6795_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14457 a_5136_34551# a_4495_35925# a_5367_34435# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14458 a_37039_36919# a_36107_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14459 a_39758_15882# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1446 a_41462_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14460 a_9363_65327# a_2840_66103# a_9280_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X14461 VSS a_8453_51727# a_10426_51549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14462 vcm_commonmode a_16362_71230# a_22386_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14463 VSS a_12727_15529# a_43774_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14464 VDD a_13005_35823# a_12641_37684# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14465 a_40762_10862# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14466 a_2083_74913# a_1586_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14467 VDD a_24959_30503# a_32779_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14468 VSS a_12947_23413# a_26706_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14469 a_23694_20902# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1447 a_6327_72917# a_6453_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14470 a_27183_43493# a_23567_43123# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X14471 a_2361_74575# a_2083_74913# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X14472 a_24714_32259# a_22399_32143# a_24632_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14473 a_30722_21906# a_12985_7663# a_30326_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14474 a_30835_39783# a_28099_42895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14475 a_26310_56170# a_12947_56817# a_26802_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14476 a_35438_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14477 a_10969_59663# a_2840_66103# a_10751_59575# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14478 a_18053_28879# a_16101_31029# a_18053_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14479 a_48794_70226# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1448 VSS a_12877_14441# a_40762_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14480 a_47486_68218# a_16746_68220# a_47394_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14481 VDD a_5607_44343# a_5043_44085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X14482 a_2672_12937# a_1591_12565# a_2325_12533# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14483 a_46390_23914# a_16362_23548# a_46482_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14484 a_20682_13874# a_12877_16911# a_20286_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14485 VSS a_20715_34717# a_20655_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14486 a_40458_8488# a_16746_8486# a_40366_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14487 a_8671_22671# a_5531_22895# a_8583_22671# VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=0p ps=0u w=650000u l=150000u
X14488 VDD a_13743_35836# a_19684_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X14489 a_23172_31573# a_5915_35943# a_23392_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1449 a_7389_22467# a_6816_19355# a_7294_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X14490 a_38754_62194# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14491 a_28295_31287# a_28618_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14492 a_2215_45021# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14493 a_40366_72234# VSS a_40458_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14494 a_45782_63198# a_15439_49525# a_45386_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14495 VSS a_12727_58255# a_42770_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14496 a_16043_38825# a_15683_39141# a_16556_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14497 a_20359_29199# a_40691_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14498 VSS a_11067_67279# a_42770_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14499 a_17507_30761# a_17554_30663# a_17943_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 a_6599_40630# a_6417_40630# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1450 VDD a_7598_36103# a_7215_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14500 VDD a_11121_23957# a_11069_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14501 VDD a_31171_27412# a_29760_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X14502 a_32730_66210# a_12983_63151# a_32334_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14503 VSS a_1586_36727# a_4259_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14504 VSS a_12516_7093# a_25702_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14505 a_2012_66415# a_1895_66628# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14506 a_17274_58178# a_10515_22671# a_17766_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14507 a_12283_42359# a_12677_42333# a_12343_42333# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X14508 a_13291_37999# a_13111_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14509 a_17670_11866# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1451 VSS a_5795_27497# a_6216_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X14510 vcm_commonmode a_16362_61190# a_29414_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14511 a_39854_24520# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14512 VDD a_11067_21583# a_43378_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14513 vcm_commonmode a_16362_15516# a_30418_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14514 VDD a_30415_50871# a_28968_50871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14515 VDD a_18197_36604# a_17803_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14516 VDD a_2011_34837# a_4762_35484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14517 a_6793_73825# a_5441_72399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14518 a_30418_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14519 VDD a_12727_15529# a_33338_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1452 a_36612_39655# a_36708_39655# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X14520 a_6835_46823# a_8643_48767# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14521 VDD VSS a_16270_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14522 a_34342_63198# a_16362_63198# a_34434_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14523 a_47886_72556# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14524 VDD a_39176_44527# a_39282_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14525 a_16385_51183# a_16219_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X14526 a_11801_64015# a_11759_63927# a_9735_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X14527 VDD a_12985_7663# a_47394_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14528 VSS a_1586_21959# a_3983_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14529 a_44474_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1453 a_2451_72373# a_4119_70741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X14530 a_41370_11866# a_16362_11500# a_41462_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14531 a_47394_62194# a_16362_62194# a_47486_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14532 a_30326_19898# a_11067_67279# a_30818_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14533 VDD a_13349_37973# a_13291_37999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14534 a_4161_25321# a_2223_28617# a_4065_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14535 VDD a_2419_48783# a_2511_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X14536 VDD a_12877_16911# a_37354_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14537 a_34834_10464# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14538 a_4903_31849# a_4702_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14539 VSS a_35932_38689# a_36579_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X1454 a_23298_18894# a_12895_13967# a_23790_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14540 a_17766_20504# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14541 VDD VDD a_24302_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14542 a_17366_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14543 VDD a_1586_66567# a_9135_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14544 a_48490_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14545 a_8643_48767# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14546 a_24394_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14547 VDD a_1952_60431# a_2727_56417# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14548 a_75445_39738# a_75541_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14549 VSS a_12983_63151# a_45782_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1455 VDD a_1586_9991# a_5639_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14550 a_7628_18365# a_7377_18012# a_7407_18038# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X14551 vcm_commonmode a_16362_69222# a_19374_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14552 a_23390_67214# a_16746_67216# a_23298_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14553 vcm_commonmode a_16362_64202# a_20378_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14554 VDD a_25015_48437# a_26187_48801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14555 a_12621_62313# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14556 a_47486_21540# a_16746_21538# a_47394_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14557 a_22294_22910# a_16362_22544# a_22386_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14558 VSS a_12901_58799# a_35742_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14559 VDD a_12355_65103# a_32334_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1456 a_4864_62581# a_2689_65103# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14560 a_2464_56989# a_2250_56989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14561 a_18278_12870# a_16362_12504# a_18370_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14562 a_3983_12879# a_1929_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X14563 a_21479_36965# a_20713_36929# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14564 a_14941_51183# a_13925_51727# a_14859_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14565 a_24331_40767# a_22632_41831# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14566 a_29269_40741# a_29943_41317# a_30816_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14567 VDD a_15439_49525# a_45386_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14568 a_37655_49667# a_35676_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14569 a_15315_52271# a_15285_52245# a_8132_53511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X1457 VSS a_3023_16341# a_3523_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X14570 a_37446_13508# a_16746_13506# a_37354_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14571 VDD a_12899_10927# a_49402_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14572 VDD a_2746_16885# a_2704_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14573 a_7563_46261# a_7368_46403# a_7873_46653# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X14574 VDD a_2939_31573# a_2926_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14575 VDD a_17449_46831# a_18243_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X14576 VSS a_2744_53511# a_2007_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14577 a_32795_36415# a_31280_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X14578 a_25798_9460# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14579 VSS a_12899_10927# a_31726_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1458 vcm_commonmode a_16362_15516# a_27406_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14580 VDD a_16244_34973# a_15345_34717# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X14581 VSS a_10515_22671# a_39758_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14582 a_33830_60508# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14583 a_36746_55166# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14584 a_3026_23805# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14585 VDD a_11865_24527# a_11574_22869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X14586 a_41462_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14587 a_11035_47893# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14588 a_2840_66103# a_34895_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14589 a_2560_45895# a_2539_42106# a_2702_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1459 VDD a_33593_31287# a_32367_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X14590 a_36395_44265# a_35463_44031# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14591 VDD a_30267_35253# a_30091_35253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14592 VDD a_2764_33609# a_2939_33535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14593 VDD a_12516_7093# a_44382_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14594 a_2787_32679# a_6655_46261# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14595 a_32730_13874# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14596 VDD a_35969_28111# a_36459_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X14597 VDD a_2411_18517# a_10475_14165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14598 a_23790_71552# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14599 a_44474_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X146 VSS a_10515_22671# a_29718_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1460 a_3668_10749# a_3417_10927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X14600 a_41370_56170# a_16362_56170# a_41462_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14601 a_19774_61512# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14602 a_37750_8854# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14603 VDD a_17358_31069# a_17507_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X14604 a_77002_40202# a_77098_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14605 a_17787_47349# a_18222_47507# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X14606 a_27406_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14607 a_29718_57174# a_10515_22671# a_29322_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14608 a_44778_66210# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14609 VDD a_7565_31751# a_7571_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1461 VDD a_12947_71576# a_44382_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14610 VDD a_4187_60673# a_4148_60547# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14611 a_42374_23914# a_12947_23413# a_42866_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14612 a_11067_66191# a_11067_46823# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X14613 a_6559_59879# a_19502_51157# a_19446_51183# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14614 a_42374_19898# a_16362_19532# a_42466_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14615 VSS a_12985_19087# a_47790_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14616 VSS a_5381_68345# a_5315_68413# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14617 a_45878_65528# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14618 a_12277_39429# a_12585_39069# a_12251_39069# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X14619 a_7573_60431# a_6559_59879# a_7449_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X1462 a_31422_13508# a_16746_13506# a_31330_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14620 a_48490_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14621 a_45386_55166# VSS a_45478_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14622 a_2592_43023# a_1757_43029# a_2620_43389# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14623 a_5297_58621# a_4918_58255# a_5225_58621# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X14624 a_35742_24918# VSS a_35346_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14625 a_31726_60186# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14626 VSS a_9305_53511# a_7764_53877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14627 a_44474_71230# a_16746_71232# a_44382_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14628 a_30418_58178# a_16746_58180# a_30326_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14629 a_31726_19898# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1463 VDD a_4674_40277# a_5074_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X14630 VSS a_10975_66407# a_21686_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14631 VDD a_22521_37692# a_22127_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14632 a_35838_57496# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14633 a_12712_59343# a_11067_13095# a_12539_59663# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14634 a_48890_17492# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14635 a_45386_14878# a_12877_14441# a_45878_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14636 VSS a_12985_7663# a_45782_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14637 a_48794_23914# a_10515_23975# a_48398_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14638 a_28011_41855# a_27245_41829# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14639 VDD a_11902_27497# a_13919_27904# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X1464 a_8836_74953# a_7921_74581# a_8489_74549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X14640 vcm_commonmode a_16362_22544# a_19374_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14641 a_28318_24918# VSS a_28810_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14642 a_23390_20536# a_16746_20534# a_23298_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14643 a_1846_57963# a_2124_57979# a_2080_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14644 a_18278_57174# a_16362_57174# a_18370_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14645 a_32826_22512# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14646 a_22386_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14647 a_4775_32687# a_4425_32687# a_4680_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X14648 a_38754_15882# a_12877_14441# a_38358_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14649 VSS a_12877_16911# a_35742_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1465 a_24768_27247# a_2235_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X14650 VSS a_17787_47349# a_3339_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X14651 a_48490_70226# a_16746_70228# a_48398_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14652 a_12218_55901# a_11141_55535# a_12056_55535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14653 VDD a_12899_11471# a_25306_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14654 a_8029_13353# a_7999_13083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14655 a_6816_19355# a_8827_17215# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X14656 a_22786_14480# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14657 a_49402_13874# a_12727_15529# a_49894_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14658 VSS a_9557_64757# a_8896_65015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14659 a_9187_10901# a_2004_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X1466 a_2882_58077# a_2124_57979# a_2319_57948# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X14660 a_20286_15882# a_16362_15516# a_20378_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14661 a_23390_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14662 a_43870_68540# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14663 a_38450_62194# a_16746_62196# a_38358_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14664 a_6444_16367# a_5529_16367# a_6097_16609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14665 VDD a_35815_31751# a_41243_30080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X14666 a_32310_49257# a_17682_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14667 a_39854_58500# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14668 vcm_commonmode a_16362_18528# a_35438_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14669 VSS a_6598_69653# a_6373_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X1467 a_44474_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14670 a_33338_14878# a_16362_14512# a_33430_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14671 VSS a_10055_58791# a_39758_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14672 a_28602_52271# a_2872_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14673 a_6614_21237# a_5671_21495# a_7170_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14674 vcm_commonmode a_16362_17524# a_48490_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14675 VSS a_12947_56817# a_28714_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14676 vcm_commonmode a_16362_8488# a_39454_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14677 a_26802_13476# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14678 a_23298_10862# a_12985_16367# a_23790_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14679 a_26706_7850# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1468 VDD a_2672_44655# a_2847_44629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14680 a_7737_74031# a_6224_73095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14681 VDD a_12985_16367# a_30326_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14682 VSS a_34759_31029# a_37589_31393# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14683 VDD VSS a_29322_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14684 VDD a_12901_66959# a_20286_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14685 a_21686_68218# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14686 a_44382_64202# a_11067_13095# a_44874_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14687 a_49494_8488# a_16746_8486# a_49402_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14688 a_5134_50639# a_4057_50645# a_4972_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14689 VDD a_28446_31375# a_38299_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1469 a_2557_72943# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14690 a_33756_31171# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14691 a_30939_31055# a_20635_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14692 VDD a_7959_15279# a_8361_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14693 a_4330_63827# a_4608_63811# a_4564_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14694 a_25398_17524# a_16746_17522# a_25306_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14695 a_30190_32143# a_30155_32375# a_29887_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14696 a_23599_38007# a_23993_37981# a_23565_38565# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X14697 VSS a_33856_40743# a_33819_41001# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X14698 a_8121_48437# a_7903_48841# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14699 a_34342_56170# a_12947_56817# a_34834_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X147 a_23790_60508# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1470 a_27406_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14700 a_29718_10862# a_12546_22351# a_29322_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14701 a_36350_70226# a_16362_70226# a_36442_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14702 a_3143_66972# a_4220_68021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14703 VDD a_20635_29415# a_31117_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14704 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14705 a_17274_66210# a_10975_66407# a_17766_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14706 VDD a_4333_22895# a_4903_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X14707 a_21782_64524# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14708 a_24302_8854# a_16362_8488# a_24394_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14709 VSS a_24683_48463# a_24673_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1471 a_29718_18894# a_12899_10927# a_29322_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14710 a_3307_18259# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14711 a_29414_16520# a_16746_16518# a_29322_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14712 vcm_commonmode a_16362_13508# a_26402_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14713 VDD a_11067_67279# a_39362_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14714 VDD a_2325_40545# a_2215_40669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14715 a_30418_11500# a_16746_11498# a_30326_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14716 VSS a_12516_7093# a_33734_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14717 a_12445_50613# a_12227_51017# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14718 VDD a_24800_43041# a_23901_43132# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X14719 a_28714_58178# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1472 a_30722_55166# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14720 a_22294_60186# a_12727_58255# a_22786_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14721 vcm_commonmode a_16362_66210# a_38450_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14722 a_28305_28879# a_28027_29217# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14723 a_13835_41001# a_13107_41317# a_13980_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14724 a_17429_32509# a_17394_32275# a_17191_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14725 a_30326_68218# a_16362_68218# a_30418_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14726 a_42466_64202# a_16746_64204# a_42374_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14727 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14728 a_13111_37999# a_13123_38231# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14729 a_2250_63517# a_2163_63293# a_1846_63403# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1473 a_31481_28585# a_30052_32117# a_30975_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14730 a_44474_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14731 a_2985_62069# a_1952_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14732 a_7841_29673# a_6649_25615# a_7841_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14733 VSS a_4191_33449# a_16587_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14734 a_33764_41831# a_32795_41855# a_33727_42089# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X14735 VSS a_12981_59343# a_36746_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14736 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14737 VDD a_2319_54684# a_2250_54813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14738 VDD config_2_in[3] a_1591_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X14739 vcm_commonmode VSS a_28410_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1474 a_43470_66210# a_16746_66212# a_43378_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14740 VSS a_1923_73087# a_2369_71677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14741 a_40762_18894# a_12899_10927# a_40366_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14742 VSS a_12901_66665# a_19678_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14743 a_33338_59182# a_16362_59182# a_33430_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14744 a_12394_25615# a_11430_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X14745 a_17366_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14746 a_47790_24918# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14747 VSS a_21479_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X14748 VSS a_9240_53877# a_9305_53511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14749 a_10615_72399# a_10509_73193# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1475 a_22530_47919# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X14750 a_6829_15279# a_5639_15279# a_6720_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X14751 VDD a_2284_36103# a_1591_36103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14752 VSS a_2847_23743# a_2781_23817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X14753 a_27333_32143# a_5363_30503# a_27417_32509# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X14754 VDD a_14735_35805# a_14761_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X14755 VDD a_7833_66415# a_8307_66415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14756 a_31741_30485# a_31659_31751# a_31898_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X14757 a_48398_9858# a_12546_22351# a_48890_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14758 a_36442_55166# VDD a_36350_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14759 a_37750_16886# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1476 VSS a_11803_55311# a_16746_58180# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X14760 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14761 a_28680_30057# a_28670_30663# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14762 vcm_commonmode VSS a_20378_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14763 a_18539_47617# a_4191_33449# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14764 VSS a_12877_14441# a_41766_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14765 a_35346_10862# a_16362_10496# a_35438_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14766 a_19374_65206# a_16746_65208# a_19282_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14767 VDD VDD a_32334_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14768 a_24302_18894# a_12895_13967# a_24794_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14769 a_21686_21906# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1477 a_27779_52271# a_27333_52271# a_27683_52271# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X14770 VSS VSS a_24698_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14771 a_18278_20902# a_16362_20536# a_18370_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14772 a_36904_28879# a_36425_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X14773 vcm_commonmode a_16362_71230# a_33430_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14774 VDD a_5381_68345# a_5411_68086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14775 VSS a_37733_37477# a_39247_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X14776 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X14777 VDD a_12947_71576# a_45386_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14778 a_17670_60186# a_12981_59343# a_17274_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14779 a_17670_19898# a_12895_13967# a_17274_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1478 a_33681_49373# a_32856_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.297e+11p pd=3.25e+06u as=0p ps=0u w=420000u l=150000u
X14780 a_38867_38591# a_38101_38565# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X14781 a_7567_64391# a_7445_63695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14782 VSS a_4528_26159# a_7571_22057# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14783 a_20378_9492# a_16746_9490# a_20286_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14784 a_7293_49525# a_7075_49929# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14785 a_28410_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14786 VSS a_12727_13353# a_27710_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14787 a_11968_28585# a_9179_22351# a_11747_28639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X14788 a_36746_63198# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14789 VSS a_21856_36513# a_22595_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X1479 a_19492_52245# a_19877_52245# a_19621_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X14790 a_31726_13874# a_12877_16911# a_31330_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14791 VSS a_2411_19605# a_4853_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14792 VSS a_4211_67655# a_1954_61677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X14793 VSS a_2944_57960# a_2882_58077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X14794 a_26319_35253# a_26495_35253# a_26447_35279# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X14795 a_9865_68047# a_3024_67191# a_8772_63927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X14796 a_39362_11866# a_16362_11500# a_39454_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14797 VSS a_1689_10396# a_1633_10422# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14798 VDD a_12985_19087# a_35346_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14799 VDD a_4528_26159# a_5337_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X148 a_26706_55166# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1480 VDD a_4864_62581# a_3016_60949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X14800 VSS a_19877_52245# a_19492_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14801 a_32334_68218# a_12727_67753# a_32826_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14802 a_43774_66210# a_12983_63151# a_43378_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14803 a_2603_64783# a_1768_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X14804 vcm_commonmode a_16362_62194# a_27406_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14805 a_28318_58178# a_10515_22671# a_28810_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14806 a_11067_67279# a_9989_46831# a_11297_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X14807 a_31422_60186# a_16746_60188# a_31330_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14808 VSS a_1775_60663# a_2300_61879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14809 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1481 a_42374_21906# a_16362_21540# a_42466_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14810 a_31422_19532# a_16746_19530# a_31330_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14811 VDD a_10515_23975# a_41370_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14812 a_28714_11866# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14813 a_29361_51727# a_28883_52031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X14814 a_41370_64202# a_16362_64202# a_41462_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14815 VSS a_4495_35925# a_8662_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X14816 VDD a_3016_60949# a_7009_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14817 a_9280_65327# a_9513_65301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14818 a_3137_16367# a_2283_15797# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14819 a_16362_11500# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X1482 a_1757_36501# a_1591_36501# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14820 VDD a_3325_49551# a_4181_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14821 vcm_commonmode a_16362_69222# a_40458_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14822 a_47790_65206# a_10975_66407# a_47394_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14823 a_38358_21906# a_11067_21583# a_38850_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14824 a_28063_32193# a_27387_32373# a_27890_32459# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.8025e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=150000u
X14825 a_8015_20175# a_7571_20291# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X14826 a_38358_17890# a_16362_17524# a_38450_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14827 VDD a_12727_15529# a_44382_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14828 a_42466_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14829 a_12709_20969# a_4792_20443# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1483 VDD a_33856_42693# a_33760_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X14830 a_45386_63198# a_16362_63198# a_45478_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14831 a_11400_26133# a_7571_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X14832 VSS a_2872_44111# a_28405_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14833 a_28113_29217# a_25269_27791# a_28027_29217# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X14834 a_37750_57174# a_10515_22671# a_37354_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14835 VSS a_5271_17999# a_5363_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14836 VSS a_28423_52245# a_28357_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14837 vcm_commonmode a_16362_68218# a_44474_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14838 VSS a_11067_13095# a_17670_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14839 a_2764_31599# a_1849_31599# a_2417_31841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1484 VDD a_12901_66665# a_48398_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14840 VDD a_8531_70543# a_35683_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14841 a_7271_53135# a_7217_53047# a_7175_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14842 a_1757_44655# a_1591_44655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14843 VSS a_8082_54599# a_7313_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14844 VDD a_12877_16911# a_48398_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14845 a_42188_43677# a_41351_42405# a_42283_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X14846 a_7615_73193# a_6453_71855# a_7257_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X14847 a_45878_10464# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14848 a_18278_65206# a_16362_65206# a_18370_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14849 VSS a_19626_31751# a_32544_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1485 a_38358_11866# a_16362_11500# a_38450_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14850 a_28688_50247# a_29147_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14851 VSS a_2686_70223# a_7063_70313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14852 a_2325_66657# a_2107_66415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X14853 a_22386_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14854 VDD a_9405_31599# a_10701_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X14855 a_19374_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14856 VSS a_11067_66191# a_12565_8545# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14857 a_22690_70226# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14858 a_21382_68218# a_16746_68220# a_21290_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14859 vcm_commonmode a_16362_59182# a_47486_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1486 VDD a_12985_19087# a_25306_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X14860 a_35602_34191# a_35425_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14861 a_8389_32937# a_6883_37019# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14862 a_7865_46805# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14863 a_20286_23914# a_16362_23548# a_20378_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14864 vcm_commonmode a_16362_64202# a_31422_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14865 a_39854_66532# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14866 a_36350_63198# a_12981_62313# a_36842_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14867 a_33338_22910# a_16362_22544# a_33430_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14868 VSS a_17191_32117# a_16917_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14869 VDD a_12355_65103# a_43378_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1487 VDD a_6260_10927# a_6435_10901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14870 a_40858_61512# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14871 VDD a_1586_21959# a_3983_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X14872 a_35438_14512# a_16746_14510# a_35346_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14873 a_39362_56170# a_16362_56170# a_39454_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14874 a_25702_61190# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14875 a_24394_59182# a_16746_59184# a_24302_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14876 vcm_commonmode a_16362_56170# a_21382_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14877 VDD a_2672_30345# a_2847_30271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14878 a_15548_30761# a_10531_31055# a_15986_30511# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X14879 a_10430_52854# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1488 a_5709_15055# a_4629_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X14880 VDD a_12257_56623# a_33338_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14881 a_2672_40303# a_1757_40303# a_2325_40545# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14882 a_44382_72234# VDD a_44874_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14883 a_11053_69135# a_10575_69439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14884 a_12202_54599# a_12231_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14885 a_44874_60508# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14886 VDD a_6224_73095# a_6559_72512# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14887 a_16362_56170# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X14888 VSS VDD a_36746_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14889 a_29718_60186# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1489 a_27314_19898# a_11067_67279# a_27806_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14890 a_28410_58178# a_16746_58180# a_28318_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14891 a_29718_19898# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14892 vcm_commonmode VSS a_25398_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14893 a_15193_42917# a_15775_42405# a_16707_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X14894 a_41766_9858# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14895 a_30722_14878# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14896 a_46786_7850# VDD a_46390_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14897 vcm_commonmode a_16362_22544# a_40458_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14898 VDD VSS a_37354_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14899 a_7071_62581# a_7199_62839# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=2.43e+06u as=0p ps=0u w=650000u l=150000u
X149 a_39454_66210# a_16746_66212# a_39362_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1490 a_31330_68218# a_12727_67753# a_31822_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X14900 a_29072_38567# a_28103_38591# a_28976_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14901 a_21782_72556# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14902 a_5823_28585# a_5449_25071# a_5906_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14903 a_17766_62516# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14904 a_17670_9858# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14905 a_6666_53609# a_3668_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14906 VDD a_12981_59343# a_21290_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14907 a_19442_28585# a_17278_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X14908 a_42770_67214# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14909 a_33430_17524# a_16746_17522# a_33338_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1491 a_48490_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14910 a_26576_50095# a_6559_59663# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X14911 a_10595_30511# a_9307_30663# a_10423_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X14912 a_3025_64783# a_1770_14441# a_2603_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X14913 a_37750_10862# a_12546_22351# a_37354_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14914 VSS a_12546_22351# a_27710_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14915 a_4266_64566# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X14916 vcm_commonmode a_16362_21540# a_44474_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14917 a_5795_27497# a_3972_25615# a_5723_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14918 a_12950_30511# a_11812_30511# a_12631_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14919 VSS a_41820_41501# a_42375_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X1492 vcm_commonmode a_16362_62194# a_26402_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14920 a_16824_28309# a_11902_27497# a_17044_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14921 VSS a_9653_69831# a_9466_69653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14922 a_42466_72234# VDD a_42374_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14923 a_38358_7850# VSS a_38450_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14924 a_33856_40743# a_32887_40767# a_33760_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X14925 vcm_commonmode a_16362_13508# a_34434_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14926 a_40176_28335# a_15607_46805# a_40086_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X14927 VSS a_8902_36469# a_8543_36469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14928 a_46882_18496# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14929 a_46786_24918# VSS a_46390_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1493 VSS a_12677_40157# a_12369_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X14930 a_43378_15882# a_12727_13353# a_43870_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14931 VDD a_2325_12533# a_2215_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14932 VDD a_16101_31029# a_18551_29451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14933 VDD a_6095_44807# a_11157_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14934 VSS a_10975_66407# a_32730_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14935 vcm_commonmode a_16362_23548# a_17366_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14936 a_8275_43255# a_4443_46607# a_8449_43361# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X14937 vcm_commonmode a_16362_12504# a_47486_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14938 a_21382_21540# a_16746_21538# a_21290_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14939 a_2012_15101# a_1895_14906# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1494 VDD a_11803_64239# a_11759_63927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14940 a_30818_23516# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14941 a_4761_48829# a_4717_48437# a_4595_48841# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X14942 a_30418_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14943 a_33135_28335# a_20635_29415# a_32772_7638# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X14944 a_24515_34789# a_20623_36595# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X14945 a_11764_65845# a_11659_66567# a_11893_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X14946 a_36746_16886# a_12727_13353# a_36350_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14947 a_6435_74005# a_6260_74031# a_6614_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X14948 a_19678_68218# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14949 a_29361_38017# a_28747_37503# a_29620_37479# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1495 a_30418_60186# a_16746_60188# a_30326_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14950 VSS a_38784_42589# a_39431_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X14951 a_49798_57174# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14952 a_9970_56118# a_5682_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X14953 a_5169_23145# a_5085_23047# a_5087_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X14954 a_49798_15882# a_12877_14441# a_49402_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X14955 a_20778_15484# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14956 VDD a_12899_10927# a_23298_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14957 a_38450_7484# VDD a_38358_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14958 VDD a_1761_52815# a_30591_37455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14959 VDD a_2686_70223# a_5245_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1496 a_30418_19532# a_16746_19530# a_30326_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14960 VDD a_10901_52245# a_10931_52598# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X14961 a_41862_69544# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14962 a_24394_12504# a_16746_12502# a_24302_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14963 a_36613_48169# a_22843_29415# a_36459_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X14964 a_36442_63198# a_16746_63200# a_36350_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14965 VDD a_5039_42167# a_14830_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14966 vcm_commonmode a_16362_9492# a_43470_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14967 a_37846_59504# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14968 a_31330_15882# a_16362_15516# a_31422_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14969 a_2177_53359# a_1899_53387# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X1497 VSS a_2473_34293# a_3803_35523# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14970 a_17003_49770# a_17095_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X14971 a_49494_62194# a_16746_62196# a_49402_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14972 result_out[6] a_1644_62581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X14973 vcm_commonmode a_16362_18528# a_46482_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14974 a_24302_69222# a_16362_69222# a_24394_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X14975 VSS a_12257_56623# a_26706_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14976 vcm_commonmode a_16362_9492# a_19374_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14977 a_30722_55166# VSS a_30326_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14978 a_5484_69455# a_5682_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14979 a_21290_11866# a_10055_58791# a_21782_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1498 a_13059_27791# a_12631_28585# a_12965_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X14980 a_8087_17289# a_7737_16917# a_7992_17277# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X14981 VDD a_19478_51959# a_19621_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14982 a_19525_51017# a_18335_50645# a_19416_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X14983 a_33819_44535# a_32887_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14984 a_29414_9492# a_16746_9490# a_29322_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X14985 a_17033_38565# a_16879_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14986 a_42374_65206# a_12355_65103# a_42866_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14987 a_28410_11500# a_16746_11498# a_28318_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14988 a_1823_54973# a_2847_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14989 VDD a_6435_10901# a_6422_11293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1499 VSS a_40783_46831# a_15607_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X14990 a_5550_52637# a_4831_52413# a_4987_52508# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X14991 VDD a_12895_13967# a_27314_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14992 a_16154_41807# a_15459_41781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X14993 VSS a_12189_46805# a_12123_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14994 a_23390_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14995 VDD a_12901_66959# a_31330_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X14996 a_9556_67503# a_8772_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X14997 a_5340_32687# a_4259_32687# a_4993_32929# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X14998 a_42770_20902# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14999 VDD a_5064_20719# a_5239_20693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15 a_25398_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X150 a_4429_14191# a_4075_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1500 a_7640_49929# a_6725_49557# a_7293_49525# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X15000 a_39468_37479# a_38499_37503# a_39372_37479# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X15001 a_45386_56170# a_12947_56817# a_45878_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15002 VDD a_24800_41953# a_25204_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15003 VSS a_12901_66665# a_40762_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15004 a_4266_64239# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15005 a_28318_66210# a_10975_66407# a_28810_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15006 VSS a_1761_30511# a_32971_35281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X15007 a_23141_52521# a_23193_52245# a_6775_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15008 a_39758_64202# a_12355_65103# a_39362_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15009 a_32826_64524# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1501 a_7758_65693# a_7039_65469# a_7195_65564# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X15010 VSS a_5039_42167# a_15483_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15011 a_22690_23914# a_10515_23975# a_22294_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15012 a_12953_53339# a_12631_52928# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15013 VSS a_8485_71855# a_9782_71311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15014 a_22786_56492# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15015 a_49402_55166# VSS a_49894_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15016 vcm_commonmode a_16362_67214# a_36442_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15017 a_11771_68021# a_11053_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15018 a_2250_56989# a_2163_56765# a_1846_56875# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15019 VSS a_12516_7093# a_44778_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1502 a_77568_39738# a_77664_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15020 a_25227_30083# a_14926_31849# a_25145_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15021 a_40458_65206# a_16746_65208# a_40366_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15022 a_12093_69135# a_12039_69367# a_10747_68565# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X15023 a_33338_60186# a_12727_58255# a_33830_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15024 a_42466_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15025 a_10975_66407# a_14524_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X15026 VSS a_3024_67191# a_9503_68841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15027 a_19678_21906# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15028 VSS a_12355_15055# a_34738_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15029 a_18848_27765# a_13390_29575# a_19071_28111# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X1503 a_2376_23047# a_1689_10396# a_2518_22895# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15030 a_49798_10862# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15031 a_6641_72765# a_6224_73095# a_6559_72512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15032 a_4906_67509# a_5024_67885# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X15033 VSS a_6646_54135# a_7755_54999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15034 VSS VDD a_17670_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15035 a_26802_55488# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15036 VDD a_9547_54421# a_7265_56053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15037 VSS a_6831_63303# a_31031_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.6875e+11p ps=4.35e+06u w=650000u l=150000u
X15038 a_4748_58255# a_4311_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15039 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1504 ctopp a_8583_33551# inp_analog VDD sky130_fd_pr__pfet_01v8 ad=2.7075e+12p pd=2.185e+07u as=1.102e+12p ps=8.76e+06u w=1.9e+06u l=220000u M=4
X15040 a_21686_70226# a_12901_66665# a_21290_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15041 VSS a_12981_59343# a_47790_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15042 a_14949_31055# a_8197_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15043 VSS a_3247_20495# a_6637_20407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15044 VDD a_21049_41245# a_20655_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15045 VDD VSS a_35346_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15046 vcm_commonmode a_16362_17524# a_22386_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15047 VSS a_12985_16367# a_26706_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15048 VSS a_2419_48783# a_2971_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X15049 a_24716_31757# a_24632_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1505 a_11964_71855# a_11049_71855# a_11617_72097# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X15050 a_8384_40303# a_7905_40553# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15051 a_25961_47919# a_25015_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15052 a_24698_61190# a_12355_15055# a_24302_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15053 a_11490_74031# a_8575_74853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15054 a_49402_72234# VSS a_49494_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X15055 a_47486_55166# VDD a_47394_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15056 a_48794_16886# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15057 a_35069_32143# a_34267_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15058 a_7737_16917# a_7571_16917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15059 vcm_commonmode VSS a_31422_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 VSS a_2689_65103# a_7637_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X15060 a_12473_36341# a_31819_35073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X15061 a_46390_10862# a_16362_10496# a_46482_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15062 a_36350_71230# a_12901_66665# a_36842_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15063 a_36842_20504# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15064 a_27535_30503# a_37287_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15065 VDD VDD a_43378_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15066 a_36442_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15067 a_27999_41495# a_1761_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15068 a_30757_37455# a_30591_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X15069 VDD a_12981_62313# a_39362_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1507 a_6662_34025# a_5691_36727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X15070 a_5957_10927# a_5913_11169# a_5791_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15071 a_39362_64202# a_16362_64202# a_39454_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15072 a_28976_38567# a_28103_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15073 VSS a_7833_66415# a_8307_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15074 a_43470_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15075 a_37919_28111# a_30788_28487# a_37830_28111# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15076 VSS a_39459_44527# a_39565_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15077 a_26402_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15078 a_28714_60186# a_12981_59343# a_28318_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15079 VSS a_12899_11471# a_25702_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1508 VSS a_37459_51183# a_37478_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X15080 a_28714_19898# a_12895_13967# a_28318_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15081 VDD a_25764_51183# a_25939_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15082 VDD a_7078_36103# a_7019_35951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X15083 a_15271_41781# a_15459_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15084 a_8643_48767# a_8468_48841# a_8822_48829# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15085 VSS a_2824_70197# a_2960_70565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+11p ps=1.6e+06u w=540000u l=150000u
X15086 a_8485_71855# a_2451_72373# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15087 a_9187_56597# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X15088 a_9275_15253# a_9379_15039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15089 a_37354_12870# a_16362_12504# a_37446_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1509 VDD a_8003_72917# a_10509_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X15090 a_33689_28111# a_28757_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15091 VSS a_18197_44220# a_17889_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15092 a_16362_64202# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X15093 VDD a_1586_18695# a_1591_19631# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15094 VSS a_12901_66959# a_37750_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15095 a_4036_54421# a_1586_51335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15096 VDD a_34759_31029# a_39029_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15097 a_30326_69222# a_12901_66959# a_30818_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15098 a_41766_67214# a_12727_67753# a_41370_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15099 vcm_commonmode a_16362_63198# a_25398_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X151 VDD a_4482_57863# a_32785_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1510 VDD a_9367_29397# a_12158_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X15100 a_7948_38377# a_5363_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=6.3375e+11p pd=4.55e+06u as=0p ps=0u w=650000u l=150000u
X15101 a_26310_59182# a_12901_58799# a_26802_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15102 a_5991_21263# a_5547_21379# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15103 VDD a_2292_17179# a_7255_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15104 vcm_commonmode a_16362_20536# a_36442_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15105 a_39454_23548# a_16746_23546# a_39362_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15106 a_43270_27791# a_41597_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15107 VDD a_6821_26311# a_6773_27805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X15108 a_17766_70548# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15109 a_13097_40719# a_12831_41085# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1511 VSS a_16510_8760# a_16746_23546# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X15110 VSS a_2163_64381# a_2124_64507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15111 a_17274_60186# a_16362_60186# a_17366_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15112 a_11542_12381# a_11416_12283# a_11138_12267# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15113 a_38754_65206# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15114 a_31422_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15115 VDD a_12251_39069# a_12277_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15116 a_27983_40871# a_22671_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15117 a_27406_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15118 VDD a_9637_30511# a_10362_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15119 a_2325_71285# a_2107_71689# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X1512 VSS a_8575_74853# a_8781_71677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15120 a_1757_9839# a_1591_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X15121 a_36350_18894# a_16362_18528# a_36442_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15122 VSS a_2596_16911# a_3166_16911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15123 VSS a_20359_29199# a_36643_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X15124 a_28115_36919# a_27183_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X15125 a_8051_52047# a_7933_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15126 vcm_commonmode a_16362_64202# a_29414_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15127 a_35742_58178# a_12901_58799# a_35346_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15128 a_37750_9858# a_12985_19087# a_37354_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15129 VDD a_20195_49793# a_20156_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1513 a_46786_65206# a_10975_66407# a_46390_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15130 a_2781_23817# a_1591_23445# a_2672_23817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15131 a_18674_68218# a_12901_66959# a_18278_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15132 a_38850_61512# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15133 a_3981_10357# a_3763_10761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X15134 a_22097_52093# a_20535_51727# a_22015_51840# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15135 a_27333_32143# a_25953_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15136 a_46482_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15137 a_43378_66210# a_16362_66210# a_43470_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15138 a_48794_57174# a_10515_22671# a_48398_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15139 VSS a_4312_19061# a_1586_9991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1514 a_18979_30287# a_35079_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X15140 VDD a_4298_58951# a_4255_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X15141 vcm_commonmode a_16362_56170# a_19374_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15142 a_24698_15882# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15143 a_20925_40743# a_19245_39747# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X15144 a_6917_24233# a_3972_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15145 a_36607_34191# a_36430_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15146 VDD a_19069_50613# a_18959_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15147 a_6423_35190# a_4811_34855# a_5964_35015# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15148 a_10476_74031# a_10239_74575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X15149 a_2104_31599# a_1987_31812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1515 VDD a_43321_29941# a_43269_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15150 a_20378_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15151 VDD a_12727_13353# a_19282_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15152 a_33734_70226# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15153 a_22259_48981# a_22084_49007# a_22438_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15154 VDD a_3751_72373# a_4031_73095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X15155 a_32426_68218# a_16746_68220# a_32334_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15156 a_15871_39913# a_16265_39868# a_15931_39859# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X15157 VSS a_16510_8760# a_16746_9490# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X15158 a_37846_67536# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15159 a_10288_53047# a_10503_52828# a_10430_52854# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X1516 vcm_commonmode a_16362_64202# a_17366_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15160 a_31330_23914# a_16362_23548# a_31422_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15161 VDD a_10975_66407# a_41370_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15162 a_47394_24918# VSS a_47886_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15163 VSS a_37939_43455# a_37885_43777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15164 a_28730_50345# a_28688_50247# a_28648_50101# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15165 a_37354_57174# a_16362_57174# a_37446_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15166 a_5173_65327# a_3983_65327# a_5064_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15167 a_34834_8456# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15168 VDD a_1591_13103# a_1768_13103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15169 a_23694_62194# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1517 a_9560_60975# a_8772_63927# a_9370_60975# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X15170 a_4985_69725# a_3325_69135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15171 a_41462_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15172 a_30722_63198# a_15439_49525# a_30326_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15173 VSS a_16928_44007# a_16891_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15174 VSS a_6795_51157# a_6753_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X15175 VSS a_10515_23975# a_37750_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15176 VDD a_12947_8725# a_44382_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15177 VSS a_12985_19087# a_40762_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15178 VDD a_9972_69831# a_9314_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15179 a_4721_45199# a_4842_45467# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1518 a_22690_23914# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15180 VDD a_12024_30199# a_11978_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15181 a_7077_62313# a_7097_63151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X15182 a_41862_14480# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15183 a_41766_20902# a_11067_67279# a_41370_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15184 a_32612_51727# a_32582_51701# a_10680_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.2245e+11p ps=7.66e+06u w=1e+06u l=150000u M=4
X15185 a_4488_60431# a_4274_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15186 a_2426_31094# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X15187 VSS a_8423_39367# a_8127_39465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15188 VDD a_12257_56623# a_44382_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15189 a_12218_65693# a_11141_65327# a_12056_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1519 a_19282_22910# a_16362_22544# a_19374_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15190 a_5156_18543# a_4241_18543# a_4809_18785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15191 a_24794_24520# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15192 a_20905_32463# a_3339_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15193 a_32334_8854# a_12985_19087# a_32826_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15194 VSS a_12707_26159# a_14073_28157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15195 a_6816_37583# a_6786_37557# a_6559_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15196 a_5588_22467# a_3339_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15197 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15198 a_27406_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15199 a_5073_27247# a_4807_27613# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X152 a_31422_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1520 a_23298_9858# a_16362_9492# a_23390_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15200 a_23747_31055# a_23303_31171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15201 a_10747_68565# a_11943_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15202 a_26706_8854# a_12947_8725# a_26310_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15203 VDD a_22577_29111# a_22535_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15204 a_19258_47375# a_18500_47491# a_18695_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X15205 a_12410_55535# a_2419_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15206 a_33155_40191# a_1761_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15207 a_4124_64391# a_4339_64521# a_4266_64566# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X15208 a_5791_10927# a_5345_10927# a_5695_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15209 a_42374_10862# a_12985_16367# a_42866_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1521 a_23390_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15210 a_2008_28487# a_2216_28309# a_2150_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15211 VDD a_10506_29967# a_15575_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u M=2
X15212 VSS a_30412_42589# a_29513_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X15213 a_22411_42359# a_21479_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X15214 a_39758_72234# VDD a_39362_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15215 a_28810_23516# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15216 VDD a_18703_29199# a_37839_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15217 a_25306_20902# a_12985_7663# a_25798_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15218 a_32826_72556# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15219 a_40762_68218# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1522 a_12355_23983# a_11865_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X15220 a_25306_16886# a_16362_16520# a_25398_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15221 a_28410_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15222 a_11753_65327# a_11709_65569# a_11587_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15223 a_12901_58799# a_10055_58791# a_12913_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15224 VSS a_13837_39860# a_16969_38365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X15225 VDD a_12901_58799# a_35346_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15226 a_7815_19319# a_7841_12167# a_7989_19425# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15227 a_32334_62194# a_16362_62194# a_32426_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X15228 a_35742_11866# a_12985_16367# a_35346_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15229 VSS a_6619_73719# a_6098_73095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1523 a_34434_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15230 a_44474_17524# a_16746_17522# a_44382_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15231 a_2107_66415# a_1757_66415# a_2012_66415# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15232 a_18770_15484# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15233 a_18674_21906# a_12985_7663# a_18278_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15234 a_37307_51339# a_35676_49525# a_37465_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15235 VDD a_12877_16911# a_22294_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15236 a_48794_10862# a_12546_22351# a_48398_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15237 a_18278_8854# a_16362_8488# a_18370_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15238 a_8127_39465# a_8021_39221# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15239 a_43774_59182# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1524 VDD a_10472_26159# a_11130_22869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X15240 a_29322_15882# a_16362_15516# a_29414_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15241 a_31905_35073# a_30757_37455# a_31819_35073# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X15242 VSS a_11311_74005# a_11245_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15243 a_23774_49871# a_23830_49525# a_23774_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X15244 a_41370_16886# a_12899_11471# a_41862_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15245 a_27329_40747# a_27263_40871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15246 a_26706_69222# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15247 a_15683_40767# a_12343_42333# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X15248 VDD a_5340_32687# a_5515_32661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15249 a_5905_44905# a_6095_44807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1525 a_36746_57174# a_10515_22671# a_36350_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15250 VSS a_12983_63151# a_30722_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15251 a_48490_16520# a_16746_16518# a_48398_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15252 a_8123_34319# a_6372_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15253 vcm_commonmode a_16362_13508# a_45478_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15254 a_7449_60431# a_6737_60431# a_7377_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15255 a_19282_11866# a_10055_58791# a_19774_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15256 VDD a_2127_4943# a_2603_4943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15257 a_8491_35727# a_5915_35943# a_8397_35727# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X15258 VDD a_3143_66972# a_7577_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15259 vcm_commonmode a_16362_23548# a_28410_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1526 a_47790_8854# a_12947_8725# a_47394_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15260 a_2012_36861# a_1761_35951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15261 a_42466_8488# a_16746_8486# a_42374_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15262 a_32426_21540# a_16746_21538# a_32334_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15263 VSS a_12901_58799# a_20682_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15264 a_16744_41605# a_15775_41317# a_16707_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X15265 a_47790_58178# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15266 VDD a_8636_63669# a_7891_64213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X15267 a_18370_8488# a_16746_8486# a_18278_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15268 vcm_commonmode a_16362_15516# a_18370_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15269 VDD a_3173_53333# a_3203_53686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1527 vcm_commonmode a_16362_68218# a_43470_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15270 VDD a_15439_49525# a_30326_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15271 VDD a_1923_59583# a_6519_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15272 a_22386_13508# a_16746_13506# a_22294_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15273 a_2121_72943# a_1643_72917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15274 VDD a_34395_31287# a_33798_31145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X15275 a_35438_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15276 a_26889_50337# a_26671_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X15277 a_47486_63198# a_16746_63200# a_47394_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15278 a_2242_24566# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X15279 VSS a_4314_40821# a_5414_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1528 a_12792_51017# a_11711_50645# a_12445_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X15280 VSS a_10515_22671# a_24698_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15281 VSS a_12901_66665# a_38754_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15282 a_21686_55166# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15283 a_1644_76181# a_1823_76181# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15284 a_34434_66210# a_16746_66212# a_34342_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15285 VSS a_11719_28023# a_12631_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15286 a_6743_29673# a_5449_25071# a_6825_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15287 a_27314_61190# a_12981_59343# a_27806_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15288 a_36442_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15289 VDD a_24931_42657# a_24755_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1529 a_19678_67214# a_12727_67753# a_19282_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15290 VDD a_35319_34191# a_35425_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15291 a_12702_25615# a_10472_26159# a_12394_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15292 VDD a_12901_66665# a_39362_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15293 a_18278_19898# a_11067_67279# a_18770_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15294 a_39454_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15295 a_32730_61190# a_12355_15055# a_32334_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15296 VSS a_31847_36893# a_31787_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15297 a_12901_66959# a_11619_56615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15298 a_38450_65206# a_16746_65208# a_38358_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15299 a_12085_64239# a_11943_63125# a_12013_64239# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X153 a_2647_31421# a_2473_34293# a_2284_31287# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1530 a_2824_70197# a_3280_70501# a_3238_70589# VSS sky130_fd_pr__nfet_01v8 ad=1.47e+11p pd=1.54e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15300 a_2882_73309# a_2163_73085# a_2319_73180# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15301 VSS VSS a_43774_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15302 a_40762_21906# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15303 VSS a_6816_19355# a_7159_22583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15304 a_2835_62215# a_3108_62043# a_3066_62069# VSS sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15305 a_37354_20902# a_16362_20536# a_37446_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15306 a_43378_57174# a_12257_56623# a_43870_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15307 a_15661_29199# a_6459_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X15308 a_32507_50959# a_4482_57863# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15309 a_11495_16341# a_11320_16367# a_11674_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1531 VSS a_8132_53511# a_9405_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15310 vcm_commonmode VSS a_21382_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15311 a_26310_67214# a_12983_63151# a_26802_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15312 VDD a_29545_28023# a_11619_3303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X15313 a_30818_65528# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15314 VSS a_12899_11471# a_33734_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15315 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15316 a_5064_45743# a_3983_45743# a_4717_45985# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X15317 VDD a_6435_74005# a_6422_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15318 a_30326_55166# VSS a_30418_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15319 VDD a_7939_30503# a_26219_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1532 a_22399_32143# a_22148_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15320 a_28607_29673# a_4811_34855# a_28513_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X15321 VSS a_12727_13353# a_46786_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15322 a_43774_12870# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15323 a_20682_24918# VSS a_20286_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15324 VSS a_20359_29199# a_35447_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X15325 a_8485_29673# a_6752_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15326 a_20778_57496# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15327 a_26706_22910# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15328 a_41370_9858# a_12546_22351# a_41862_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15329 a_8480_37039# a_5915_35943# a_8177_37013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X1533 VDD a_27411_50069# a_27869_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15330 a_30326_14878# a_12877_14441# a_30818_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15331 VSS a_12985_7663# a_30722_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15332 a_34342_59182# a_12901_58799# a_34834_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15333 a_15575_28879# a_12631_28585# a_15829_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15334 a_17274_9858# a_12546_22351# a_17766_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15335 a_35932_37601# a_35647_38053# a_36579_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X15336 a_47394_58178# a_10515_22671# a_47886_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15337 VSS a_12899_10927# a_19678_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15338 a_5871_47594# a_5963_47349# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15339 vcm_commonmode VSS a_29414_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1534 a_49798_56170# a_12257_56623# a_49402_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15340 a_23694_15882# a_12877_14441# a_23298_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15341 VSS a_12877_16911# a_20682_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15342 VDD a_7000_43541# a_14655_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15343 a_47790_11866# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15344 VSS a_24959_30503# a_34062_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15345 VDD a_4647_63937# a_4608_63811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15346 a_35907_31055# a_27535_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X15347 a_30079_47375# a_27869_50095# a_29987_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X15348 a_27806_9460# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15349 VSS a_12355_15055# a_45782_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1535 VSS a_31551_31751# a_30155_32375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X15350 VDD a_12755_53030# a_12901_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15351 a_28963_28853# a_4811_34855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15352 VDD a_16744_40517# a_16265_39868# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X15353 a_30542_51433# a_28881_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15354 VSS a_2319_54684# a_2250_54813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15355 a_23390_62194# a_16746_62196# a_23298_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15356 a_3238_70589# a_2960_70565# a_3166_70589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15357 a_24794_58500# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15358 vcm_commonmode a_16362_18528# a_20378_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15359 a_11396_60975# a_7773_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X1536 VSS a_1586_40455# a_5179_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15360 VSS a_8583_33551# a_33479_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15361 a_6010_56989# a_5291_56765# a_5447_56860# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X15362 a_27710_14878# a_12727_15529# a_27314_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15363 VSS a_10055_58791# a_24698_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15364 VSS a_12481_54447# a_12407_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15365 vcm_commonmode a_16362_17524# a_33430_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15366 VDD VSS a_46390_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15367 VSS a_28089_31157# a_28446_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X15368 VDD a_11067_13095# a_15660_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15369 a_4328_10761# a_3413_10389# a_3981_10357# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X1537 a_18413_47919# a_18243_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X15370 VDD a_2411_18517# a_10659_9813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15371 a_10317_67191# a_9513_65301# a_10480_67075# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15372 VDD a_8273_42479# a_8827_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15373 a_24910_31599# a_23747_31055# a_24591_31599# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u w=650000u l=150000u
X15374 a_23271_50943# a_23096_51017# a_23450_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15375 VSS a_11067_13095# a_36746_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15376 VSS a_18045_38017# a_19283_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15377 a_13615_48579# a_5039_42167# a_13543_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15378 a_39758_8854# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15379 VSS a_12231_55509# a_12165_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1538 VSS a_12899_10927# a_28714_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15380 a_34834_21508# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15381 a_34434_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15382 VSS a_3983_12015# a_4065_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15383 VDD a_2944_57960# a_2882_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15384 a_3413_10389# a_3247_10389# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15385 a_37354_65206# a_16362_65206# a_37446_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15386 a_14049_40693# a_13067_38517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15387 a_41462_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15388 a_47886_20504# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15389 a_47486_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1539 a_6725_45205# a_6559_45205# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X15390 VSS a_12985_19087# a_49798_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15391 a_21290_70226# a_16362_70226# a_21382_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15392 a_10791_15529# a_10673_15055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15393 a_13357_32143# a_7695_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15394 vcm_commonmode a_16362_69222# a_49494_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15395 a_37846_12472# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15396 VDD a_1689_10396# a_1633_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X15397 a_35346_13874# a_16362_13508# a_35438_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15398 VDD a_12546_22351# a_41370_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15399 VSS a_27175_47375# a_27509_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X154 VSS vcm_commonmode VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u M=80
X1540 a_3049_14343# a_2873_13879# a_3212_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15400 a_12993_50345# a_9963_50959# a_12993_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15401 VDD a_11067_67279# a_24302_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15402 a_48398_12870# a_16362_12504# a_48490_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15403 a_27406_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15404 a_21178_52047# a_19576_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15405 a_44778_61190# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15406 a_43470_59182# a_16746_59184# a_43378_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15407 vcm_commonmode a_16362_56170# a_40458_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15408 a_37446_24552# VDD a_37354_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15409 a_10299_11703# a_9491_12297# a_10473_11809# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1541 VSS a_12981_62313# a_41766_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15410 a_27710_71230# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15411 a_26402_69222# a_16746_69224# a_26310_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15412 vcm_commonmode a_16362_66210# a_23390_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15413 VSS a_2989_45717# a_2923_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15414 VSS a_17927_31573# a_17488_48731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15415 a_25306_24918# VSS a_25398_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15416 a_24223_31171# a_15548_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15417 VDD a_11851_64391# a_11803_64239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15418 VDD a_12983_63151# a_35346_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15419 VDD a_23271_50943# a_22989_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X1542 a_38450_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15420 a_46390_7850# VDD a_46882_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15421 a_25398_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15422 a_28318_60186# a_16362_60186# a_28410_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15423 VSS a_12981_59343# a_21686_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15424 vcm_commonmode VSS a_44474_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15425 a_18370_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15426 VDD a_4528_26159# a_6993_23555# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15427 VSS a_22132_44129# a_25263_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15428 VDD a_15557_52245# a_15285_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X15429 vcm_commonmode a_16362_65206# a_27406_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1543 a_10073_23439# a_8569_24527# a_9971_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15430 VDD a_12985_16367# a_18278_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15431 VDD a_8273_42479# a_8123_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15432 VDD a_21273_30485# a_21012_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15433 a_25939_51157# a_25764_51183# a_26118_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X15434 a_11399_18543# a_10883_18543# a_11304_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X15435 a_29322_23914# a_16362_23548# a_29414_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15436 a_36842_62516# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15437 a_28714_7850# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15438 a_2886_46831# a_2656_45895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15439 a_41370_67214# a_16362_67214# a_41462_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1544 a_2041_61519# a_1954_61677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15440 a_46786_58178# a_12901_58799# a_46390_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15441 VDD a_12981_59343# a_40366_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15442 a_12360_21263# a_12263_20969# a_11763_21237# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15443 vcm_commonmode a_16362_57174# a_17366_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15444 a_23739_29245# a_23685_29111# a_23643_29245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15445 a_29718_68218# a_12901_66959# a_29322_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15446 a_49894_61512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15447 a_2107_39049# a_1757_38677# a_2012_39037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15448 a_21382_55166# VDD a_21290_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15449 a_22690_16886# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1545 a_9215_61127# a_9424_60949# a_9382_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X15450 VSS a_3987_19623# a_7571_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15451 a_9435_65327# a_7803_55509# a_9363_65327# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X15452 a_20286_10862# a_16362_10496# a_20378_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15453 VSS a_5211_24759# a_9135_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15454 a_9179_22351# a_8671_22671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15455 a_21829_48161# a_21611_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X15456 a_17983_41855# a_16744_41605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X15457 a_4595_45743# a_4149_45743# a_4499_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15458 a_4811_34855# a_23685_29111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X15459 a_22105_30761# a_15548_30761# a_22014_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1546 a_21686_70226# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15460 VDD a_2787_30503# a_24714_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15461 VDD VDD a_33338_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15462 a_34738_69222# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15463 VDD a_35033_38780# a_34639_38825# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15464 VDD a_12947_71576# a_30326_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15465 VDD a_12355_15055# a_26310_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15466 a_25953_32143# a_25605_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X15467 a_5475_74895# a_5441_72399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15468 VSS a_2163_63293# a_2124_63419# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15469 a_5823_28585# a_6162_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1547 vcm_commonmode a_16362_59182# a_46482_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15470 VSS a_4482_57863# a_33071_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X15471 a_2847_15039# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15472 VSS a_27183_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X15473 a_2693_68021# a_2475_68425# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15474 a_2284_31287# a_2473_34293# a_2426_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15475 a_35346_58178# a_16362_58178# a_35438_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15476 VDD a_2040_43401# a_2216_42997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15477 a_23753_51433# a_23487_50095# a_23193_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15478 a_2203_15113# a_1757_14741# a_2107_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15479 VSS a_3305_38671# a_3705_40079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X1548 a_20378_68218# a_16746_68220# a_20286_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15480 a_21686_63198# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15481 vcm_commonmode a_16362_22544# a_49494_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15482 a_18278_68218# a_16362_68218# a_18370_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15483 a_31822_7452# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15484 a_48398_57174# a_16362_57174# a_48490_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15485 VSS a_9863_51420# a_9794_51549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15486 a_11898_10205# a_11179_9981# a_11335_10076# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X15487 a_35346_17890# a_12899_10927# a_35838_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15488 VSS a_12947_23413# a_35742_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15489 a_2503_34319# a_2473_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X1549 VDD a_3016_60949# a_5089_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X15490 a_24302_11866# a_16362_11500# a_24394_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15491 VSS a_12546_22351# a_20682_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15492 VDD a_12899_10927# a_42374_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15493 a_1761_35951# a_1591_35951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15494 a_43470_12504# a_16746_12502# a_43378_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15495 VDD a_36464_49783# a_36465_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X15496 a_15259_46805# a_15607_46805# a_15541_46831# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X15497 VSS a_33641_29967# a_34613_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15498 a_26402_22544# a_16746_22542# a_26310_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15499 a_22995_30663# a_7939_30503# a_23169_30539# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X155 a_41766_22910# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1550 a_17039_51157# a_19439_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X15500 vcm_commonmode a_16362_70226# a_35438_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15501 a_75199_38962# a_75111_39506# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15502 a_28195_35327# a_27429_35301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X15503 VSS a_7210_55081# a_7115_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X15504 a_25398_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15505 a_39362_16886# a_12899_11471# a_39854_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15506 a_43003_30761# a_33641_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15507 a_40366_11866# a_10055_58791# a_40858_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15508 VSS a_28817_29111# a_28817_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15509 VSS a_12983_63151# a_28714_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1551 a_6921_72943# a_8003_72917# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X15510 a_25702_64202# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15511 a_1761_50639# a_1591_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X15512 result_out[13] a_1644_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15513 a_23298_21906# a_11067_21583# a_23790_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15514 a_26221_29423# a_26191_29397# a_26137_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15515 a_38315_38053# a_37076_37253# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X15516 a_23298_17890# a_16362_17524# a_23390_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15517 VDD a_12727_58255# a_33338_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15518 a_17366_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15519 a_1757_43029# a_1591_43029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1552 a_32371_32117# a_32367_28309# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X15520 vcm_commonmode a_16362_61190# a_38450_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15521 a_30326_63198# a_16362_63198# a_30418_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15522 VSS a_12901_58799# a_18674_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15523 a_42466_18528# a_16746_18526# a_42374_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15524 VDD a_12901_58799# a_46390_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15525 a_22690_57174# a_10515_22671# a_22294_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15526 a_4233_25321# a_3325_18543# a_4161_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15527 VDD a_38628_47349# a_29927_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15528 VDD a_1923_54591# a_5132_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15529 a_46786_11866# a_12985_16367# a_46390_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1553 a_39362_8854# a_16362_8488# a_39454_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15530 a_2969_41909# a_2751_42313# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15531 a_5531_53903# a_5258_54223# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15532 a_34342_67214# a_12983_63151# a_34834_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15533 a_11491_60975# a_10975_60975# a_11396_60975# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X15534 a_29814_15484# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15535 vcm_commonmode a_16362_10496# a_17366_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15536 a_29718_21906# a_12985_7663# a_29322_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15537 a_26310_12870# a_12877_16911# a_26802_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15538 a_2847_49855# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15539 a_30818_10464# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1554 a_35346_24918# VSS a_35838_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15540 VDD a_33080_37149# a_32181_36893# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X15541 a_47394_66210# a_10975_66407# a_47886_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15542 a_4127_50069# a_2840_66103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X15543 a_17003_49770# a_17095_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X15544 a_18907_48829# a_18653_48502# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15545 a_19678_55166# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15546 vcm_commonmode a_16362_14512# a_43470_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15547 a_19678_13874# a_12877_16911# a_19282_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15548 a_3186_25321# a_2315_24540# a_3104_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15549 a_34738_22910# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1555 a_34342_7850# VDD a_34834_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15550 vcm_commonmode a_16362_59182# a_32426_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15551 a_22386_9492# a_16746_9490# a_22294_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15552 vcm_commonmode VSS a_26402_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15553 a_24953_47753# a_23763_47381# a_24844_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15554 VSS a_32611_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X15555 a_41862_56492# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15556 a_17696_29967# a_16228_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X15557 VDD a_12516_7093# a_27314_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15558 a_24794_66532# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15559 a_2100_24759# a_2315_24540# a_2242_24566# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X1556 VSS a_28011_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X15560 a_10607_29423# a_8485_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X15561 a_21290_63198# a_12981_62313# a_21782_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15562 a_19374_60186# a_16746_60188# a_19282_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15563 VDD a_12985_19087# a_37354_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15564 a_19374_19532# a_16746_19530# a_19282_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15565 VSS a_24892_38237# a_23993_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X15566 a_20378_14512# a_16746_14510# a_20286_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15567 a_24302_56170# a_16362_56170# a_24394_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15568 VDD a_11710_58487# a_11711_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15569 a_22639_50639# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X1557 a_29942_30663# a_30052_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15570 a_30181_38571# a_30115_38695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15571 a_33543_39095# a_32611_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15572 VSS VDD a_36746_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15573 a_8095_40303# a_6372_38279# a_7905_40553# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X15574 a_29118_50639# a_28959_49783# a_29038_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X15575 a_40762_70226# a_12901_66665# a_40366_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15576 VDD a_4043_44343# a_2656_45895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X15577 a_28810_65528# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15578 a_25306_62194# a_12355_15055# a_25798_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15579 VSS a_8753_66103# a_7987_64213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1558 VSS a_32887_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X15580 VSS a_4968_60405# a_4906_60431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15581 VSS a_5013_20473# a_4947_20541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15582 a_17651_30485# a_17415_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15583 VSS a_12901_66665# a_49798_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15584 a_45478_66210# a_16746_66212# a_45386_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15585 a_47486_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15586 a_18770_57496# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15587 a_1761_35407# a_1591_35407# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X15588 a_22285_47919# a_21095_47919# a_22176_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15589 VDD VSS a_22294_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1559 a_29718_13874# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15590 VSS a_12985_7663# a_28714_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15591 VSS a_1586_51335# a_1591_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15592 VSS a_30716_51701# a_30663_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X15593 a_43774_61190# a_12355_15055# a_43378_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15594 a_35346_9858# a_16362_9492# a_35438_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15595 VSS a_12899_10927# a_40762_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15596 a_18915_42089# a_17983_41855# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X15597 VDD a_7931_10357# a_7862_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15598 a_26706_71230# a_12947_71576# a_26310_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15599 a_15959_44031# a_15193_44005# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X156 a_16746_56172# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X1560 a_19026_31375# a_3339_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X15600 VSS a_9989_46831# a_13461_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15601 a_49494_65206# a_16746_65208# a_49402_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15602 VSS a_12877_16911# a_18674_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15603 a_45478_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15604 a_48398_20902# a_16362_20536# a_48490_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15605 a_13867_37782# a_13909_37571# a_13867_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15606 a_22690_10862# a_12546_22351# a_22294_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15607 a_5909_71855# a_4719_71855# a_5800_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X15608 a_2369_12925# a_2325_12533# a_2203_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15609 a_39454_57174# a_16746_57176# a_39362_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1561 a_49494_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15610 a_5778_43933# a_4701_43567# a_5616_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15611 a_47790_60186# a_12981_59343# a_47394_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15612 a_47790_19898# a_12895_13967# a_47394_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15613 VSS a_12899_11471# a_44778_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15614 a_41766_13874# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15615 a_7896_18695# a_8104_18517# a_8038_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15616 result_out[1] a_1644_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15617 a_8689_17999# a_5535_18012# a_8111_18825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15618 a_42466_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15619 a_11981_20495# a_3987_19623# a_11763_20407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1562 a_38358_56170# a_16362_56170# a_38450_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15620 VDD a_11067_67279# a_32334_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15621 a_31822_18496# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15622 a_31726_24918# VSS a_31330_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15623 a_11413_25321# a_9955_20969# a_11340_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15624 a_25398_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15625 VSS a_32134_49159# a_32135_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15626 vcm_commonmode a_16362_12504# a_32426_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15627 vcm_commonmode a_16362_63198# a_44474_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15628 a_45386_59182# a_12901_58799# a_45878_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15629 VSS a_12895_13967# a_17670_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1563 a_44874_7452# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15630 VDD a_38436_29941# a_38883_29217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15631 a_21686_16886# a_12727_13353# a_21290_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15632 a_30991_35307# a_26433_39631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15633 a_36842_70548# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15634 a_42283_38007# a_41351_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15635 a_33430_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15636 VSS a_1586_69367# a_1959_68053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15637 VDD a_33591_32375# a_28547_51175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X15638 a_4274_60431# a_4187_60673# a_3870_60563# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X15639 VSS a_43227_28309# a_43175_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1564 a_40762_7850# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15640 a_33734_69222# a_12516_7093# a_33338_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15641 a_22535_28879# a_18053_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15642 VSS a_2163_59585# a_2124_59459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15643 a_16746_12502# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X15644 a_21382_63198# a_16746_63200# a_21290_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15645 a_19596_42919# a_18627_42943# a_19500_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X15646 a_46482_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15647 a_19282_70226# a_16362_70226# a_19374_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15648 a_22786_59504# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15649 VSS a_8583_33551# a_32743_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1565 a_10899_28879# a_10648_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15650 a_25013_31599# a_23119_31599# a_24910_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15651 a_18674_14878# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15652 VSS a_5915_30287# a_7825_36815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X15653 a_21387_38591# a_19780_39429# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X15654 VSS VDD a_38754_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15655 vcm_commonmode a_16362_18528# a_31422_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15656 a_43774_9858# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15657 a_20964_31029# a_20905_32143# a_21356_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15658 a_21371_50959# a_13643_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X15659 a_48794_7850# VDD a_48398_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1566 a_7910_38671# a_3949_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=5.72e+06u as=0p ps=0u w=1e+06u l=150000u
X15660 VDD a_3327_9308# a_8117_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X15661 a_9945_47919# a_9779_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15662 a_37750_68218# a_12901_66959# a_37354_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15663 VSS a_12355_65103# a_34738_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15664 a_39299_48783# a_20635_29415# a_39210_48783# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X15665 VDD a_12899_11471# a_34342_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15666 a_12663_40871# a_32555_43777# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X15667 VDD a_4987_52508# a_4918_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15668 a_19678_9858# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15669 a_14553_28585# a_9731_22895# a_14471_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1567 a_11611_12252# a_11416_12283# a_11921_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X15670 VSS a_11067_13095# a_47790_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15671 VDD a_1683_27399# a_1683_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15672 VDD a_32672_49007# a_33681_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15673 a_45878_21508# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15674 a_45478_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15675 VSS a_12546_22351# a_29718_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15676 a_48398_65206# a_16362_65206# a_48490_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15677 VSS a_12947_56817# a_37750_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15678 VDD a_8459_71285# a_7707_70741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15679 a_30326_56170# a_12947_56817# a_30818_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1568 VDD a_12139_18517# a_7377_18012# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15680 VDD a_12727_13353# a_38358_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15681 a_35838_13476# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15682 VSS a_4417_22671# a_9253_24011# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15683 a_24698_64202# a_12355_65103# a_24302_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15684 a_22577_29111# a_2235_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15685 a_9307_30663# a_6773_27805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15686 a_39454_10496# a_16746_10494# a_39362_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15687 a_41967_31375# a_41427_52263# a_41795_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15688 a_29483_42943# a_28717_42917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X15689 a_46390_13874# a_16362_13508# a_46482_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1569 VDD a_12899_11471# a_32334_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15690 VSS a_11480_23957# a_11424_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15691 a_25398_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15692 a_9278_55311# a_7210_55081# a_9468_55311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15693 a_15941_31849# a_16087_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15694 VSS a_39244_41953# a_38345_42044# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X15695 a_42770_62194# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15696 a_4212_15823# a_3998_15823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15697 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X15698 a_20496_49551# a_20282_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15699 a_39362_67214# a_16362_67214# a_39454_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X157 a_38358_21906# a_16362_21540# a_38450_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1570 a_31726_62194# a_12981_62313# a_31330_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15700 a_25702_72234# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15701 vcm_commonmode a_16362_67214# a_21382_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15702 a_6606_16733# a_5529_16367# a_6444_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15703 a_22148_32259# a_20905_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15704 VDD a_12727_67753# a_33338_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15705 a_26310_8854# a_12985_19087# a_26802_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15706 a_43870_24520# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15707 a_10509_62985# a_9319_62613# a_10400_62985# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15708 a_33430_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15709 VDD a_12983_63151# a_46390_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1571 a_3295_62083# a_3983_59887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X15710 VDD a_40783_46831# a_15607_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15711 vcm_commonmode a_16362_9492# a_45478_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15712 VDD a_2292_43291# a_6655_46261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15713 a_16362_67214# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X15714 VSS a_3987_19623# a_5547_21379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15715 a_18674_55166# a_18602_55312# a_18278_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15716 VDD a_1867_32839# a_1867_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15717 a_46482_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15718 VSS a_12981_59343# a_32730_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15719 a_33734_22910# a_11067_21583# a_33338_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1572 VDD a_6372_38279# a_6786_37557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X15720 a_29414_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15721 a_7657_64489# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15722 a_9649_61225# a_7210_55081# a_9215_61127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15723 a_2216_16885# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15724 VDD a_12985_16367# a_29322_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15725 VDD VSS a_20286_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15726 VDD a_12901_66959# a_19282_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15727 a_44382_20902# a_12985_7663# a_44874_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15728 VSS a_18197_36604# a_17889_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15729 a_44382_16886# a_16362_16520# a_44474_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1573 a_21387_39679# a_19596_40743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X15730 a_19678_63198# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15731 a_5418_48829# a_2595_47653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15732 a_47886_62516# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15733 a_7905_40553# a_7097_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15734 a_17211_49373# a_16587_49007# a_17103_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X15735 vcm_commonmode a_16362_57174# a_28410_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15736 a_4947_20541# a_3987_19623# a_4584_20407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15737 VDD a_5595_63125# a_5553_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X15738 a_34342_12870# a_12877_16911# a_34834_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15739 a_37750_21906# a_12985_7663# a_37354_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1574 a_2122_20719# a_1945_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15740 a_32426_55166# VDD a_32334_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15741 a_33734_16886# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15742 a_17274_22910# a_10515_23975# a_17766_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15743 a_31330_10862# a_16362_10496# a_31422_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15744 a_21290_71230# a_12901_66665# a_21782_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15745 VSS a_19442_28585# a_19541_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X15746 a_21782_20504# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15747 a_21382_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15748 VDD a_12981_62313# a_24302_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15749 VSS a_32795_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X1575 a_39362_23914# a_12947_23413# a_39854_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15750 a_24302_64202# a_16362_64202# a_24394_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15751 a_45782_69222# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15752 VSS a_7707_70741# a_7624_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15753 VSS a_15968_36061# a_15069_35805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X15754 vcm_commonmode VSS a_34434_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15755 a_10117_14013# a_9083_13879# a_10045_14013# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15756 a_5357_62313# a_4797_62063# a_5274_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X15757 a_28192_48783# a_26514_47375# a_28108_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15758 vcm_commonmode a_16362_23548# a_47486_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15759 a_40315_31849# a_7295_44647# a_40233_31605# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1576 a_39362_19898# a_16362_19532# a_39454_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15760 a_6980_45565# a_6361_44655# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15761 VDD a_1586_9991# a_1591_16917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15762 a_6921_72943# a_8003_72917# a_7615_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X15763 a_25306_70226# a_12516_7093# a_25798_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15764 a_46390_58178# a_16362_58178# a_46482_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15765 VDD a_12727_15529# a_27314_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15766 a_23669_49257# a_23019_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15767 VDD a_6738_19783# a_6743_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X15768 a_22294_12870# a_16362_12504# a_22386_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15769 a_51936_39932# a_49876_37608# a_51714_39886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.24e+12p ps=9.24e+06u w=2e+06u l=150000u M=2
X1577 a_43378_72234# VDD a_43870_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15770 VSS a_12901_66959# a_22690_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15771 a_49798_68218# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15772 a_11901_63151# a_11053_62607# a_11829_63151# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15773 a_43539_29967# a_43680_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15774 a_18351_37503# a_17585_37477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X15775 vcm_commonmode a_16362_15516# a_37446_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15776 a_46390_17890# a_12899_10927# a_46882_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15777 a_27793_51733# a_27627_51733# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X15778 a_41462_13508# a_16746_13506# a_41370_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15779 a_12671_37782# a_12343_36893# a_12671_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1578 a_19878_49683# a_20195_49793# a_20153_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X15780 VSS a_3417_31599# a_3799_31063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15781 a_24394_23548# a_16746_23546# a_24302_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15782 VDD a_33868_47349# a_33802_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15783 vcm_commonmode a_16362_20536# a_21382_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15784 a_12831_41085# a_12651_41085# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15785 a_37446_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15786 a_28810_10464# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15787 a_39758_18894# a_12899_10927# a_39362_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15788 VSS a_10515_22671# a_43774_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15789 a_40762_55166# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1579 a_43870_21508# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15790 a_33957_49007# a_32856_48463# a_33857_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.47e+11p ps=1.54e+06u w=420000u l=150000u
X15791 a_9418_12342# a_3327_9308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15792 vcm_commonmode a_16362_70226# a_46482_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15793 VSS a_12727_67753# a_26706_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15794 a_23694_65206# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15795 VDD a_1915_20394# a_1867_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15796 VSS a_21479_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X15797 a_16375_41807# a_15931_39859# a_16012_41959# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X15798 a_22671_43439# a_1761_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15799 a_21290_18894# a_16362_18528# a_21382_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X158 VSS a_14926_31849# a_25145_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X1580 a_43470_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15800 a_37354_19898# a_11067_67279# a_37846_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15801 a_27745_27275# a_23928_28585# a_27659_27275# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X15802 a_41370_68218# a_12727_67753# a_41862_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15803 vcm_commonmode a_16362_62194# a_36442_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15804 VSS a_12447_29199# a_40139_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X15805 VDD a_15193_42917# a_16648_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X15806 a_40458_60186# a_16746_60188# a_40366_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15807 VDD a_12727_58255# a_44382_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15808 a_40458_19532# a_16746_19530# a_40366_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15809 a_1761_25071# a_1591_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1581 VSS a_5671_21495# a_11981_20495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X15810 a_20682_58178# a_12901_58799# a_20286_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15811 a_14831_50095# a_14445_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X15812 a_19282_63198# a_12981_62313# a_19774_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15813 a_4487_64239# a_4339_64521# a_4124_64391# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X15814 VSS a_12901_58799# a_29718_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15815 a_23790_61512# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15816 a_26706_56170# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15817 a_29207_36415# a_28441_36389# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X15818 a_18145_31849# a_16917_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15819 VDD a_7000_43541# a_15575_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1582 a_40366_14878# a_16362_14512# a_40458_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15820 a_31422_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15821 a_18370_14512# a_16746_14510# a_18278_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15822 a_27806_16488# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15823 VSS a_19807_28111# a_36459_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15824 a_45386_67214# a_12983_63151# a_45878_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15825 vcm_commonmode a_16362_10496# a_28410_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15826 VDD a_1803_19087# a_30855_41809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X15827 a_27417_32509# a_27387_32373# a_27333_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15828 a_6662_34025# a_6372_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X15829 a_19416_51017# a_18501_50645# a_19069_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1583 a_25987_41317# a_25221_41281# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X15830 a_33430_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15831 a_4035_11989# a_4211_11989# a_4163_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X15832 a_4680_32687# a_4563_32900# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15833 a_45782_22910# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15834 a_18278_69222# a_12901_66959# a_18770_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15835 VSS a_16012_41959# a_15189_39889# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15836 a_22786_67536# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15837 VDD a_2235_30503# a_7030_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15838 a_23592_52271# a_23193_52245# a_22921_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X15839 a_32334_24918# a_12899_3855# a_32826_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1584 VDD a_40691_47375# a_20359_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X15840 a_22294_57174# a_16362_57174# a_22386_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15841 a_21800_36165# a_20927_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X15842 VSS a_12899_10927# a_38754_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15843 a_9613_48981# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X15844 a_42770_15882# a_12877_14441# a_42374_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15845 a_15697_28335# a_14912_27497# a_15599_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X15846 VSS a_8540_42167# a_8383_43255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15847 a_4605_64061# a_4127_63669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15848 VSS a_10515_23975# a_22690_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15849 VSS a_4124_64391# a_4075_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1585 a_30052_32117# a_30203_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15850 a_19374_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15851 a_49798_21906# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15852 a_5693_39465# a_5490_41365# a_5259_39367# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X15853 a_12283_36919# a_12677_36893# a_12343_36893# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X15854 a_2672_51183# a_1591_51183# a_2325_51425# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X15855 VDD a_77285_39738# a_77098_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X15856 a_16891_43177# a_15959_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15857 a_4211_11989# a_1929_12131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15858 a_26465_48463# a_26187_48801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X15859 VSS VDD a_47790_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1586 VSS VDD a_26706_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15860 a_4499_48841# a_4149_48469# a_4404_48829# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X15861 a_4404_20719# a_3969_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15862 a_43870_58500# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15863 a_39758_13874# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15864 VSS a_10055_58791# a_43774_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15865 a_7994_42479# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15866 a_9418_12015# a_3327_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15867 a_7373_62927# a_6515_62037# a_7071_62581# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X15868 a_2926_31965# a_1849_31599# a_2764_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15869 VSS a_11067_21583# a_26706_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1587 a_36520_39429# a_35647_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X15870 a_7301_30511# a_5993_32687# a_7229_30511# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15871 a_41766_62194# a_12981_62313# a_41370_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15872 a_29814_57496# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15873 a_2369_19631# a_2325_19873# a_2203_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15874 VSS a_7862_34025# a_26985_31605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15875 a_6666_53359# a_5541_53609# a_6666_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X15876 a_24698_72234# VDD a_24302_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15877 VDD a_2191_68565# a_4075_63151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15878 VDD a_12901_58799# a_20286_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15879 a_30663_49257# a_30609_49159# a_30567_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1588 a_28714_60186# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15880 VDD a_4417_22671# a_8113_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15881 a_20682_11866# a_12985_16367# a_20286_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15882 a_20778_9460# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15883 VSS a_12877_16911# a_29718_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15884 VSS a_5239_48767# a_5173_48841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X15885 a_38754_60186# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15886 a_37446_58178# a_16746_58180# a_37354_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15887 a_38754_19898# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15888 a_2939_33535# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15889 a_40366_70226# a_16362_70226# a_40458_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1589 a_27406_58178# a_16746_58180# a_27314_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15890 VSS a_35493_43421# a_35185_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15891 a_11881_67325# a_11659_66567# a_11793_67325# VSS sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X15892 a_12605_54991# a_12371_53903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15893 a_32730_64202# a_12355_65103# a_32334_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15894 VSS a_11999_67477# a_12805_68367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15895 a_2834_29967# a_1757_29973# a_2672_30345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15896 a_40219_48783# a_20635_29415# a_40050_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15897 a_33430_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15898 a_39854_22512# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15899 VSS a_1952_60431# a_4692_55541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X159 a_37951_42089# a_38011_42035# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.57899e+15p ps=1.51821e+10u w=800000u l=150000u M=2
X1590 a_28714_19898# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15900 vcm_commonmode a_16362_18528# a_29414_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15901 VDD a_11067_67279# a_43378_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15902 vcm_commonmode a_16362_13508# a_30418_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15903 a_18674_63198# a_15439_49525# a_18278_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15904 VSS a_2595_47653# a_4761_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15905 a_2781_44655# a_1591_44655# a_2672_44655# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15906 a_46482_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15907 a_43378_61190# a_16362_61190# a_43470_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15908 a_36842_8456# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15909 a_14902_48783# a_5039_42167# a_14524_48437# VSS sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X1591 VDD a_33155_35839# a_33015_36161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15910 a_26310_71230# a_16362_71230# a_26402_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15911 a_32730_58178# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15912 VDD a_10055_58791# a_33338_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X15913 vcm_commonmode a_16362_66210# a_42466_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15914 a_38239_32375# a_36507_31573# a_38382_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15915 a_2467_28662# a_2216_28309# a_2008_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15916 a_9150_71311# a_9024_71427# a_8746_71443# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X15917 a_32310_49257# a_28108_48463# a_32218_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15918 VDD a_12343_36893# a_12369_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X15919 VDD a_12947_8725# a_46390_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1592 a_19678_9858# a_12985_19087# a_19282_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15920 VSS a_12985_19087# a_42770_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15921 a_44382_24918# VSS a_44474_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15922 a_1803_20719# a_1626_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X15923 a_47886_70548# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15924 a_4174_52854# a_3668_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X15925 a_44474_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15926 a_9613_48981# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15927 a_20378_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15928 a_2215_71311# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15929 a_44778_69222# a_12516_7093# a_44382_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1593 a_34613_31375# a_32970_31145# a_34395_31287# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X15930 a_47394_60186# a_16362_60186# a_47486_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15931 VSS a_12985_19087# a_18674_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15932 a_38239_32375# a_38210_30199# a_38299_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X15933 a_32426_63198# a_16746_63200# a_32334_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15934 VDD config_1_in[1] a_1591_9295# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X15935 VSS a_3143_22364# a_3529_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15936 VSS a_12707_26159# a_13251_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X15937 VSS a_12901_66665# a_23694_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15938 VDD a_12985_16367# a_37354_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15939 a_33045_49871# a_6831_63303# a_32318_48695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1594 a_30326_70226# a_16362_70226# a_30418_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15940 a_28714_8854# a_12947_8725# a_28318_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15941 a_25221_41281# a_24423_40229# a_25355_40183# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X15942 a_21382_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15943 VDD a_12901_66665# a_24302_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15944 a_17366_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15945 VDD a_3143_22364# a_4233_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15946 a_51422_39932# a_51714_39886# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X15947 VDD a_13669_39605# a_13613_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X15948 a_24394_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15949 a_48794_68218# a_12901_66959# a_48398_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1595 a_33830_13476# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15950 VSS a_12355_65103# a_45782_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15951 a_34639_42089# a_35033_42044# a_34699_42035# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X15952 vcm_commonmode a_16362_67214# a_19374_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15953 a_11017_16367# a_10973_16609# a_10851_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X15954 a_23390_65206# a_16746_65208# a_23298_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15955 vcm_commonmode a_16362_56170# a_49494_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15956 a_15305_38543# a_15039_38909# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15957 a_23535_50247# a_22989_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15958 a_11138_12267# a_11455_12157# a_11413_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15959 VSS a_23901_43132# a_23593_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1596 a_31726_9858# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X15960 a_22294_20902# a_16362_20536# a_22386_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15961 a_25447_43447# a_24515_43493# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15962 VDD a_12981_62313# a_32334_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15963 VSS a_12257_56623# a_35742_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15964 VDD a_3491_42239# a_3478_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X15965 VSS a_32181_36893# a_31873_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15966 VDD a_12355_15055# a_45386_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15967 a_37589_31393# a_32970_31145# a_37503_31393# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X15968 a_37446_11500# a_16746_11498# a_37354_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15969 VDD a_12727_13353# a_49402_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1597 VSS a_10975_66407# a_18674_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X15970 VSS a_14258_34191# a_18851_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X15971 vcm_commonmode a_16362_8488# a_34434_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X15972 a_26402_56170# a_16746_56172# a_26310_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15973 a_27710_17890# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15974 VDD a_12895_13967# a_36350_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15975 a_25798_7452# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15976 a_21686_7850# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15977 a_29545_28023# a_28963_28853# a_29708_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X15978 VSS a_12727_13353# a_31726_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15979 a_2672_23817# a_1757_23445# a_2325_23413# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1598 VDD a_4831_58497# a_4792_58371# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15980 a_35647_40229# a_33856_40743# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X15981 a_40762_63198# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15982 a_37354_68218# a_16362_68218# a_37446_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15983 a_44474_8488# a_16746_8486# a_44382_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15984 VDD a_4571_26677# a_7921_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15985 VDD a_15439_49525# a_18278_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15986 a_4163_12015# a_3327_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15987 a_9190_74941# a_8575_74853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15988 a_25299_30083# a_25263_29981# a_25227_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X15989 a_9945_47919# a_9779_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1599 a_31551_31751# a_31659_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X15990 a_31117_28879# a_30788_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15991 a_14293_41807# a_13867_42134# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15992 VSS a_29545_40193# a_29863_39913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X15993 VDD a_12135_69109# a_12093_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15994 a_8060_58799# a_8199_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15995 VSS a_38499_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X15996 VSS a_2011_34837# a_4263_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15997 result_out[12] a_1644_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X15998 a_32334_58178# a_10515_22671# a_32826_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X15999 a_7075_42479# a_6559_42479# a_6980_42479# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X16 a_17033_38565# a_16879_37999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X160 a_33641_29967# a_33363_30305# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X1600 a_9221_24847# a_7203_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X16000 VDD a_12727_67753# a_44382_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16001 a_32730_11866# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16002 a_2426_31421# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16003 a_24184_47741# a_7479_54439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16004 a_29322_10862# a_16362_10496# a_29414_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16005 a_2203_19631# a_1757_19631# a_2107_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16006 a_22213_37479# a_22521_37692# a_20827_37737# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X16007 a_19282_71230# a_12901_66665# a_19774_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16008 VSS a_2437_28309# a_2371_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16009 VDD a_2011_34837# a_4522_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1601 a_76365_40202# a_76461_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16010 a_44474_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16011 a_3357_22649# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16012 VSS a_12355_15055# a_30722_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16013 a_14001_28157# a_11902_27497# a_13919_27904# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16014 a_27406_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16015 a_29718_55166# VSS a_29322_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16016 VSS a_1923_59583# a_4365_64061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16017 a_44778_64202# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16018 a_7155_55509# a_7479_67075# a_7681_67279# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X16019 a_32795_44031# a_31004_44869# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X1602 VDD a_2163_73085# a_2124_73211# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X16020 a_44778_22910# a_11067_21583# a_44382_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16021 a_5064_65327# a_4149_65327# a_4717_65569# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16022 a_42374_21906# a_11067_21583# a_42866_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16023 a_42374_17890# a_16362_17524# a_42466_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16024 VDD a_40403_37683# a_40429_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X16025 a_9263_24501# a_7377_18012# a_9959_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X16026 a_22793_51005# a_22749_50613# a_22627_51017# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16027 a_17366_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16028 VDD VSS a_31330_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16029 a_34738_56170# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1603 a_22690_64202# a_12355_65103# a_22294_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16030 vcm_commonmode a_16362_58178# a_26402_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16031 a_17670_66210# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16032 a_4220_57685# a_4674_57685# a_4612_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X16033 a_3595_37583# a_2971_37589# a_3487_37961# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X16034 VSS a_7815_42453# a_7749_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16035 VSS a_11067_13095# a_21686_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16036 a_35838_55488# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16037 a_48890_15484# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16038 a_45386_12870# a_12877_16911# a_45878_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16039 a_48794_21906# a_12985_7663# a_48398_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1604 VDD VSS a_36350_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16040 vcm_commonmode a_16362_20536# a_19374_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16041 a_3280_70501# a_1586_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X16042 a_22294_65206# a_16362_65206# a_22386_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16043 a_1761_2767# a_1591_2767# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16044 a_28318_22910# a_10515_23975# a_28810_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16045 a_9305_53511# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16046 a_34434_61190# a_16746_61192# a_34342_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16047 a_18278_55166# VSS a_18370_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16048 vcm_commonmode VSS a_23390_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16049 a_32826_20504# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1605 a_16362_19532# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X16050 a_32426_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16051 VDD a_24667_31055# a_24746_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16052 a_3484_61493# a_3938_61493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16053 a_17366_71230# a_16746_71232# a_17274_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16054 a_38754_13874# a_12877_16911# a_38358_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16055 VSS a_12985_16367# a_35742_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16056 a_41351_42405# a_40585_42369# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16057 vcm_commonmode VSS a_45478_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16058 a_18278_14878# a_12877_14441# a_18770_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16059 VDD a_7862_34025# a_26311_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1606 a_20778_72556# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16060 VSS a_18539_47617# a_18500_47491# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16061 a_19282_18894# a_16362_18528# a_19374_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16062 VDD a_12877_14441# a_25306_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16063 a_22786_12472# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16064 a_49402_11866# a_10055_58791# a_49894_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16065 a_20286_13874# a_16362_13508# a_20378_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16066 a_39362_68218# a_12727_67753# a_39854_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16067 a_43530_28585# a_43495_28487# a_43227_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16068 a_43870_66532# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16069 a_40366_63198# a_12981_62313# a_40858_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1607 a_46882_12472# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16070 a_43378_9858# a_12546_22351# a_43870_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16071 VSS a_3173_46805# a_3107_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16072 a_38450_60186# a_16746_60188# a_38358_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16073 a_38450_19532# a_16746_19530# a_38358_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16074 VDD a_26889_50337# a_26779_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16075 vcm_commonmode a_16362_16520# a_35438_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16076 a_33338_12870# a_16362_12504# a_33430_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16077 a_33008_28853# a_30788_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X16078 VDD a_20713_39105# a_22260_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16079 a_17008_49007# a_16891_49220# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1608 VDD a_1586_40455# a_1591_49557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X16080 a_9669_26703# a_9289_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X16081 VSS a_32031_37683# a_31971_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16082 VSS a_33264_37601# a_33727_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X16083 a_12447_29199# a_13353_30511# a_18944_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16084 a_19282_9858# a_12546_22351# a_19774_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16085 a_5639_27247# a_3972_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16086 vcm_commonmode a_16362_15516# a_48490_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16087 a_22386_24552# VDD a_22294_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16088 a_19621_52521# a_19576_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16089 a_9135_25321# a_6162_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 VDD a_12985_7663# a_20286_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16090 a_17709_48761# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16091 a_35438_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16092 a_26802_11468# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16093 a_2672_23817# a_1591_23445# a_2325_23413# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16094 VSS a_39836_38567# a_39449_39868# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X16095 a_29814_9460# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16096 VDD a_2417_31841# a_2307_31965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16097 VDD a_12983_63151# a_20286_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16098 a_44382_62194# a_12355_15055# a_44874_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16099 a_1954_61677# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X161 a_37750_61190# a_12355_15055# a_37354_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1610 VDD a_10975_66407# a_19282_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16100 VDD a_7479_57175# a_6515_62037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16101 a_10391_67477# a_10216_67503# a_10570_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16102 a_30412_34337# a_29943_34789# a_30816_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16103 a_33080_37149# a_32795_36415# a_33727_36649# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16104 VSS a_5993_32687# a_7295_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16105 a_25398_15516# a_16746_15514# a_25306_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16106 a_48398_19898# a_11067_67279# a_48890_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16107 a_32730_72234# VDD a_32334_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16108 a_12651_41085# a_12663_40871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16109 a_17274_64202# a_11067_13095# a_17766_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1611 a_44382_13874# a_16362_13508# a_44474_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16110 a_1586_40455# a_4535_43031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16111 a_21782_62516# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16112 a_2867_15279# a_2830_15431# a_1895_14906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16113 a_22169_52093# a_19478_51959# a_22097_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16114 a_31726_58178# a_12901_58799# a_31330_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16115 a_45782_71230# a_12947_71576# a_45386_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16116 VDD a_3805_30083# a_4248_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16117 a_40458_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16118 a_29414_14512# a_16746_14510# a_29322_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16119 a_18907_48502# a_18413_47919# a_18835_48502# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1612 a_1757_26159# a_1591_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16120 vcm_commonmode a_16362_11500# a_26402_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16121 a_6989_24233# a_5531_22895# a_6917_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16122 a_25798_19500# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16123 a_11433_69921# a_11215_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X16124 a_27415_36341# a_12473_37429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16125 a_25015_48437# a_25019_47679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16126 a_2409_72399# a_2322_72631# a_1895_71482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16127 VDD a_12257_56623# a_27314_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16128 VDD a_6393_34837# a_6423_35190# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16129 VDD a_34759_31029# a_38209_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1613 VDD a_26020_30199# a_25971_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X16130 a_12671_41807# a_12417_42134# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16131 a_6369_74031# a_5179_74031# a_6260_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X16132 vcm_commonmode a_16362_64202# a_38450_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16133 a_16154_42134# a_15459_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X16134 VSS a_7467_61751# a_3938_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16135 a_5489_69135# a_4345_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16136 a_43774_23914# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16137 a_44474_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16138 a_7681_67279# a_3143_66972# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16139 a_2163_54589# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1614 a_23390_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16140 a_9613_13077# a_1929_12131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16141 a_21231_30511# a_20911_31055# a_21123_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16142 a_20286_58178# a_16362_58178# a_20378_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16143 a_34342_71230# a_16362_71230# a_34434_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16144 VSS a_12895_13967# a_36746_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16145 a_32121_44545# a_32795_44031# a_33668_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16146 a_10229_66237# a_2840_66103# a_10147_65984# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16147 a_40762_16886# a_12727_13353# a_40366_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16148 a_5970_43567# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16149 a_20282_49551# a_20195_49793# a_19878_49683# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X1615 a_29814_22512# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16150 a_33338_57174# a_16362_57174# a_33430_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16151 VSS a_12899_10927# a_49798_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16152 a_20286_17890# a_12899_10927# a_20778_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16153 VSS a_12947_23413# a_20682_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16154 VDD a_7755_54999# a_7210_55081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16155 a_17366_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16156 a_8583_22671# a_4798_23759# a_8671_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16157 VSS a_4903_31849# a_10317_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16158 a_36831_49257# a_28881_52271# a_36735_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16159 a_10614_53942# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1616 a_20286_62194# a_16362_62194# a_20378_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16160 VSS a_32370_50871# a_32091_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16161 VSS a_9011_74879# a_8945_74953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16162 a_41862_59504# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16163 a_48398_7850# VDD a_48890_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16164 a_37750_14878# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16165 a_3749_37949# a_3705_37557# a_3583_37961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16166 VSS a_2606_41079# a_19128_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16167 vcm_commonmode a_16362_70226# a_20378_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16168 a_8994_63927# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X16169 a_32672_49007# a_32135_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X1617 a_28817_28111# a_13643_28327# a_28599_28023# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16170 a_17654_51183# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16171 a_26706_17890# a_12899_11471# a_26310_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16172 VSS a_13143_29575# a_13643_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16173 VDD a_2672_21807# a_2847_21781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16174 VSS a_1950_59887# a_10147_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X16175 VDD a_12901_66665# a_32334_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16176 a_24302_16886# a_12899_11471# a_24794_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16177 a_49750_39288# a_42165_36367# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.394e+11p pd=2.82e+06u as=0p ps=0u w=420000u l=150000u M=2
X16178 a_1950_59887# a_1920_59861# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X16179 a_1761_35951# a_1591_35951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1618 a_41766_67214# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16180 a_12815_16519# a_12580_15939# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X16181 VSS a_10317_67191# a_10010_68021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16182 a_12641_43124# a_12671_42134# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16183 a_4993_32929# a_4775_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X16184 vcm_commonmode a_16362_61190# a_23390_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16185 VDD a_41211_28023# a_39727_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X16186 VDD a_20009_48981# a_20039_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16187 VDD a_12901_58799# a_31330_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16188 VDD a_1923_54591# a_9187_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16189 VSS a_12727_15529# a_27710_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1619 VSS a_6738_19783# a_6743_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X16190 a_11644_30761# a_10899_28879# a_11183_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16191 a_31726_11866# a_12985_16367# a_31330_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16192 VDD a_29927_29199# a_36401_46859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16193 VDD a_12947_71576# a_18278_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16194 a_21627_49373# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16195 VDD a_7563_46261# a_7494_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16196 a_77285_40202# a_77381_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16197 a_12341_3311# a_12171_3311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16198 VDD VDD a_35346_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16199 a_2939_31573# a_2764_31599# a_3118_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X162 a_4831_58497# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1620 a_19374_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16200 a_18370_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16201 VSS a_10975_66407# a_39758_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16202 a_32334_66210# a_10975_66407# a_32826_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16203 VSS a_2191_68565# a_4075_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16204 a_43774_64202# a_12355_65103# a_43378_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16205 vcm_commonmode a_16362_60186# a_27406_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16206 vcm_commonmode a_16362_19532# a_27406_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16207 a_37846_23516# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16208 a_2989_45717# a_2656_45895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16209 a_37446_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1621 a_7458_10515# a_7736_10499# a_7692_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16210 VSS a_1586_45431# a_4535_43031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16211 VDD a_12985_7663# a_41370_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16212 a_41766_7850# VDD a_41370_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16213 VDD a_7155_55509# a_6646_54135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16214 a_30139_36649# a_29207_36415# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16215 a_44474_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16216 a_41370_62194# a_16362_62194# a_41462_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16217 a_4032_53047# a_1823_53885# a_4174_52854# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X16218 a_1761_27791# a_1591_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16219 VDD a_38327_44759# a_38140_44501# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1622 a_2203_23817# a_1757_23445# a_2107_23817# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X16220 a_36199_32143# a_35815_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16221 a_33734_56170# a_12257_56623# a_33338_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16222 a_29718_63198# a_15439_49525# a_29322_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16223 a_17670_7850# VDD a_17274_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16224 VSS a_23447_28853# a_23298_28487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16225 a_44778_72234# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16226 vcm_commonmode a_16362_67214# a_40458_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16227 a_9613_13077# a_1929_12131# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16228 VDD a_11763_21237# a_11480_23957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16229 a_12885_37782# a_12343_36893# a_12671_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1623 a_33338_61190# a_16362_61190# a_33430_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X16230 VSS a_12546_22351# a_22690_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16231 a_2847_26133# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16232 VSS a_28441_36389# a_29127_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X16233 a_38358_15882# a_16362_15516# a_38450_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16234 VDD a_2787_32679# a_7942_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.5e+11p ps=2.7e+06u w=1e+06u l=150000u
X16235 a_2058_34102# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16236 VDD a_10055_58791# a_44382_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16237 a_8543_36469# a_5363_30503# a_8762_36815# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16238 a_42466_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16239 VDD a_31223_36369# a_31083_36395# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1624 a_36746_10862# a_12546_22351# a_36350_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16240 VDD a_14963_39783# a_19417_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X16241 a_2965_47753# a_1775_47381# a_2856_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X16242 a_9972_69831# a_1586_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16243 a_8449_43361# a_8383_43255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16244 a_37750_55166# VSS a_37354_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16245 VSS VDD a_21686_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16246 a_18703_29199# a_33694_30761# a_42715_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X16247 a_2847_40277# a_2672_40303# a_3026_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16248 a_48490_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16249 a_14076_35077# a_13107_34789# a_13980_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X1625 a_4887_36495# a_4443_36611# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16250 a_2121_56623# a_1643_56597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16251 a_15681_27497# a_11430_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16252 a_33864_28111# a_25787_28327# a_33689_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X16253 a_30418_66210# a_16746_66212# a_30326_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16254 VDD a_12985_16367# a_48398_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16255 a_7561_36495# a_5915_35943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16256 a_3026_69501# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16257 a_8289_52047# a_4298_58951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16258 VDD a_12901_66959# a_38358_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16259 a_18278_63198# a_16362_63198# a_18370_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1626 a_25263_39913# a_25300_39655# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X16260 a_32426_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16261 VDD a_14298_32143# a_8491_41383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16262 a_12815_53609# a_4351_67279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16263 vcm_commonmode a_16362_58178# a_34434_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16264 a_19374_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16265 a_13835_36649# a_15775_36965# a_16707_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16266 vcm_commonmode a_16362_68218# a_17366_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16267 VSS a_16152_43677# a_15253_43421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X16268 vcm_commonmode a_16362_57174# a_47486_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16269 VSS a_2959_47113# a_35039_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1627 VDD a_9653_69831# a_9466_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16270 VSS a_30412_34337# a_30875_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16271 VSS a_18045_41281# a_18915_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16272 a_33430_7484# VDD a_33338_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16273 a_11851_64391# a_11521_66567# a_12085_64239# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16274 VSS a_2143_15271# a_11711_12559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16275 a_40366_71230# a_12901_66665# a_40858_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16276 a_39854_64524# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16277 a_36350_61190# a_12981_59343# a_36842_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16278 a_33338_20902# a_16362_20536# a_33430_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16279 VSS a_76365_39738# a_76178_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1628 vcm_commonmode a_16362_21540# a_43470_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16280 a_77922_40050# a_75475_38962# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16281 VDD a_12981_62313# a_43378_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16282 a_4057_50645# a_3891_50645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X16283 a_2882_56989# a_2163_56765# a_2319_56860# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16284 VSS a_12355_15055# a_28714_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16285 VDD a_11709_61217# a_11599_61341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16286 a_24394_57174# a_16746_57176# a_24302_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16287 a_25702_18894# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16288 a_5051_43567# a_4535_43567# a_4956_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16289 a_1644_58773# a_1823_58773# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1629 a_46482_24552# VDD a_46390_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16290 a_12877_14441# a_11067_13095# a_12723_14191# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16291 VSS a_2744_46983# a_2467_47893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16292 a_7171_45577# a_6725_45205# a_7075_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16293 a_24394_9492# a_16746_9490# a_24302_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16294 a_44382_70226# a_12516_7093# a_44874_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16295 a_16648_42693# a_15775_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16296 a_48398_68218# a_16362_68218# a_48490_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16297 VSS a_12901_66959# a_41766_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16298 a_5239_20693# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16299 VDD a_15439_49525# a_29322_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X163 a_32730_7850# VDD a_32334_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1630 a_19774_14480# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16300 a_6737_27907# a_5085_23047# a_6641_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16301 VSS a_5085_23047# a_6559_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16302 a_30326_59182# a_12901_58799# a_30818_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16303 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16304 a_26225_47919# a_4891_47388# a_25879_48169# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16305 a_27683_52271# a_27333_52271# a_27588_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X16306 VSS a_4528_26159# a_7203_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16307 VSS a_2011_34837# a_4762_35484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16308 a_8074_38991# a_5363_30503# a_7755_38991# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u w=650000u l=150000u
X16309 VDD a_13669_38517# a_13613_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1631 a_19678_20902# a_11067_67279# a_19282_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16310 a_17274_72234# VDD a_17766_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16311 vcm_commonmode a_16362_20536# a_40458_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16312 a_43470_23548# a_16746_23546# a_43378_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16313 a_18977_28111# a_18126_28023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16314 VSS a_39468_37479# a_39431_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X16315 a_21782_70548# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16316 a_42466_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16317 VDD a_1761_34319# a_33155_35839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16318 a_17766_60508# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16319 a_25398_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1632 a_17274_15882# a_16362_15516# a_17366_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16320 VSS a_2689_65103# a_4119_70741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X16321 VDD a_37520_49783# a_36464_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X16322 VDD a_2325_51425# a_2215_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16323 a_5353_43343# a_3987_19623# a_4842_45467# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16324 a_6913_72399# a_6559_72512# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16325 a_42770_65206# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16326 VSS a_23901_42044# a_23593_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16327 a_33430_15516# a_16746_15514# a_33338_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16328 VSS a_29207_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X16329 a_16746_71232# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X1633 VDD a_10055_58791# a_23298_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16330 a_42866_17492# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16331 a_31422_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16332 a_40366_18894# a_16362_18528# a_40458_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16333 a_5052_14709# a_5755_14709# a_5709_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16334 VDD a_8575_74853# a_8459_71285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16335 VSS a_1586_18695# a_1591_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16336 a_2744_53511# a_2952_53333# a_2886_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16337 vcm_commonmode VSS a_38450_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16338 a_8355_18870# a_8104_18517# a_7896_18695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16339 a_7939_27497# a_6773_27805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1634 vcm_commonmode a_16362_66210# a_32426_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16340 a_42466_70226# a_16746_70228# a_42374_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16341 a_22690_68218# a_12901_66959# a_22294_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16342 VSS a_12901_58799# a_48794_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16343 a_45782_56170# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16344 a_37354_9858# a_16362_9492# a_37446_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16345 vcm_commonmode a_16362_11500# a_34434_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16346 a_46882_16488# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16347 a_43378_13874# a_12727_15529# a_43870_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16348 a_28714_66210# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16349 VSS a_11067_13095# a_32730_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1635 a_21382_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16350 a_4433_55581# a_3295_62083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16351 a_33830_19500# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16352 vcm_commonmode a_16362_21540# a_17366_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16353 a_26310_23914# a_12947_23413# a_26802_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16354 vcm_commonmode a_16362_10496# a_47486_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16355 a_26310_19898# a_16362_19532# a_26402_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16356 a_47486_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16357 a_30818_21508# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16358 a_30418_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16359 a_14945_37479# a_15253_37692# a_14919_37683# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1636 a_28318_7850# VSS a_28410_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16360 a_4345_69679# a_2952_66139# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16361 VSS a_40457_27765# a_40402_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X16362 a_7369_24233# a_6989_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X16363 VSS a_19885_50095# a_20914_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16364 a_20267_30503# a_33694_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X16365 a_33338_65206# a_16362_65206# a_33430_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X16366 a_36746_14878# a_12727_15529# a_36350_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16367 a_7407_18038# a_6816_19355# a_7407_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16368 a_45478_61190# a_16746_61192# a_45386_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16369 a_25702_59182# a_12727_58255# a_25306_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1637 a_21267_52047# a_19478_51959# a_21178_52047# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X16370 VSS a_12947_56817# a_22690_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16371 a_49798_55166# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16372 a_19774_18496# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16373 a_19678_24918# VSS a_19282_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16374 VDD a_12727_13353# a_23298_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16375 a_49798_13874# a_12877_16911# a_49402_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16376 a_20778_13476# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16377 VDD a_11902_27497# a_19525_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16378 a_7755_23145# a_4528_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16379 a_37354_69222# a_12901_66959# a_37846_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1638 a_9863_51420# a_9668_51451# a_10173_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X16380 VSS a_10883_11177# a_11898_10205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16381 a_41862_67536# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16382 a_24394_10496# a_16746_10494# a_24302_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16383 VDD a_3799_31063# a_2473_34293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16384 VSS a_8005_53333# a_2952_53333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X16385 VSS a_35676_49525# a_37512_50755# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16386 a_31330_13874# a_16362_13508# a_31422_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16387 a_32795_42943# a_31648_43781# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X16388 a_49494_60186# a_16746_60188# a_49402_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16389 vcm_commonmode a_16362_16520# a_46482_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1639 a_41862_63520# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16390 a_49494_19532# a_16746_19530# a_49402_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16391 VDD a_6473_40277# a_6417_40630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X16392 a_24302_67214# a_16362_67214# a_24394_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16393 VSS VSS a_26706_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16394 a_39305_32463# a_12907_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16395 a_10244_26159# a_6162_28487# a_10138_26159# VSS sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X16396 a_6614_47919# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16397 VSS a_10515_23975# a_41766_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16398 a_38450_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16399 a_25939_51157# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X164 VSS a_12899_10927# a_34738_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1640 VSS a_17488_48731# a_18430_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X16400 a_27806_68540# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16401 VSS a_13669_38517# a_13613_38870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16402 a_13809_48463# a_13461_48579# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X16403 a_33597_48829# a_32672_49007# a_33515_48576# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16404 a_6800_20291# a_5825_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16405 VDD a_12983_63151# a_31330_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16406 VDD a_27652_38237# a_26753_37981# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X16407 a_24844_47753# a_23929_47381# a_24497_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X16408 VSS a_1586_69367# a_2971_73493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16409 a_31422_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1641 a_36442_16520# a_16746_16518# a_36350_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16410 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16411 a_25300_39655# a_24331_39679# a_25204_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16412 a_45782_9858# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16413 a_48890_57496# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16414 a_36746_71230# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16415 a_35438_69222# a_16746_69224# a_35346_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16416 a_43774_72234# VDD a_43378_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16417 VDD a_7499_74031# a_7901_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16418 a_28318_64202# a_11067_13095# a_28810_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16419 a_2108_10749# a_1761_9295# a_1887_10422# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1642 a_45878_18496# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16420 VDD a_5535_18012# a_12360_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16421 a_32826_62516# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16422 a_16012_41959# a_15931_39859# a_16154_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X16423 a_6641_63401# a_2927_68565# a_6559_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16424 a_8857_14709# a_8639_15113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X16425 VSS a_2847_69439# a_2781_69513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X16426 VSS a_8325_18517# a_8259_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16427 VSS a_12947_23413# a_18674_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16428 VDD a_1923_73087# a_3588_70589# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16429 VSS a_12877_16911# a_48794_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1643 a_41510_29673# a_28757_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X16430 a_22690_21906# a_12985_7663# a_22294_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16431 a_38436_29941# a_32823_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X16432 a_18278_56170# a_12947_56817# a_18770_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16433 a_30599_28023# a_12907_27023# a_30745_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X16434 a_44177_28879# a_41842_27221# a_43495_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16435 a_17321_49249# a_17103_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X16436 VDD a_10515_22671# a_25306_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16437 a_39454_68218# a_16746_68220# a_39362_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16438 vcm_commonmode a_16362_65206# a_36442_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16439 VDD a_4036_54421# a_3295_54421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X1644 a_4032_53047# a_4240_53083# a_4174_53181# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16440 VSS a_31171_27412# a_29760_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X16441 a_41766_24918# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16442 a_38358_23914# a_16362_23548# a_38450_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16443 a_7933_51433# a_7073_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16444 VDD a_4972_51017# a_5147_50943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16445 a_30722_69222# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16446 VDD a_27195_32375# a_27167_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16447 a_33385_46805# a_22291_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16448 a_22176_47919# a_21261_47919# a_21829_48161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16449 a_25702_12870# a_10055_58791# a_25306_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1645 vcm_commonmode VSS a_42466_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16450 a_37750_63198# a_15439_49525# a_37354_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16451 a_1929_10651# a_2847_9813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16452 a_32730_9858# a_12985_19087# a_32334_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16453 VSS a_12727_58255# a_34738_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16454 VDD a_77002_39738# a_76744_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16455 a_10472_54135# a_10680_52245# a_10614_53942# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16456 VSS a_11067_67279# a_34738_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16457 vcm_commonmode a_16362_23548# a_32426_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16458 VDD a_14293_39631# a_19769_38793# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X16459 VSS a_12516_7093# a_17670_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1646 VSS a_11067_23759# a_16362_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X16460 VSS a_40403_37683# a_40343_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16461 a_23685_38341# a_23993_37981# a_23565_38565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X16462 a_31330_58178# a_16362_58178# a_31422_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16463 a_45386_71230# a_16362_71230# a_45478_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16464 VSS a_12895_13967# a_47790_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16465 a_30657_29967# a_30052_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16466 a_16955_52047# a_12907_27023# a_37922_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16467 a_11877_50645# a_11711_50645# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16468 a_1849_52271# a_1683_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16469 VDD a_10391_67477# a_10378_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1647 VSS a_35517_34954# a_26550_40871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X16470 vcm_commonmode a_16362_15516# a_22386_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16471 VDD a_11067_21583# a_35346_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16472 a_31330_17890# a_12899_10927# a_31822_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16473 VSS a_4311_58229# a_1823_65853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16474 a_4031_73095# a_2686_70223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16475 VSS a_6473_40277# a_6417_40630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16476 VSS a_21187_29415# a_32401_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16477 VSS a_10649_58947# a_10607_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X16478 a_28318_8854# a_12985_19087# a_28810_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16479 a_20972_28335# a_20027_27221# a_5915_35943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X1648 a_49494_15516# a_16746_15514# a_49402_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16480 a_7821_22057# a_4571_26677# a_7749_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16481 a_35487_49871# a_28881_52271# a_35379_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16482 VDD a_2216_28309# a_4095_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16483 vcm_commonmode a_16362_9492# a_47486_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16484 a_22386_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16485 a_49402_70226# a_16362_70226# a_49494_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16486 a_24698_18894# a_12899_10927# a_24302_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16487 a_48794_14878# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16488 vcm_commonmode a_16362_70226# a_31422_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16489 a_27214_28335# a_3339_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1649 vcm_commonmode a_16362_12504# a_46482_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16490 a_39854_72556# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16491 a_19121_48502# a_4482_57863# a_18907_48502# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X16492 VDD a_12901_66665# a_43378_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16493 a_36442_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16494 VDD a_12981_59343# a_39362_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16495 a_39362_62194# a_16362_62194# a_39454_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16496 a_11763_20407# a_3987_19623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X16497 a_22294_19898# a_11067_67279# a_22786_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16498 vcm_commonmode a_16362_62194# a_21382_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16499 a_43470_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X165 VDD a_4427_25071# a_5918_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.25e+11p ps=2.45e+06u w=1e+06u l=150000u
X1650 a_20378_21540# a_16746_21538# a_20286_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16500 VSS a_1954_61677# a_3983_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16501 VSS a_33593_31287# a_32367_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16502 a_11945_23777# a_11480_23957# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16503 a_7987_15431# a_9275_15253# a_9221_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16504 a_26402_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16505 a_7192_58255# a_7107_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16506 a_9835_69513# a_9485_69141# a_9740_69501# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X16507 a_8938_61519# a_7210_55081# a_8635_61751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16508 VSS a_12877_14441# a_25702_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16509 a_1761_34319# a_1591_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1651 a_35438_9492# a_16746_9490# a_35346_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16510 result_out[2] a_1644_56053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16511 VDD a_10103_11079# a_9455_11079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16512 a_35438_22544# a_16746_22542# a_35346_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16513 VDD a_11430_26159# a_14482_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.55e+11p ps=5.31e+06u w=1e+06u l=150000u
X16514 VDD VDD a_16270_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16515 VSS a_21879_30663# a_21057_30669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X16516 VDD a_7213_62215# a_7539_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16517 a_26523_29199# a_2787_30503# a_27132_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16518 VDD a_29667_31055# a_30203_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X16519 VDD a_13576_42589# a_12677_42333# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X1652 a_5235_71855# a_4719_71855# a_5140_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X16520 VDD a_12947_71576# a_29322_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16521 VSS a_12983_63151# a_37750_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16522 VDD a_20827_37737# a_22213_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16523 a_26778_29473# a_26191_29397# a_26694_29473# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16524 VSS a_29513_34428# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X16525 a_30326_67214# a_12983_63151# a_30818_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16526 a_41766_65206# a_10975_66407# a_41370_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16527 a_3541_19385# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16528 VDD a_12473_37429# a_12885_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16529 VSS a_76365_40202# a_76178_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1653 a_35742_58178# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16530 a_29414_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16531 a_21686_8854# a_12947_8725# a_21290_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16532 VSS a_22448_39429# a_22411_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16533 VDD a_2223_28617# a_3186_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16534 a_39454_21540# a_16746_21538# a_39362_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16535 a_27183_40229# a_26417_40193# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X16536 a_28410_66210# a_16746_66212# a_28318_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16537 a_12680_53511# a_12953_53339# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16538 VDD a_1952_60431# a_4441_62327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16539 a_14049_40693# a_13067_38517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1654 VDD a_12985_16367# a_27314_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16540 a_30722_22910# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16541 a_5081_34025# a_4893_33821# a_4999_33781# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16542 a_27314_21906# a_16362_21540# a_27406_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16543 a_2847_19605# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16544 VDD a_15439_49525# a_37354_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16545 VSS a_9751_25071# a_12263_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16546 a_44778_56170# a_12257_56623# a_44382_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16547 a_27323_30083# a_25321_29673# a_27251_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16548 VSS a_12899_10927# a_23694_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16549 VSS a_4149_24527# a_5449_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1655 VDD a_2847_18517# a_3325_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16550 a_10053_69109# a_9835_69513# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X16551 a_4057_13647# a_3677_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16552 a_9359_60214# a_9177_60214# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16553 VDD a_37459_51183# a_37534_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X16554 VSS a_8399_49159# a_8399_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X16555 a_33430_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16556 a_6340_61225# a_2952_66139# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16557 a_2882_59343# a_2124_59459# a_2319_59317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16558 vcm_commonmode a_16362_59182# a_41462_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16559 VDD a_2325_23413# a_2215_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1656 VSS a_4333_22895# a_4903_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X16560 a_35550_27791# a_21187_29415# a_35478_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X16561 a_35647_38053# a_32031_37683# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16562 a_46482_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16563 VSS VDD a_32730_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16564 VSS a_6435_47893# a_6369_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16565 VSS a_14511_50069# a_14445_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16566 a_3417_33231# a_2939_33535# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16567 VDD a_12516_7093# a_36350_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16568 a_35676_49525# a_29361_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16569 a_24698_13874# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1657 VDD a_12901_66959# a_17274_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16570 a_3019_46070# a_2539_42106# a_2560_45895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16571 a_3339_30503# a_24768_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16572 a_5064_65327# a_3983_65327# a_4717_65569# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16573 a_36442_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16574 a_6260_47919# a_5179_47919# a_5913_48161# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16575 VDD a_12901_66959# a_49402_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16576 a_49798_63198# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16577 a_12481_54447# a_12203_54475# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X16578 a_19374_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16579 vcm_commonmode a_16362_58178# a_45478_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1658 a_3541_9593# a_1689_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16580 a_2012_40303# a_1895_40516# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16581 vcm_commonmode a_16362_68218# a_28410_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16582 a_34342_23914# a_12947_23413# a_34834_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16583 a_10073_23439# a_8569_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16584 a_22411_36919# a_21479_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16585 a_34342_19898# a_16362_19532# a_34434_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16586 a_17507_52047# a_37427_47893# a_37195_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16587 a_37846_65528# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16588 a_8569_49007# a_8399_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16589 a_32371_32117# a_32367_28309# a_32802_32463# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X1659 a_18674_68218# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16590 a_47394_22910# a_10515_23975# a_47886_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16591 a_37354_55166# VSS a_37446_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16592 VSS a_12981_62313# a_26706_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16593 VSS a_28789_50613# a_19478_51959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X16594 a_23694_60186# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16595 a_22386_58178# a_16746_58180# a_22294_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16596 a_36442_71230# a_16746_71232# a_36350_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16597 a_23694_19898# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16598 a_5089_53903# a_3325_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16599 VDD a_28639_49551# a_28814_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X166 a_7640_42479# a_6559_42479# a_7293_42721# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X1660 a_12899_3855# a_11067_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X16600 a_37354_14878# a_12877_14441# a_37846_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16601 VSS a_12985_7663# a_37750_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16602 a_8177_38991# a_3949_41935# a_8074_38991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16603 a_41862_12472# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16604 a_8201_62839# a_7803_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X16605 VSS a_1923_73087# a_5957_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16606 VDD a_5535_18012# a_12066_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X16607 VSS a_12473_37429# a_12892_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16608 a_24794_22512# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16609 VSS a_23731_28023# a_23051_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1661 a_7622_57711# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X16610 a_31422_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16611 a_19770_51005# a_2872_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16612 a_41462_24552# VDD a_41370_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16613 VDD a_12899_11471# a_17274_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16614 VDD a_9963_29967# a_10506_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X16615 a_13005_35823# a_12579_35862# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16616 a_2672_18543# a_1591_18543# a_2325_18785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16617 a_28318_72234# VDD a_28810_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16618 a_39758_70226# a_12901_66665# a_39362_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16619 a_28810_21508# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1662 a_35463_42943# a_33856_42693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16620 a_28410_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16621 VSS a_33264_37601# a_32365_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X16622 a_32826_70548# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16623 a_25306_14878# a_16362_14512# a_25398_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16624 VDD a_8367_44343# a_8308_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X16625 a_40858_18496# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16626 a_4312_19061# a_1586_18695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X16627 VDD a_31543_51335# a_30947_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16628 a_5175_27791# a_4995_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16629 a_32334_60186# a_16362_60186# a_32426_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1663 a_48794_57174# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16630 VDD a_30625_52245# a_30573_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16631 a_44474_15516# a_16746_15514# a_44382_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16632 vcm_commonmode a_16362_12504# a_41462_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16633 a_18770_13476# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16634 VSS a_10475_14165# a_9083_13879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16635 VDD a_12985_16367# a_22294_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16636 VDD a_4792_20443# a_10401_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16637 a_4771_56597# a_4974_56875# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16638 a_31096_38341# a_30127_38053# a_31059_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16639 a_33603_47081# a_26523_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1664 a_2713_35925# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16640 VDD a_42188_37149# a_42224_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16641 a_43774_57174# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16642 a_29322_13874# a_16362_13508# a_29414_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16643 a_26706_67214# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16644 a_49402_63198# a_12981_62313# a_49894_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16645 a_17366_17524# a_16746_17522# a_17274_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16646 VSS a_12355_65103# a_30722_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16647 a_1823_67668# a_1915_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16648 a_16746_68220# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X16649 a_48490_14512# a_16746_14510# a_48398_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1665 a_28410_7484# VDD a_28318_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16650 vcm_commonmode a_16362_11500# a_45478_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16651 a_21663_42943# a_20897_42917# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X16652 a_11659_66567# a_12231_65301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16653 a_22786_9460# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16654 a_44874_19500# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16655 vcm_commonmode a_16362_21540# a_28410_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16656 VSS a_4495_35925# a_4903_31849# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16657 a_28248_52271# a_27167_52271# a_27901_52513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16658 a_8031_24527# a_4351_26703# a_8113_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X16659 a_6567_25615# a_5085_24759# a_6649_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X1666 a_40858_69544# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16660 VSS a_12257_56623# a_20682_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16661 VSS a_23567_44211# a_23507_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16662 a_26802_63520# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16663 VSS a_5105_47673# a_5039_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16664 vcm_commonmode a_16362_13508# a_18370_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16665 VDD a_12355_15055# a_30326_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16666 a_11964_18543# a_10883_18543# a_11617_18785# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16667 a_22386_11500# a_16746_11498# a_22294_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16668 a_8080_47607# a_6559_22671# a_8222_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X16669 a_48398_69222# a_12901_66959# a_48890_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1667 a_35438_63198# a_16746_63200# a_35346_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16670 VDD a_12895_13967# a_21290_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16671 VSS a_1586_9991# a_3247_10389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16672 VDD a_30007_38695# a_13669_39605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X16673 a_3854_29977# a_2216_28309# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16674 a_17709_48761# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16675 a_22294_68218# a_16362_68218# a_22386_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16676 a_13795_35606# a_13613_35606# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16677 a_5629_21379# a_2317_28892# a_5547_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16678 a_28747_37503# a_27981_37477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16679 a_34434_64202# a_16746_64204# a_34342_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1668 a_30412_34337# a_29943_34789# a_30875_34743# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X16680 a_5993_32687# a_5515_32661# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16681 a_38850_8456# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16682 a_34738_8854# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16683 a_11711_28111# a_9179_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16684 a_36442_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16685 VDD a_13975_34191# a_14081_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16686 VDD a_30762_49641# a_30809_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X16687 VDD a_1643_64213# a_1591_64239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16688 a_10073_23439# a_9263_24501# a_10253_23759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X16689 VSS a_10751_59575# a_10649_58947# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1669 vcm_commonmode a_16362_9492# a_33430_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16690 a_13516_29673# a_10899_28879# a_13173_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16691 VDD a_12947_8725# a_48398_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16692 VSS a_12985_19087# a_44778_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16693 a_49494_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16694 a_25798_69544# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16695 VDD a_15607_46805# a_40599_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16696 a_32560_27907# a_21187_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16697 a_32730_18894# a_12899_10927# a_32334_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16698 VDD a_2319_64476# a_2250_64605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X16699 a_20505_29967# a_20103_30287# a_20341_30287# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X167 vcm_commonmode VSS a_44474_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1670 a_6260_10927# a_5345_10927# a_5913_11169# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X16700 VDD config_2_in[10] a_1591_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X16701 a_25306_59182# a_16362_59182# a_25398_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16702 VDD a_27891_41495# a_23789_39100# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X16703 a_18811_38053# a_18045_38017# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16704 a_39758_24918# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16705 VSS a_9642_10357# a_9583_10703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16706 a_45782_17890# a_12899_11471# a_45386_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16707 a_26495_41781# a_12473_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16708 a_43378_55166# VSS a_43870_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16709 a_23195_29967# a_22922_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1671 a_40366_59182# a_16362_59182# a_40458_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16710 a_26310_65206# a_12355_65103# a_26802_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16711 a_2196_47741# a_2079_47546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X16712 a_42099_43177# a_41167_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16713 a_11396_55535# a_8199_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X16714 VSS a_12877_14441# a_33734_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16715 vcm_commonmode a_16362_61190# a_42466_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16716 a_29322_58178# a_16362_58178# a_29414_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16717 VSS VSS a_16666_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16718 VDD a_10286_26311# a_10771_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16719 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1672 a_49894_19500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16720 vcm_commonmode a_16362_71230# a_25398_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16721 VSS a_12727_15529# a_46786_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16722 a_38295_29967# a_38210_30199# a_38077_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16723 a_43774_10862# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16724 a_10426_51549# a_9668_51451# a_9863_51420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16725 VDD a_12947_71576# a_37354_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16726 a_20778_55488# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16727 a_29322_17890# a_12899_10927# a_29814_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16728 a_46390_8854# a_16362_8488# a_46482_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16729 VSS a_12947_23413# a_29718_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1673 a_12985_19087# a_12815_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X16730 a_26706_20902# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16731 VSS a_2411_26133# a_2369_39037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16732 a_10673_15055# a_9865_14441# a_10589_15055# VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16733 a_38499_37503# a_37733_37477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16734 a_15285_52245# a_7050_53333# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16735 a_41370_7850# VDD a_41862_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16736 a_30326_12870# a_12877_16911# a_30818_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16737 a_38101_38565# a_38315_39141# a_39247_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X16738 a_9253_30511# a_8117_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16739 VSS a_24755_42325# a_16152_43677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1674 a_18770_64524# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16740 VSS a_9276_12167# a_9227_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16741 a_17274_7850# VDD a_17766_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16742 a_25006_47375# a_23929_47381# a_24844_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16743 VSS a_12727_13353# a_19678_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16744 VSS a_9275_15253# a_10117_14013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16745 a_36890_34191# a_36713_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16746 a_17843_48981# a_17668_49007# a_18022_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X16747 vcm_commonmode a_16362_70226# a_29414_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16748 a_23694_13874# a_12877_16911# a_23298_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16749 VSS a_12985_16367# a_20682_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1675 a_7030_31055# a_5449_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.55e+11p pd=5.31e+06u as=0p ps=0u w=1e+06u l=150000u
X16750 VSS a_11619_63151# a_11797_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16751 VSS a_2748_68565# result_out[10] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X16752 vcm_commonmode VSS a_30418_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16753 a_40387_31849# a_8491_41383# a_40315_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16754 a_27806_7452# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16755 a_23694_7850# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16756 a_29791_52436# a_25419_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16757 a_43378_72234# VSS a_43470_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16758 a_48794_63198# a_15439_49525# a_48398_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16759 VSS a_12727_58255# a_45782_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1676 a_10379_66389# a_10391_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16760 VSS a_11067_67279# a_45782_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16761 a_13919_27904# a_11602_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16762 a_24302_68218# a_12727_67753# a_24794_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16763 a_5411_12791# a_5775_12649# a_5710_12675# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16764 a_46482_8488# a_16746_8486# a_46390_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16765 a_35742_66210# a_12983_63151# a_35346_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16766 vcm_commonmode a_16362_62194# a_19374_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16767 VDD a_27359_43985# a_27219_44011# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16768 a_11667_63303# a_11943_63125# a_11901_63151# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16769 a_23390_60186# a_16746_60188# a_23298_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1677 a_23298_69222# a_16362_69222# a_23390_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16770 VDD a_10515_23975# a_33338_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16771 VDD a_12727_58255# a_27314_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16772 vcm_commonmode a_16362_16520# a_20378_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16773 a_23390_19532# a_16746_19530# a_23298_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16774 VDD a_8772_63927# a_8773_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16775 a_19807_27247# a_11902_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X16776 VDD a_2606_41079# a_19121_48502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16777 VDD a_11067_21583# a_46390_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16778 vcm_commonmode a_16362_15516# a_33430_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16779 a_20378_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1678 VDD a_12981_62313# a_22294_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16780 VDD a_1923_73087# a_1643_72917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16781 a_3670_70589# a_3452_70537# a_3588_70589# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16782 VDD a_12727_15529# a_36350_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16783 a_5510_18543# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16784 a_3983_24233# a_2315_24540# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16785 a_34434_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16786 VDD a_11067_46823# a_36519_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16787 a_2672_44655# a_1757_44655# a_2325_44897# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16788 VDD VSS a_19282_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16789 VSS a_14646_29423# a_20964_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1679 VSS a_12257_56623# a_25702_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X16790 a_37354_63198# a_16362_63198# a_37446_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16791 a_31422_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16792 a_47486_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16793 a_2012_12925# a_1895_12730# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16794 a_3972_25615# a_3529_25731# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X16795 a_33338_19898# a_11067_67279# a_33830_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16796 a_33080_37149# a_32795_36415# a_33668_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X16797 a_8746_71443# a_9063_71553# a_9021_71677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16798 a_23169_30539# a_3339_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16799 VDD a_28841_29575# a_29829_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X168 a_7215_36201# a_7019_35951# a_5490_41365# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.96e+12p pd=1.792e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X1680 a_9971_23439# a_9263_24501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16800 vcm_commonmode a_16362_67214# a_49494_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16801 a_37846_10464# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16802 a_15959_35327# a_14735_35805# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X16803 a_30722_71230# a_12947_71576# a_30326_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16804 a_34257_48169# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16805 a_11883_58575# a_11521_66567# a_11794_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16806 a_31184_36165# a_30311_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16807 a_2781_69513# a_1591_69141# a_2672_69513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X16808 VSS a_12727_67753# a_35742_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16809 a_6422_48285# a_5345_47919# a_6260_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1681 a_48890_9460# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16810 a_10614_54269# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16811 a_27406_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16812 vcm_commonmode a_16362_59182# a_39454_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16813 vcm_commonmode VSS a_25398_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16814 a_32795_38053# a_31096_38341# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X16815 a_43470_57174# a_16746_57176# a_43378_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16816 a_44778_18894# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16817 VSS a_3143_66972# a_7657_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X16818 a_26402_67214# a_16746_67216# a_26310_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16819 a_11883_58575# a_4351_67279# a_11711_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X1682 VSS a_75445_39738# a_75258_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16820 vcm_commonmode a_16362_64202# a_23390_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16821 a_29062_52093# a_2872_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16822 VSS a_12680_53511# a_11303_53511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X16823 a_25306_22910# a_16362_22544# a_25398_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16824 a_2952_66139# a_4075_69143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16825 VDD a_12355_65103# a_35346_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16826 a_37554_27247# a_30052_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16827 a_7803_11703# a_1929_10651# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16828 a_40458_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16829 a_14983_51157# a_17475_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X1683 VSS a_34759_31029# a_36193_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16830 VSS a_2163_57853# a_2124_57979# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16831 a_17670_61190# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16832 a_45386_9858# a_12546_22351# a_45878_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16833 VDD a_15439_49525# a_48398_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16834 VDD a_8082_56775# a_7169_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X16835 VSS a_12895_13967# a_21686_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16836 a_10873_27497# a_8935_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16837 a_3325_29967# a_2847_30271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X16838 a_26359_38007# a_26753_37981# a_13909_38659# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X16839 a_34725_38567# a_35033_38780# a_34699_38771# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1684 a_31611_43447# a_31648_43781# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X16840 a_7929_40125# a_4685_37583# a_7847_39872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16841 a_8453_64757# a_6515_62037# a_8957_65103# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X16842 VSS a_38454_34191# a_39331_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X16843 a_6791_70455# a_2952_66139# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X16844 VDD a_4941_35727# a_5693_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16845 a_36842_60508# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16846 VDD a_28881_52271# a_34895_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16847 VDD a_14919_37683# a_14945_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16848 VSS a_2375_48084# a_2079_47546# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X16849 a_49402_71230# a_12901_66665# a_49894_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1685 VDD a_23192_27791# a_27659_27275# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16850 a_44474_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16851 vcm_commonmode VSS a_17366_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16852 a_12120_54019# a_6095_44807# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X16853 a_22690_14878# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16854 a_4999_33781# a_2011_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16855 a_8395_37289# a_6372_38279# a_8177_37013# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16856 a_5457_13103# a_5399_13255# a_5023_13255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16857 VSS a_8273_42479# a_10607_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16858 a_13445_51335# a_12993_50345# a_13608_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X16859 VDD a_4433_55581# a_4533_55799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1686 a_16648_40517# a_16744_40517# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X16860 a_41370_24918# VSS a_41862_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16861 a_19678_58178# a_12901_58799# a_19282_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16862 a_7067_30663# a_2787_32679# a_7301_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16863 a_11307_57711# a_10957_57711# a_11212_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X16864 a_17449_46831# a_17171_46859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X16865 a_26802_71552# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16866 a_34738_67214# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16867 a_47486_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16868 VDD a_12985_19087# a_32334_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16869 a_12355_15055# a_15660_49257# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1687 VSS a_28841_29575# a_28799_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X16870 result_out[9] a_1644_66933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X16871 a_47790_66210# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16872 a_30735_49257# a_30005_48463# a_30663_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16873 a_45386_23914# a_12947_23413# a_45878_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16874 a_45386_19898# a_16362_19532# a_45478_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16875 VSS a_9179_13737# a_8815_13879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X16876 a_10689_29745# a_8273_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16877 a_34434_72234# VDD a_34342_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16878 vcm_commonmode a_16362_20536# a_49494_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16879 a_4427_25071# a_3983_25321# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1688 a_41370_65206# a_12355_65103# a_41862_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16880 VSS a_3325_49551# a_4073_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16881 VSS a_12947_56817# a_41766_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16882 a_35346_15882# a_12727_13353# a_35838_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16883 a_38850_18496# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16884 a_38754_24918# VSS a_38358_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16885 VSS a_11067_21583# a_35742_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16886 a_47486_71230# a_16746_71232# a_47394_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16887 VDD a_12727_13353# a_42374_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16888 a_27710_69222# a_12516_7093# a_27314_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16889 VSS a_10975_66407# a_24698_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1689 a_27406_11500# a_16746_11498# a_27314_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16890 a_28089_31157# a_25313_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16891 vcm_commonmode a_16362_12504# a_39454_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16892 VDD a_12215_31573# a_12161_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16893 a_3668_56311# a_4307_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X16894 a_9382_58255# a_6515_62037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X16895 a_48398_14878# a_12877_14441# a_48890_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16896 a_22786_23516# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16897 VDD a_28248_52271# a_28423_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16898 a_22386_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16899 a_49402_18894# a_16362_18528# a_49494_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X169 VSS a_5490_41365# a_5098_41391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1690 a_10901_54201# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16900 a_43470_10496# a_16746_10494# a_43378_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16901 a_23767_48463# a_23579_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X16902 a_26402_20536# a_16746_20534# a_26310_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16903 a_10421_14735# a_9865_14441# a_10339_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16904 VSS a_10615_72399# a_10949_72719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X16905 a_25398_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16906 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X16907 VSS a_21479_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X16908 a_8364_62723# a_7803_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16909 VSS a_12355_65103# a_28714_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1691 VDD a_12895_13967# a_26310_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16910 a_40458_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16911 VDD a_2437_28309# a_2467_28662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16912 a_33830_69544# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16913 VDD a_12899_11471# a_28318_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16914 a_27247_43047# a_12725_44527# a_27421_42923# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X16915 a_25798_14480# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16916 VSS a_2473_34293# a_5087_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16917 VSS a_6775_53877# a_4240_53083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16918 VSS a_25300_38567# a_25263_38825# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X16919 a_23298_15882# a_16362_15516# a_23390_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1692 a_44382_58178# a_16362_58178# a_44474_58178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16920 a_26402_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16921 a_29667_31055# a_29416_31171# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X16922 a_46882_68540# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16923 VDD a_10984_58487# a_6417_62215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16924 VDD a_22132_44129# a_21233_44220# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X16925 vcm_commonmode a_16362_18528# a_38450_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16926 VSS a_12257_56623# a_18674_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16927 a_11851_64391# a_11521_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16928 VSS a_3541_9593# a_3475_9661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16929 a_42466_16520# a_16746_16518# a_42374_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1693 a_30722_63198# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X16930 a_38115_52263# a_38524_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X16931 a_22690_55166# VSS a_22294_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16932 a_2012_51183# a_1867_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16933 a_30801_41835# a_12357_37999# a_30715_41835# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X16934 a_34342_65206# a_12355_65103# a_34834_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16935 VSS a_6795_51157# a_10045_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16936 a_29814_13476# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16937 a_26310_10862# a_12985_16367# a_26802_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16938 a_41766_58178# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16939 VDD a_12901_66959# a_23298_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1694 a_19282_60186# a_12727_58255# a_19774_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16940 VDD a_3572_56311# a_2419_55687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16941 a_1761_8751# a_1591_8751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X16942 a_47394_64202# a_11067_13095# a_47886_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16943 a_9869_49525# a_9651_49929# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16944 VDD a_12901_58799# a_19282_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16945 a_30323_44265# a_29391_44031# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16946 VSS a_5331_18517# a_5265_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16947 VDD a_11955_69653# a_11942_70045# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X16948 VDD a_2744_66103# a_1915_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16949 a_19678_11866# a_12985_16367# a_19282_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1695 vcm_commonmode a_16362_71230# a_40458_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X16950 a_12892_41807# a_12641_42036# a_12671_42134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X16951 a_34738_20902# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16952 vcm_commonmode a_16362_57174# a_32426_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16953 a_10265_10927# a_9642_10357# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16954 a_37354_56170# a_12947_56817# a_37846_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16955 a_11399_71855# a_11049_71855# a_11304_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X16956 VDD a_12727_67753# a_27314_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16957 a_1920_59861# a_2099_59861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X16958 a_11760_46983# a_7571_26151# a_11902_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16959 a_24794_64524# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1696 a_27314_68218# a_16362_68218# a_27406_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16960 a_21290_61190# a_12981_59343# a_21782_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16961 VDD VDD a_37354_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X16962 VSS VDD a_33734_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16963 a_8117_12559# a_1929_12131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16964 VDD a_2283_15797# a_1908_17141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X16965 a_43774_7850# VDD a_43378_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16966 a_30035_40767# a_29269_40741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X16967 a_4065_16617# a_3301_16617# a_3983_16617# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X16968 a_19680_31849# a_19626_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X16969 VDD a_4578_40455# a_4693_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1697 a_7635_64015# a_7213_62215# a_7445_63695# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X16970 a_27710_22910# a_11067_21583# a_27314_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16971 VSS a_12516_7093# a_36746_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16972 a_7657_66415# a_7387_66781# a_7567_66781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X16973 VSS a_5963_36585# a_5594_36727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16974 a_25306_60186# a_12727_58255# a_25798_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16975 a_34434_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16976 a_2380_68413# a_2263_68218# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X16977 a_10673_15055# a_10339_14735# a_10589_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=0p ps=0u w=1e+06u l=150000u
X16978 VDD a_32397_28023# a_31263_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X16979 a_33338_68218# a_16362_68218# a_33430_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1698 a_26157_31605# a_25263_29981# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X16980 a_8570_34319# a_6372_38279# a_7939_30503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X16981 a_45478_64202# a_16746_64204# a_45386_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16982 VSS a_49876_37608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.84e+07u l=3.9e+06u
X16983 a_2107_15113# a_1757_14741# a_2012_15101# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X16984 VDD a_41636_37601# a_42224_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X16985 VDD a_2319_57948# a_2250_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X16986 VSS a_12546_22351# a_24698_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16987 a_30479_48576# a_17682_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16988 a_47486_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16989 VSS a_41636_37601# a_40737_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X1699 a_39454_64202# a_16746_64204# a_39362_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16990 a_18770_55488# a_18602_55312# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16991 VDD a_12349_25847# a_12394_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16992 a_26505_31599# a_26157_31605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X16993 VSS a_12981_59343# a_39758_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16994 a_35438_56170# a_16746_56172# a_35346_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16995 a_36746_17890# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16996 a_22197_31171# a_20881_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X16997 a_41462_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X16998 a_43774_18894# a_12899_10927# a_43378_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16999 VSS a_12727_13353# a_40762_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_3173_66169# a_2840_66103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X170 a_31330_56170# a_16362_56170# a_31422_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1700 VDD a_27267_39605# a_1799_29556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X17000 a_35346_7850# VSS a_35438_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17001 a_8113_24527# a_5449_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17002 a_10846_60797# a_1950_59887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17003 VSS a_12985_16367# a_18674_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17004 a_45478_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17005 VSS a_17039_51157# a_22793_51005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17006 vcm_commonmode a_16362_62194# a_40458_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17007 a_41370_58178# a_10515_22671# a_41862_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17008 a_39454_55166# VDD a_39362_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17009 a_17493_50639# a_16902_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1701 a_10325_66415# a_9513_65301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17010 vcm_commonmode VSS a_23390_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17011 VSS a_12877_14441# a_44778_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17012 a_41766_11866# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17013 VSS a_20359_29199# a_30021_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17014 a_38358_10862# a_16362_10496# a_38450_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17015 a_10575_69439# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17016 a_30722_56170# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17017 a_5547_21379# a_4792_20443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17018 a_27600_36165# a_26631_35877# a_27504_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X17019 VDD VDD a_35346_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1702 a_44382_17890# a_12899_10927# a_44874_17492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17020 a_27314_18894# a_12895_13967# a_27806_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17021 VSS VSS a_27710_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17022 a_9260_25045# a_9167_24011# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17023 VDD a_41820_41501# a_40921_41245# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X17024 a_21290_8854# a_12985_19087# a_21782_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17025 a_31822_16488# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17026 a_6243_30662# a_5906_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X17027 VDD a_12947_71576# a_48398_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17028 vcm_commonmode a_16362_9492# a_40458_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17029 vcm_commonmode a_16362_10496# a_32426_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1703 VSS a_12947_23413# a_44778_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17030 a_18370_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17031 a_7293_45173# a_7075_45577# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X17032 a_2163_54589# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17033 VSS a_12899_11471# a_17670_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17034 a_48490_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17035 VSS a_2127_4943# a_2603_4943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17036 a_77002_39738# a_77098_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17037 a_21686_14878# a_12727_15529# a_21290_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17038 a_29220_50639# a_29055_49525# a_29118_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17039 a_30418_61190# a_16746_61192# a_30326_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1704 a_7363_62063# a_2840_53511# a_7267_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X17040 a_8443_47741# a_8295_47388# a_8080_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17041 a_14711_27247# a_12349_25847# a_14577_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X17042 a_2107_49929# a_1757_49557# a_2012_49917# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X17043 a_22294_69222# a_12901_66959# a_22786_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17044 a_33734_67214# a_12727_67753# a_33338_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17045 a_26402_9492# a_16746_9490# a_26310_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17046 vcm_commonmode a_16362_63198# a_17366_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17047 a_18278_59182# a_12901_58799# a_18770_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17048 a_13251_28111# a_11602_25071# a_13155_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17049 a_7000_43541# a_7847_40847# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1705 a_41766_20902# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17050 a_33313_51157# a_33697_50359# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17051 VDD a_8003_72917# a_9707_73807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17052 a_46786_66210# a_12983_63151# a_46390_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17053 vcm_commonmode a_16362_16520# a_31422_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17054 VDD a_10515_23975# a_44382_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17055 a_7377_32259# a_7281_29423# a_7295_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17056 a_33785_49007# a_33515_49007# a_33681_49373# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17057 a_10501_65871# a_10147_65984# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17058 a_12687_34191# a_12510_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17059 VSS a_16265_39868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X1706 VSS a_2284_36103# a_1591_36103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17060 a_23390_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17061 a_1761_37039# a_1591_37039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17062 a_28108_48783# a_27509_47695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17063 a_5713_74895# a_5441_72399# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17064 a_19374_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17065 VDD a_2325_18785# a_2215_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17066 VSS a_2928_22583# a_2007_20149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17067 vcm_commonmode a_16362_69222# a_43470_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17068 VDD a_12877_14441# a_34342_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17069 VSS a_7373_40847# a_8191_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X1707 a_11889_69679# a_10699_69679# a_11780_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17070 a_37076_37253# a_36107_36965# a_37039_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17071 VSS a_21663_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17072 a_11803_67503# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17073 a_45478_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17074 VDD a_11495_16341# a_11482_16733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17075 a_26020_30199# a_14926_31849# a_26251_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17076 a_26919_41271# a_25987_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17077 VDD a_4215_51157# a_27627_51733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X17078 a_41141_32143# a_35815_31751# a_41059_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17079 a_34906_47491# a_34062_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1708 a_5259_39367# a_5831_39189# a_5604_39215# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X17080 a_48398_63198# a_16362_63198# a_48490_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17081 a_38450_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17082 a_35346_66210# a_16362_66210# a_35438_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17083 a_21686_71230# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17084 VSS a_4792_20443# a_12541_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17085 a_20378_69222# a_16746_69224# a_20286_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17086 vcm_commonmode a_16362_68218# a_47486_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17087 a_35838_11468# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17088 VDD a_3016_60949# a_5245_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17089 a_3578_25625# a_2223_28617# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1709 VDD a_11067_67279# a_12901_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17090 VSS a_18127_35797# a_17939_36129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17091 a_2856_47753# a_1941_47381# a_2509_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X17092 a_39362_9858# a_16362_9492# a_39454_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17093 a_12013_64239# a_11710_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17094 VSS a_2292_43291# a_2369_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17095 VSS a_4711_54965# a_4642_54991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X17096 a_25398_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17097 a_49494_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17098 a_42770_60186# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17099 a_31669_51433# a_28881_52271# a_31871_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_2461_33597# a_2417_33205# a_2295_33609# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1710 a_21382_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17100 a_41462_58178# a_16746_58180# a_41370_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17101 a_42770_19898# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17102 VSS a_9707_51325# a_9668_51451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17103 a_28524_47919# a_26397_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17104 a_25702_70226# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17105 VDD a_5682_69367# a_10239_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X17106 a_24394_68218# a_16746_68220# a_24302_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17107 vcm_commonmode a_16362_65206# a_21382_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17108 VDD a_12677_42333# a_12283_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17109 VDD a_10717_53113# a_10747_52854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1711 a_1761_32143# a_1591_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17110 a_23298_23914# a_16362_23548# a_23390_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17111 VDD a_10975_66407# a_33338_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17112 a_39362_24918# VSS a_39854_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17113 a_18626_47375# a_18500_47491# a_18222_47507# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17114 a_43870_22512# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17115 VDD a_1586_18695# a_10883_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X17116 a_33430_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17117 VDD a_12355_65103# a_46390_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17118 a_22690_63198# a_15439_49525# a_22294_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17119 a_4287_65540# a_4167_64783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1712 VSS a_12727_13353# a_34738_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17120 a_19626_31751# a_19459_29423# a_19697_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X17121 a_28714_61190# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17122 a_27406_59182# a_16746_59184# a_27314_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17123 a_30326_71230# a_16362_71230# a_30418_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17124 a_33830_14480# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17125 a_33734_20902# a_11067_67279# a_33338_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17126 VSS a_12895_13967# a_32730_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17127 VDD a_12257_56623# a_36350_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17128 a_16762_24520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17129 a_2244_22583# config_1_in[13] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1713 a_37750_18894# a_12899_10927# a_37354_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17130 a_47394_72234# VDD a_47886_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17131 VDD a_11067_21583# a_20286_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17132 VDD a_12983_63151# a_19282_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17133 a_29829_49257# a_17682_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17134 a_44382_14878# a_16362_14512# a_44474_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17135 a_31551_31751# a_27535_30503# a_31725_31627# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17136 a_47886_60508# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17137 a_14611_46859# a_5039_42167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17138 a_19374_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17139 a_9215_58487# a_8592_58255# a_9560_58575# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X1714 a_24844_47753# a_23763_47381# a_24497_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X17140 a_9581_71855# a_7707_70741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X17141 vcm_commonmode VSS a_28410_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17142 a_7369_24233# a_6989_24233# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17143 a_34342_10862# a_12985_16367# a_34834_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17144 a_12831_35645# a_12651_35645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17145 a_11909_63695# a_11803_64239# a_9735_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17146 a_33734_14878# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17147 vcm_commonmode a_16362_22544# a_43470_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17148 VSS a_3016_60949# a_2960_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17149 a_17274_20902# a_12985_7663# a_17766_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1715 vcm_commonmode a_16362_70226# a_44474_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17150 a_24794_72556# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17151 a_1757_66415# a_1591_66415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17152 a_17274_16886# a_16362_16520# a_17366_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17153 a_21382_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17154 a_6459_38377# a_6372_38279# a_6377_38133# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17155 a_47790_9858# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17156 VDD a_12981_59343# a_24302_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17157 a_9556_49917# a_8569_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X17158 a_24302_62194# a_16362_62194# a_24394_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17159 a_45782_67214# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1716 a_12885_42134# a_12713_41923# a_12671_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X17160 a_10145_60405# a_9927_60809# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17161 a_36442_17524# a_16746_17522# a_36350_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17162 a_4031_73095# a_3751_72373# a_4429_72943# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X17163 VSS a_3247_20495# a_7628_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17164 a_7755_23145# a_4571_26677# a_8009_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X17165 a_2401_41941# a_2235_41941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17166 a_20378_22544# a_16746_22542# a_20286_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17167 vcm_commonmode a_16362_21540# a_47486_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17168 a_35742_59182# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17169 VDD a_10055_58791# a_27314_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1717 a_3215_68351# a_3040_68425# a_3394_68413# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17170 a_45478_72234# VDD a_45386_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17171 a_18674_69222# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17172 VSS a_2843_71829# a_5241_72765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17173 VSS a_12983_63151# a_22690_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17174 a_37751_49667# a_28881_52271# a_37655_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17175 VSS a_11771_23671# a_10286_26311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X17176 a_49894_18496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17177 vcm_commonmode a_16362_13508# a_37446_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17178 a_49798_24918# VSS a_49402_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17179 a_46390_15882# a_12727_13353# a_46882_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1718 a_10287_56118# a_8123_56399# a_9828_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X17180 a_8126_46287# a_7407_46529# a_7563_46261# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X17181 a_41462_11500# a_16746_11498# a_41370_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17182 VDD a_12895_13967# a_40366_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17183 a_24394_21540# a_16746_21538# a_24302_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17184 a_39758_58178# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17185 VDD a_4351_26159# a_4528_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X17186 VDD a_2656_45895# a_3983_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X17187 a_39758_16886# a_12727_13353# a_39362_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17188 a_36708_39655# a_35739_39679# a_36671_39913# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17189 VDD a_15439_49525# a_22294_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1719 a_21782_17492# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17190 VSS a_17039_51157# a_19913_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17191 a_7557_49007# a_7387_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17192 VDD a_5877_54421# a_5336_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17193 a_2369_23805# a_2325_23413# a_2203_23817# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17194 VDD a_12899_10927# a_26310_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17195 a_2834_22173# a_1757_21807# a_2672_21807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17196 a_36116_44765# a_35463_44031# a_36395_44265# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17197 a_8516_29199# a_6162_28487# a_8396_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X17198 a_15775_44581# a_13984_43781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X17199 VSS a_12889_39889# a_12921_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 a_45782_21906# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1720 a_21686_23914# a_10515_23975# a_21290_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17200 a_44874_69544# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17201 result_out[8] a_1644_65845# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17202 a_41370_66210# a_10975_66407# a_41862_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17203 a_27406_12504# a_16746_12502# a_27314_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17204 a_39454_63198# a_16746_63200# a_39362_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17205 vcm_commonmode a_16362_60186# a_36442_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17206 vcm_commonmode a_16362_19532# a_36442_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17207 a_4312_51005# a_3983_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X17208 a_9218_25071# a_5449_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17209 VDD a_32795_29967# a_33515_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1721 a_9747_67503# a_9301_67503# a_9651_67503# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X17210 a_1757_36501# a_1591_36501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17211 a_44382_59182# a_16362_59182# a_44474_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17212 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17213 VSS a_8994_63927# a_8636_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17214 VSS a_8543_36469# a_8423_39367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17215 VDD a_7841_12167# a_7959_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17216 a_19282_61190# a_12981_59343# a_19774_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17217 VSS a_21387_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17218 VSS a_1591_16367# a_1768_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17219 a_27314_69222# a_16362_69222# a_27406_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1722 VDD a_24755_42325# a_16152_43677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17220 VSS a_12257_56623# a_29718_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17221 vcm_commonmode a_16362_9492# a_49494_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17222 a_18487_28487# a_7571_29199# a_18661_28363# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17223 a_31422_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17224 a_2497_61519# a_2141_61635# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17225 a_1644_72373# a_1823_72381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17226 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17227 VDD a_12516_7093# a_21290_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17228 a_45386_65206# a_12355_65103# a_45878_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17229 a_4711_54965# a_4555_55233# a_4856_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X1723 VDD a_2693_68021# a_2583_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X17230 VSS a_12585_39069# a_12277_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17231 a_21382_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17232 a_4119_70741# a_3668_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X17233 a_12479_9633# a_11067_67279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17234 a_12345_26409# a_9955_20969# a_12263_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17235 vcm_commonmode a_16362_58178# a_30418_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17236 vcm_commonmode a_16362_71230# a_44474_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17237 a_75728_40202# a_75824_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17238 a_11396_65327# a_8999_61493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X17239 a_35346_57174# a_12257_56623# a_35838_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1724 vcm_commonmode a_16362_62194# a_34434_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17240 VDD a_12947_8725# a_41370_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17241 a_28011_41855# a_27245_41829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X17242 VDD a_7749_37903# a_8679_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17243 a_45782_20902# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17244 VSS a_12947_23413# a_48794_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17245 a_36520_42693# a_35647_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17246 a_18278_67214# a_12983_63151# a_18770_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17247 a_8625_20175# a_8015_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X17248 a_48398_56170# a_12947_56817# a_48890_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17249 a_22786_65528# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1725 a_35346_58178# a_10515_22671# a_35838_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17250 a_6559_63401# a_4119_70741# a_6641_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17251 VDD a_12947_8725# a_17274_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17252 a_32334_22910# a_10515_23975# a_32826_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17253 a_16060_28585# a_13390_29575# a_15599_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17254 VSS config_2_in[10] a_1591_44111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17255 VDD a_35676_49525# a_35598_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17256 a_2965_13967# a_2873_13879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17257 a_22294_55166# VSS a_22386_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17258 VSS a_12727_13353# a_38754_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17259 a_35742_12870# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1726 a_32334_21906# a_11067_21583# a_32826_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17260 a_16746_20534# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X17261 a_5541_53609# a_1952_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17262 a_21382_71230# a_16746_71232# a_21290_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17263 a_42770_13874# a_12877_16911# a_42374_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17264 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17265 a_23694_8854# a_12947_8725# a_23298_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17266 a_18674_22910# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17267 a_10531_31055# a_10280_31171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X17268 a_25702_23914# a_10515_23975# a_25306_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17269 a_22294_14878# a_12877_14441# a_22786_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1727 a_32334_17890# a_16362_17524# a_32426_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17270 VSS a_12985_7663# a_22690_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17271 a_21140_28335# a_20027_27221# a_5915_35943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17272 a_25798_56492# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17273 VSS a_27869_50095# a_29561_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X17274 a_6913_64239# a_6375_64489# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17275 a_4495_35925# a_5405_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X17276 a_16008_28111# a_13390_29575# a_15851_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.9325e+11p ps=2.51e+06u w=650000u l=150000u
X17277 a_2325_51425# a_2107_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X17278 a_16746_18526# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X17279 VSS a_41842_27221# a_20267_30503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1728 VDD a_3983_68591# a_1923_73087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X17280 VSS a_12516_7093# a_47790_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17281 VSS a_6417_62215# a_6365_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17282 a_39362_58178# a_10515_22671# a_39854_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17283 VSS a_2411_18517# a_10713_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17284 VSS a_29513_34428# a_29205_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17285 a_8733_29967# a_3339_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X17286 a_12879_38517# a_13067_38517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17287 a_12671_42134# a_12641_42036# a_12599_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17288 a_39758_11866# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17289 a_45478_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1729 VDD a_12727_58255# a_42374_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17290 a_9828_56311# a_7479_54439# a_9970_56118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17291 a_3478_41935# a_2401_41941# a_3316_42313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17292 a_1803_19087# a_1626_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17293 a_10394_19605# a_5671_21495# a_11564_19631# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X17294 VDD a_22989_48437# a_23019_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X17295 a_29943_41317# a_28980_41831# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X17296 VSS a_12355_15055# a_37750_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17297 a_41766_60186# a_12981_59343# a_41370_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17298 a_41766_19898# a_12895_13967# a_41370_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17299 a_10513_48161# a_10295_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X173 a_6559_59663# a_26662_48981# a_26610_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X1730 vcm_commonmode VSS a_17366_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17300 a_29814_55488# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17301 a_24698_70226# a_12901_66665# a_24302_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17302 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17303 VSS a_6372_38279# a_8480_38127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17304 a_9493_54447# a_7803_55509# a_7265_56053# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17305 a_25398_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17306 a_28410_61190# a_16746_61192# a_28318_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17307 VDD VSS a_38358_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17308 a_8662_28111# a_3607_34639# a_8576_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17309 vcm_commonmode a_16362_17524# a_25398_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1731 a_11902_47158# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X17310 a_20778_7452# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17311 a_4985_61021# a_1823_62589# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17312 VSS a_27155_40871# a_15459_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X17313 VSS a_12985_16367# a_29718_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17314 a_2847_45503# a_2672_45577# a_3026_45565# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17315 a_9198_53903# a_6515_62037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17316 VSS a_7623_13621# a_6738_19783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17317 a_12300_22895# a_11574_22869# a_11130_22869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X17318 a_5871_47594# a_5963_47349# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17319 a_2865_58799# a_2695_58799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1732 VSS a_12877_14441# a_38754_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17320 VDD a_3112_19319# a_3063_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17321 a_14951_39997# a_14963_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17322 a_33430_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17323 vcm_commonmode a_16362_16520# a_29414_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17324 a_39854_20504# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17325 VDD VDD a_46390_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17326 a_39454_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17327 a_9765_32143# a_9318_32509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17328 vcm_commonmode a_16362_11500# a_30418_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17329 a_40458_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1733 a_35742_11866# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17330 VSS a_24800_43041# a_23901_43132# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X17331 a_7009_33231# a_3607_34639# a_6883_37019# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17332 a_2375_48084# a_2467_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17333 a_46482_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17334 a_29414_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17335 a_26319_42869# a_12549_44212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17336 a_10754_62973# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17337 a_3026_71677# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17338 vcm_commonmode a_16362_64202# a_42466_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17339 VDD a_12546_22351# a_33338_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1734 a_21382_70226# a_16746_70228# a_21290_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17340 a_27937_27247# a_27659_27275# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17341 a_17691_27791# a_12631_28585# a_17774_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17342 VSS a_23901_35516# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17343 a_2111_38279# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17344 a_44382_22910# a_16362_22544# a_44474_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17345 VSS a_6786_37557# a_7749_37903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17346 a_19374_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17347 VSS a_52778_39936# a_53260_40156# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17348 a_33338_69222# a_12901_66959# a_33830_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17349 VDD a_19410_43439# a_26267_43983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1735 vcm_commonmode a_16362_61190# a_47486_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17350 a_12631_52928# a_12755_53030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17351 a_44778_67214# a_12727_67753# a_44382_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17352 vcm_commonmode a_16362_63198# a_28410_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17353 a_19678_71230# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17354 a_18370_69222# a_16746_69224# a_18278_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17355 a_9943_69135# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17356 a_26162_49007# a_26218_48981# a_6559_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X17357 VSS a_27183_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17358 a_17274_24918# VSS a_17366_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17359 a_2989_45717# a_2656_45895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X1736 a_7624_68021# a_7155_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X17360 VDD a_11145_60431# a_11449_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17361 a_22132_40865# a_21479_40229# a_22411_40183# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17362 a_21382_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17363 a_34738_59182# a_12727_58255# a_34342_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17364 VSS a_6895_15253# a_6829_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17365 a_17366_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17366 a_23205_51017# a_22015_50645# a_23096_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17367 a_27797_29423# a_27422_29789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17368 a_6637_20407# a_3247_20495# a_6800_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17369 a_22260_39655# a_21387_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1737 VDD a_2663_43541# a_2419_48783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X17370 a_33669_48829# a_32856_48463# a_33597_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17371 vcm_commonmode a_16362_65206# a_19374_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17372 a_24698_24918# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17373 a_9751_25071# a_9218_25321# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X17374 VSS a_27560_34337# a_26661_34428# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X17375 a_30722_17890# a_12899_11471# a_30326_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17376 a_38754_58178# a_12901_58799# a_38358_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17377 VSS VSS a_35742_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17378 VSS a_33694_30761# a_35581_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17379 VDD a_12981_59343# a_32334_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1738 a_24698_56170# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17380 a_3325_69135# a_2847_69439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17381 VDD a_7407_46529# a_7368_46403# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X17382 a_49494_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17383 a_46390_66210# a_16362_66210# a_46482_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17384 a_10969_71631# a_10949_72719# a_10981_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X17385 a_9832_60797# a_9424_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17386 VDD a_35517_34954# a_26550_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X17387 a_7289_62607# a_7619_62581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17388 a_27710_15882# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17389 a_5462_18038# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1739 a_18674_21906# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17390 a_17417_31171# a_17358_31069# a_17322_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17391 VSS a_8268_35381# a_7078_36103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X17392 VSS a_12727_15529# a_31726_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17393 a_3983_30761# a_3417_33231# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X17394 a_7295_32259# a_6883_37019# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17395 a_24794_9460# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17396 VDD a_26523_29199# a_44177_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17397 VDD a_12947_71576# a_22294_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17398 a_40458_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17399 a_19559_44535# a_18627_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X174 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u M=33
X1740 a_48794_10862# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17400 a_36453_31599# a_28446_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17401 VDD a_12355_15055# a_18278_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17402 VSS a_10975_66407# a_43774_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17403 a_7691_12265# a_3327_9308# a_7583_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17404 a_41862_23516# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17405 a_41462_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17406 a_9556_49917# a_8569_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17407 VDD a_10975_66407# a_44382_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17408 a_9963_29967# a_8739_28879# a_10045_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X17409 a_5441_72399# a_5087_72512# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1741 a_35383_28111# a_21187_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.8675e+11p pd=3.79e+06u as=0p ps=0u w=650000u l=150000u
X17410 a_2141_61635# a_1823_72381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17411 a_26706_62194# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17412 a_44474_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17413 VSS a_12727_58255# a_30722_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17414 VSS a_11067_67279# a_30722_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17415 a_2325_40545# a_2107_40303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17416 VSS a_1915_21482# a_1867_21263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17417 VSS a_2952_66139# a_6641_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X17418 a_20682_66210# a_12983_63151# a_20286_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17419 VDD a_10515_22671# a_34342_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1742 a_22294_13874# a_12727_15529# a_22786_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17420 a_3018_47375# a_1941_47381# a_2856_47753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17421 a_11763_21237# a_12166_21501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17422 VDD a_12659_54965# a_12631_52928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17423 VDD a_12899_11471# a_47394_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17424 a_44874_14480# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17425 a_44778_20902# a_11067_67279# a_44382_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17426 VDD a_26112_30663# a_26063_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X17427 a_1761_47919# a_1591_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17428 a_42374_15882# a_16362_15516# a_42466_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17429 a_18370_22544# a_16746_22542# a_18278_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1743 a_36395_36649# a_35463_36415# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X17430 a_27806_24520# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17431 VSS a_12985_19087# a_46786_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17432 a_17366_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17433 VDD a_11067_21583# a_31330_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17434 VSS a_4314_40821# a_6653_36611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17435 a_34738_12870# a_10055_58791# a_34342_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17436 a_16224_27791# a_12985_25615# a_15851_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17437 a_17670_64202# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17438 vcm_commonmode a_16362_23548# a_41462_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17439 VDD a_12727_15529# a_21290_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1744 VSS a_7987_40821# a_7000_43541# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.053e+12p ps=1.104e+07u w=650000u l=150000u M=4
X17440 VDD a_11067_13095# a_12712_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17441 a_48890_13476# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17442 a_45386_10862# a_12985_16367# a_45878_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17443 VDD a_1645_42453# a_1593_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17444 a_13975_34191# a_13798_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17445 a_5132_52637# a_4918_52637# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17446 VDD a_12901_66959# a_42374_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17447 a_22294_63198# a_16362_63198# a_22386_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17448 a_28318_20902# a_12985_7663# a_28810_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17449 a_43774_68218# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 a_25798_55488# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17450 a_28318_16886# a_16362_16520# a_28410_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17451 VSS a_15009_47919# a_15617_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17452 a_34434_18528# a_16746_18526# a_34342_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17453 VDD a_12901_58799# a_38358_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17454 VSS a_22448_38341# a_22521_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X17455 a_32426_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17456 VSS a_15959_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17457 a_38754_11866# a_12985_16367# a_38358_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17458 a_47486_17524# a_16746_17522# a_47394_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17459 a_27710_56170# a_12257_56623# a_27314_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1746 VDD a_53260_40156# a_53218_40254# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17460 a_12164_25321# a_9955_20969# a_12082_25077# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17461 a_18278_12870# a_12877_16911# a_18770_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17462 VDD a_12877_16911# a_25306_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17463 a_22786_10464# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17464 VDD a_3143_66972# a_5756_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X17465 a_39362_66210# a_10975_66407# a_39854_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17466 a_38171_43983# a_37994_43983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17467 a_48398_8854# a_16362_8488# a_48490_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17468 VSS a_12727_67753# a_20682_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17469 a_43870_64524# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1747 VDD a_51714_39886# a_52590_39936# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X17470 a_46786_59182# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17471 a_43378_7850# VDD a_43870_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17472 a_40366_61190# a_12981_59343# a_40858_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17473 vcm_commonmode a_16362_14512# a_35438_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17474 VDD a_8051_52047# a_8453_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17475 a_7097_63151# a_6559_63401# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17476 vcm_commonmode a_16362_59182# a_24394_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17477 vcm_commonmode VSS a_18370_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17478 a_24928_36391# a_24055_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X17479 a_19282_7850# VDD a_19774_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1748 a_30039_47919# a_26417_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17480 vcm_commonmode a_16362_13508# a_48490_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17481 a_33830_56492# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17482 VDD a_5199_11791# a_5601_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17483 a_35438_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17484 a_4987_58229# a_4792_58371# a_5297_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17485 VSS a_8635_61751# a_8039_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17486 a_5153_34025# a_2011_34837# a_5081_34025# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17487 a_29814_7452# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17488 a_25702_7850# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17489 VDD a_12355_65103# a_20286_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1749 a_33430_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17490 a_5547_31599# a_4495_35925# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X17491 a_36401_46859# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17492 a_44382_60186# a_12727_58255# a_44874_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17493 VSS a_2847_71615# a_2781_71689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X17494 a_6327_72917# a_6453_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17495 a_48490_8488# a_16746_8486# a_48398_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17496 a_25987_41317# a_25221_41281# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X17497 a_10497_10703# a_9642_10357# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17498 a_1757_29973# a_1591_29973# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17499 a_25398_13508# a_16746_13506# a_25306_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X175 a_7281_29423# a_6743_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1750 a_4792_41167# a_3949_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=0p ps=0u w=650000u l=150000u M=2
X17500 a_18012_32143# a_17798_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17501 a_32730_70226# a_12901_66665# a_32334_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17502 a_17274_62194# a_12355_15055# a_17766_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17503 a_1950_59887# a_1920_59861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17504 a_7815_45503# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17505 VSS a_4891_47388# a_27175_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17506 a_21782_60508# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17507 VSS a_10515_22671# a_27710_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17508 a_37446_66210# a_16746_66212# a_37354_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17509 a_30720_51183# a_30762_49641# a_30530_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1751 a_6614_21237# a_5535_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17510 a_5281_11791# a_4429_14191# a_5199_11791# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17511 VSS a_1586_21959# a_10883_18007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17512 a_36350_21906# a_16362_21540# a_36442_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17513 a_39454_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17514 a_5449_25071# a_5085_23047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X17515 a_6825_29423# a_5441_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17516 a_4555_55233# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17517 a_35742_61190# a_12355_15055# a_35346_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17518 a_31083_36395# a_26433_39631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17519 a_2873_52271# a_1683_52271# a_2764_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1752 a_24394_61190# a_16746_61192# a_24302_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17520 vcm_commonmode VSS a_42466_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17521 a_18674_71230# a_12947_71576# a_18278_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17522 a_32426_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17523 VSS VSS a_46786_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17524 a_43774_21906# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17525 a_32730_66210# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17526 a_46390_57174# a_12257_56623# a_46882_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17527 a_13097_36367# a_12671_36694# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17528 a_7199_62839# a_7077_62313# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X17529 VDD a_9414_10383# a_9490_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1753 VDD a_12899_3311# a_34342_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17530 a_30326_23914# a_12947_23413# a_30818_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17531 a_30326_19898# a_16362_19532# a_30418_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17532 a_4987_58229# a_4831_58497# a_5132_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X17533 VSS a_12899_11471# a_36746_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17534 VSS a_1643_72917# a_1591_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17535 a_33203_34191# a_33026_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17536 a_8205_75369# a_7901_74281# a_8059_74746# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17537 a_40762_14878# a_12727_15529# a_40366_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17538 a_34434_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17539 vcm_commonmode VSS a_27406_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1754 vcm_commonmode a_16362_17524# a_21382_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17540 a_5265_23145# a_5085_24759# a_5169_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17541 a_33338_55166# VSS a_33430_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17542 VDD a_35431_31751# a_25787_28327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X17543 a_28103_38591# a_27337_38565# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X17544 a_7295_56399# a_7265_56053# a_7201_56399# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X17545 VSS a_12727_13353# a_49798_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17546 a_46786_12870# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17547 a_23790_18496# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17548 a_23694_24918# VSS a_23298_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17549 VSS a_29483_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X1755 a_2875_61225# a_2497_61519# a_2657_60949# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17550 a_20286_15882# a_12727_13353# a_20778_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17551 VSS a_11067_21583# a_20682_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17552 a_17366_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17553 a_32426_71230# a_16746_71232# a_32334_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17554 VDD a_35932_41953# a_35033_42044# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X17555 VDD a_14681_50247# a_14511_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17556 vcm_commonmode a_16362_12504# a_24394_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17557 a_33338_14878# a_12877_14441# a_33830_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17558 a_7775_10625# a_1586_18695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17559 VSS a_3949_41935# a_4578_40455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1756 a_20964_31029# a_5915_35943# a_21184_31375# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X17560 a_10473_47713# a_10407_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17561 a_37354_59182# a_12901_58799# a_37846_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17562 a_31819_35073# a_30757_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17563 a_29943_34789# a_29177_34753# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X17564 vcm_commonmode a_16362_62194# a_49494_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17565 a_47394_9858# a_12546_22351# a_47886_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17566 VDD a_1586_36727# a_2971_37589# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X17567 a_26706_15882# a_12877_14441# a_26310_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17568 VDD a_1761_31055# a_32327_35839# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X17569 VSS a_12981_62313# a_35742_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1757 VDD a_13123_38231# a_13111_37999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17570 a_23501_42583# a_23597_42325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17571 a_27683_52271# a_27167_52271# a_27588_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17572 VDD a_14963_39783# a_18949_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X17573 a_19621_52521# a_4758_45369# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17574 a_33856_44869# a_32887_44581# a_33819_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17575 a_38450_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17576 a_6393_34837# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17577 a_16012_41959# a_15193_41781# a_16154_41807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17578 a_31822_68540# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17579 a_26402_62194# a_16746_62196# a_26310_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1758 VSS a_4685_37583# a_8268_35381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X17580 a_27806_58500# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17581 VDD a_2411_18517# a_11756_12381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17582 vcm_commonmode a_16362_18528# a_23390_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17583 a_12381_35836# a_32003_35307# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X17584 a_6749_66959# a_2952_66139# a_6156_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17585 VSS a_1683_27399# a_1683_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17586 VSS a_10055_58791# a_27710_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17587 a_31904_30511# a_30790_30663# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X17588 a_14912_27497# a_14287_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17589 a_7195_65564# a_7000_65595# a_7505_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X1759 a_28714_13874# a_12877_16911# a_28318_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17590 VSS a_39727_27765# a_39673_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17591 a_40458_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17592 VDD VSS a_49402_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17593 a_33797_28585# a_4811_34855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X17594 a_25961_48169# a_4891_47388# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17595 a_5504_37815# a_4314_40821# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17596 a_32397_28023# a_21187_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17597 a_40762_71230# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17598 a_4124_64391# a_1768_13103# a_4266_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17599 VSS a_11067_13095# a_39758_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X176 a_51330_39932# a_49876_41198# a_51422_39932# VDD sky130_fd_pr__pfet_01v8 ad=1.24e+12p pd=9.24e+06u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u M=2
X1760 VSS a_12985_16367# a_25702_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X17600 a_32334_64202# a_11067_13095# a_32826_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17601 VDD a_7707_70741# a_9333_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X17602 a_37846_21508# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17603 a_37446_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17604 a_22164_51157# a_22015_51840# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17605 VSS a_2411_26133# a_2369_30333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X17606 a_26779_50461# a_26155_50095# a_26671_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17607 a_44474_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17608 a_41370_60186# a_16362_60186# a_41462_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17609 a_8459_71285# a_8746_71443# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1761 a_2107_71689# a_1591_71317# a_2012_71677# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X17610 a_22294_56170# a_12947_56817# a_22786_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17611 VDD a_6514_37191# a_5701_37013# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17612 VSS a_29927_29199# a_38067_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17613 VSS a_29943_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17614 a_44778_70226# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17615 a_43470_68218# a_16746_68220# a_43378_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17616 VSS a_3339_30503# a_26350_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X17617 vcm_commonmode a_16362_65206# a_40458_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17618 a_1761_8751# a_1591_8751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X17619 VSS a_5085_23047# a_7939_27497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1762 a_10430_16950# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X17620 a_42374_23914# a_16362_23548# a_42466_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17621 VSS a_12677_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17622 a_6791_70455# a_7063_70313# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17623 a_38358_13874# a_16362_13508# a_38450_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17624 VDD a_12546_22351# a_44382_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17625 VSS a_5024_67885# a_6515_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17626 a_17366_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17627 VSS a_12263_4391# a_12815_4399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17628 VDD a_2509_47349# a_2399_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17629 VSS a_18307_27791# a_18848_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1763 VSS a_31223_36369# a_31169_36395# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17630 a_34738_62194# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17631 a_3417_10927# a_3247_10927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17632 VDD a_11709_55777# a_11599_55901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17633 a_23385_28585# a_23298_28487# a_23303_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17634 a_17670_72234# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17635 VSS a_1867_32839# a_1867_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17636 a_13867_35606# a_13097_36367# a_13795_35606# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X17637 VSS a_12516_7093# a_21686_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17638 a_47790_61190# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17639 VDD a_4528_26159# a_7343_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X1764 a_10173_51183# a_9794_51549# a_10101_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17640 a_46482_59182# a_16746_59184# a_46390_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17641 vcm_commonmode a_16362_56170# a_43470_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17642 a_2228_61879# a_2041_61519# a_2141_61635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X17643 VSS a_4220_57685# a_2944_57960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X17644 a_2672_69513# a_1757_69141# a_2325_69109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X17645 VDD a_6921_72943# a_7755_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X17646 a_29414_69222# a_16746_69224# a_29322_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17647 vcm_commonmode a_16362_66210# a_26402_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17648 a_30418_64202# a_16746_64204# a_30326_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17649 a_4887_36495# a_4443_36611# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1765 a_5449_32687# a_4259_32687# a_5340_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17650 a_28318_24918# VSS a_28410_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17651 a_42466_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17652 a_53714_40254# a_52778_39936# a_53260_40156# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17653 VDD a_12983_63151# a_38358_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17654 a_35838_63520# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17655 a_32426_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17656 a_4956_43567# a_4839_43780# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X17657 VDD a_3143_66972# a_7567_66781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X17658 a_7107_58487# a_5024_67885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17659 a_32397_28023# a_32167_29611# a_32560_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1766 a_48398_72234# VSS a_48490_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17660 a_38450_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17661 a_18370_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17662 VSS a_12981_59343# a_24698_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17663 a_20378_56170# a_16746_56172# a_20286_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17664 a_21686_17890# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17665 a_2012_18543# a_1895_18756# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17666 VSS a_28757_27247# a_31033_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17667 vcm_commonmode VSS a_47486_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17668 a_2475_68425# a_1959_68053# a_2380_68413# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X17669 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1767 a_2464_54813# a_2250_54813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17670 a_14761_36165# a_15069_35805# a_14735_35805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X17671 a_5320_18231# a_5535_18012# a_5462_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17672 VSS a_38239_32375# a_39305_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17673 a_43870_72556# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17674 a_39854_62516# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17675 VDD a_32143_35281# a_32003_35307# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17676 a_49798_58178# a_12901_58799# a_49402_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17677 VDD a_12981_59343# a_43378_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17678 a_43678_31029# a_43680_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17679 VSS a_12727_58255# a_28714_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1768 a_27411_50069# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17680 a_24394_55166# VDD a_24302_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17681 a_25702_16886# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17682 VSS a_11067_67279# a_28714_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17683 a_2899_16367# a_2283_15797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17684 a_6722_65579# a_7000_65595# a_6956_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17685 VDD a_6098_73095# a_6559_72512# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17686 a_9167_24011# a_6559_22671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17687 a_23298_10862# a_16362_10496# a_23390_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17688 a_18637_29451# a_13390_29575# a_18551_29451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X17689 VDD a_28789_50613# a_19478_51959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1769 a_29322_68218# a_12727_67753# a_29814_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17690 VDD VDD a_20286_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17691 VDD a_12792_51017# a_12967_50943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17692 a_37750_69222# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17693 VSS a_27183_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17694 a_5537_37039# a_5449_37191# a_5455_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17695 VSS a_12983_63151# a_41766_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17696 VSS a_1929_12131# a_5867_11995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17697 VDD a_12355_15055# a_29322_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17698 result_out[11] a_1644_70197# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X17699 VSS a_24959_30503# a_33135_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 a_48398_57174# a_12257_56623# a_48890_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1770 a_21356_31055# a_14646_29423# a_21101_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X17700 VSS a_2235_30503# a_25462_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X17701 vcm_commonmode a_16362_23548# a_39454_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17702 a_8296_54697# a_8199_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X17703 VSS a_2317_28892# a_3801_24643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X17704 a_43470_21540# a_16746_21538# a_43378_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17705 a_17274_70226# a_12516_7093# a_17766_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17706 a_38358_58178# a_16362_58178# a_38450_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17707 a_40762_9858# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17708 a_25313_31599# a_24746_31849# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X17709 a_45782_7850# VDD a_45386_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1771 a_30326_63198# a_12981_62313# a_30818_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17710 VDD a_7050_53333# a_15505_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X17711 a_4989_42255# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17712 a_3588_70589# a_3452_70537# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17713 VDD a_1923_59583# a_2464_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17714 a_38358_17890# a_12899_10927# a_38850_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17715 a_27314_11866# a_16362_11500# a_27406_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17716 a_33430_13508# a_16746_13506# a_33338_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17717 a_42866_15484# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17718 VDD a_12899_10927# a_45386_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17719 a_4789_52271# a_4311_52245# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1772 a_28410_60186# a_16746_60188# a_28318_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17720 a_31726_66210# a_12983_63151# a_31330_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17721 a_36643_27247# a_22291_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17722 a_5147_50943# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17723 a_7115_58575# a_6467_55527# a_6978_58487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X17724 a_46482_12504# a_16746_12502# a_46390_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17725 a_27981_37477# a_27183_36965# a_28115_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X17726 VSS a_12546_22351# a_26706_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17727 VDD a_6831_63303# a_32311_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17728 a_3392_73853# a_3275_73658# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X17729 a_29414_22544# a_16746_22542# a_29322_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1773 a_49798_7850# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X17730 a_36717_47375# a_36448_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17731 vcm_commonmode a_16362_70226# a_38450_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17732 VDD a_6752_29941# a_6825_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17733 VSS a_12727_67753# a_18674_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17734 a_9370_69831# a_9466_69653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17735 VSS a_12257_56623# a_48794_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17736 VSS a_1923_73087# a_3670_70589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17737 a_37354_7850# VSS a_37446_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17738 a_32038_29575# a_30788_28487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X17739 a_43378_11866# a_10055_58791# a_43870_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1774 a_28410_19532# a_16746_19530# a_28318_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17740 a_2107_26159# a_1757_26159# a_2012_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X17741 a_2672_69513# a_1591_69141# a_2325_69109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17742 a_28714_64202# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17743 a_26310_21906# a_11067_21583# a_26802_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17744 VDD a_12516_7093# a_40366_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17745 a_26310_17890# a_16362_17524# a_26402_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17746 VDD a_12727_58255# a_36350_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17747 a_47486_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17748 a_10378_67869# a_9301_67503# a_10216_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17749 a_30418_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1775 VDD a_10515_23975# a_38358_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X17750 a_8289_14741# a_8123_14741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17751 a_33338_63198# a_16362_63198# a_33430_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17752 a_18674_56170# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17753 a_5784_16367# a_5533_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17754 a_45478_18528# a_16746_18526# a_45386_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17755 VDD a_12901_58799# a_49402_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17756 a_5915_35943# a_20027_27221# a_20794_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X17757 a_23390_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17758 a_20286_66210# a_16362_66210# a_20378_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17759 a_25702_57174# a_10515_22671# a_25306_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1776 vcm_commonmode a_16362_16520# a_25398_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17760 a_19774_16488# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17761 a_10753_12559# a_10351_12879# a_10589_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X17762 vcm_commonmode a_16362_68218# a_32426_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17763 a_49798_11866# a_12985_16367# a_49402_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17764 a_20778_11468# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17765 VDD a_16265_39868# a_15871_39913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17766 a_37354_67214# a_12983_63151# a_37846_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17767 a_20575_47713# a_4443_46607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17768 VDD config_1_in[12] a_1626_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17769 a_41862_65528# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1777 a_35838_20504# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17770 a_23298_8854# a_12985_19087# a_23790_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17771 a_5121_35407# a_5079_35639# a_5025_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X17772 VSS a_15095_41781# a_15009_40193# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17773 VSS a_1915_20394# a_1867_20175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17774 vcm_commonmode a_16362_9492# a_42466_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17775 a_12935_31287# a_11719_28023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X17776 vcm_commonmode a_16362_14512# a_46482_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17777 a_37750_22910# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17778 VSS a_12381_43957# a_26495_42869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17779 VSS a_12985_7663# a_41766_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1778 a_35438_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17780 VSS a_26319_36341# a_19096_36513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17781 a_44874_56492# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17782 a_10862_10091# a_11140_10107# a_11096_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17783 a_24302_24918# VSS a_24794_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17784 VSS a_7000_43541# a_15575_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17785 a_28410_9492# a_16746_9490# a_28318_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17786 a_27806_66532# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17787 VDD a_12355_65103# a_31330_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17788 VDD a_77285_40202# a_77098_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17789 a_33748_51727# a_33360_51701# a_32582_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X1779 a_3972_25615# a_3529_25731# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17790 a_5172_54223# a_3016_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17791 a_27314_56170# a_16362_56170# a_27406_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17792 a_16735_51183# a_16385_51183# a_16640_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X17793 a_9651_67503# a_9135_67503# a_9556_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17794 VDD a_12257_56623# a_21290_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17795 VSS VDD a_39758_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17796 a_35438_67214# a_16746_67216# a_35346_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17797 a_32334_72234# VDD a_32826_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17798 VSS a_12818_52521# a_12680_53511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17799 a_43774_70226# a_12901_66665# a_43378_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X178 a_12901_52521# a_12202_54599# a_12818_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1780 a_26350_28585# a_2787_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X17800 VDD a_18053_28879# a_23447_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.646e+11p ps=2.94e+06u w=420000u l=150000u
X17801 VSS a_33839_28309# a_35616_27765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17802 a_28318_62194# a_12355_15055# a_28810_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17803 a_32826_60508# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17804 vcm_commonmode a_16362_17524# a_44474_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17805 VSS a_11067_21583# a_18674_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17806 a_33734_62194# a_12981_62313# a_33338_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17807 VSS a_12985_16367# a_48794_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17808 VDD VSS a_25306_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17809 a_16666_72234# VDD a_16270_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1781 a_38358_64202# a_16362_64202# a_38450_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17810 VDD a_2012_33927# a_2093_28918# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X17811 a_46786_61190# a_12355_15055# a_46390_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17812 a_29943_39141# a_29072_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X17813 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X17814 a_29718_71230# a_12947_71576# a_29322_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17815 a_30722_67214# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17816 a_21382_17524# a_16746_17522# a_21290_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17817 vcm_commonmode a_16362_8488# a_31422_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17818 a_16615_41001# a_15683_40767# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X17819 a_25702_10862# a_12546_22351# a_25306_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1782 a_7295_44647# a_17651_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X17820 a_7183_45199# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17821 vcm_commonmode a_16362_21540# a_32426_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17822 a_20442_28111# a_20027_27221# a_20359_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X17823 a_4399_48084# a_4491_47893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X17824 a_20682_59182# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17825 a_48490_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17826 a_2882_63517# a_2124_63419# a_2319_63388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17827 VSS a_12899_11471# a_47790_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17828 a_30418_72234# VDD a_30326_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17829 a_10961_19087# a_10791_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1783 VDD a_1923_54591# a_4035_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17830 a_18351_37503# a_17585_37477# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X17831 a_45478_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17832 a_35838_71552# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17833 a_4333_22351# a_3143_22364# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17834 a_3173_53333# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17835 a_4490_10383# a_3413_10389# a_4328_10761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X17836 VDD a_11067_67279# a_35346_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17837 vcm_commonmode a_16362_13508# a_22386_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17838 VSS a_35033_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X17839 a_9215_58487# a_8491_57487# a_9382_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1784 a_20881_28111# a_20359_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17840 a_31330_15882# a_12727_13353# a_31822_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17841 a_3452_70537# a_3372_70197# a_3856_70589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17842 VSS a_16917_31573# a_11719_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X17843 a_4149_45743# a_3983_45743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17844 a_38450_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17845 a_35346_61190# a_16362_61190# a_35438_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17846 VSS a_4215_51157# a_16219_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17847 vcm_commonmode a_16362_63198# a_47486_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17848 VSS a_5535_18012# a_8581_18319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17849 a_18278_71230# a_16362_71230# a_18370_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1785 a_27201_48169# a_22989_48437# a_27105_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X17850 a_48398_59182# a_12901_58799# a_48890_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17851 a_10151_21379# a_10045_21379# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17852 a_24698_58178# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17853 vcm_commonmode a_16362_66210# a_34434_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17854 a_24698_16886# a_12727_13353# a_24302_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X17855 a_8201_62839# a_7676_61493# a_8364_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17856 a_2781_71689# a_1591_71317# a_2672_71689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X17857 a_39854_70548# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17858 a_36442_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17859 a_7825_36815# a_5915_35943# a_7479_36495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1786 a_42466_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17860 a_24055_36415# a_22448_37253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X17861 a_36746_69222# a_12516_7093# a_36350_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17862 a_39362_60186# a_16362_60186# a_39454_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17863 VDD a_23487_49007# a_23579_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17864 VDD a_37888_43983# a_37994_43983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17865 a_17691_27791# a_13390_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17866 a_24394_63198# a_16746_63200# a_24302_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17867 vcm_commonmode a_16362_60186# a_21382_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17868 a_25798_59504# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17869 a_49494_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1787 a_38557_32143# a_38288_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17870 vcm_commonmode a_16362_19532# a_21382_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17871 a_25388_35077# a_24515_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17872 a_35438_20536# a_16746_20534# a_35346_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17873 result_out[15] a_1644_76181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17874 VSS a_12355_65103# a_37750_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17875 a_4407_51017# a_3891_50645# a_4312_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X17876 a_30326_65206# a_12355_65103# a_30818_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17877 a_49798_9858# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17878 a_7803_55509# a_8307_66415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17879 a_33939_43439# a_33762_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1788 a_10589_14735# a_9083_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17880 a_1644_53877# a_1823_53885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17881 a_35438_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17882 VDD a_17939_36129# a_17763_35797# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X17883 a_17321_49249# a_17103_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X17884 VDD a_6619_16341# a_5535_18012# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X17885 VDD a_23928_28585# a_28607_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17886 a_35447_27247# a_22015_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17887 a_30762_49641# a_30520_50345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X17888 a_10337_10927# a_9219_11471# a_10265_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17889 a_34759_31029# a_39035_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1789 a_25398_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17890 a_4607_46109# a_3983_45743# a_4499_45743# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X17891 a_28410_64202# a_16746_64204# a_28318_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17892 a_20286_57174# a_12257_56623# a_20778_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17893 VDD a_4495_35925# a_4275_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X17894 VDD a_15607_46805# a_41510_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17895 VSS config_1_in[1] a_1591_9295# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X17896 a_30722_20902# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17897 VDD a_12355_15055# a_37354_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17898 a_33338_56170# a_12947_56817# a_33830_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17899 a_42466_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X179 a_32334_23914# a_12947_23413# a_32826_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1790 a_2748_68565# a_2927_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17900 VDD a_2411_18517# a_10935_11989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17901 a_1586_21959# a_1643_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X17902 a_18370_56170# a_16746_56172# a_18278_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17903 a_19678_17890# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17904 VSS a_12727_13353# a_23694_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17905 a_20682_12870# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17906 VSS a_7571_29199# a_12263_26409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17907 VSS a_35319_34191# a_35425_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17908 VDD a_2143_15271# a_4065_16617# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17909 a_1681_5175# a_1591_7119# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1791 a_11179_9981# a_1586_18695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17910 a_19517_31751# a_4674_40277# a_19680_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17911 a_45782_62194# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17912 a_5025_35407# a_4578_40455# a_4941_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17913 a_3173_53333# a_2840_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X17914 vcm_commonmode a_16362_57174# a_41462_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17915 a_28714_72234# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17916 VSS a_5085_24759# a_6162_28487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X17917 VSS a_12516_7093# a_32730_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17918 a_24302_58178# a_10515_22671# a_24794_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17919 a_21479_40229# a_20713_40193# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X1792 vcm_commonmode a_16362_69222# a_37446_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17920 VDD a_12727_67753# a_36350_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17921 a_24698_11866# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17922 a_30418_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17923 a_46882_24520# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17924 VSS a_6224_73095# a_6377_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X17925 a_36442_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17926 VDD a_2775_46025# a_2875_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17927 VDD a_12983_63151# a_49402_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17928 VSS a_12355_15055# a_22690_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17929 a_19374_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1793 a_2847_21781# a_2672_21807# a_3026_21807# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X17930 a_49494_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17931 VDD a_32920_34191# a_33026_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X17932 a_18222_47507# a_18539_47617# a_18497_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17933 VDD a_7000_43541# a_13615_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17934 a_36746_22910# a_11067_21583# a_36350_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17935 a_34342_21906# a_11067_21583# a_34834_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17936 a_34342_17890# a_16362_17524# a_34434_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17937 a_22595_42089# a_21663_41855# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17938 VDD a_12727_15529# a_40366_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17939 a_10571_74031# a_10055_74031# a_10476_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1794 a_41462_67214# a_16746_67216# a_41370_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17940 a_15911_31784# a_16087_31751# a_16297_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X17941 VDD a_8117_30287# a_8297_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17942 VDD VSS a_23298_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17943 a_47394_20902# a_12985_7663# a_47886_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17944 VDD a_5254_67503# a_9490_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X17945 a_47394_16886# a_16362_16520# a_47486_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17946 vcm_commonmode a_16362_58178# a_18370_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17947 a_10614_52271# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17948 a_33830_8456# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17949 a_34423_30287# a_26523_29199# a_32038_29575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1795 VSS a_5541_53609# a_6666_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17950 a_20341_30287# a_14625_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17951 a_37354_12870# a_12877_16911# a_37846_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17952 VSS a_7644_46805# a_8126_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17953 a_1815_10422# a_1633_10422# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X17954 a_21781_49007# a_21737_49249# a_21615_49007# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X17955 a_41862_10464# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17956 VDD a_12947_8725# a_43378_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17957 a_24794_20504# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17958 VDD a_10515_23975# a_27314_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17959 a_11753_60975# a_11709_61217# a_11587_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1796 a_11711_58255# a_11521_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X17960 a_24394_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17961 VDD VDD a_31330_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17962 a_5041_64061# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17963 a_11521_58951# a_11943_63125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X17964 a_27314_64202# a_16362_64202# a_27406_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17965 VSS a_5691_36727# a_6713_37903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17966 a_48794_69222# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17967 a_14081_35606# a_13909_35395# a_13867_35606# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X17968 a_14088_38543# a_13837_38772# a_13867_38870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X17969 a_31422_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1797 a_24643_28335# a_23195_29967# a_4811_34855# VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X17970 a_5825_20495# a_5963_20149# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17971 a_31753_47919# a_31186_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17972 vcm_commonmode VSS a_37446_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17973 a_12158_32143# a_10515_32143# a_12412_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X17974 VDD a_12877_14441# a_17274_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17975 a_10597_32143# a_4903_31849# a_10515_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X17976 VSS a_35932_38689# a_35033_38780# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X17977 a_25702_8854# a_12947_8725# a_25306_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17978 a_9424_60949# a_9643_63125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X17979 a_28318_70226# a_12516_7093# a_28810_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1798 a_13888_43781# a_13984_43781# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X17980 a_2325_18785# a_2107_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X17981 VSS a_12901_58799# a_42770_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17982 a_28410_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17983 a_36350_18894# a_12895_13967# a_36842_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17984 a_25306_12870# a_16362_12504# a_25398_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17985 a_11747_28639# a_9179_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17986 a_10589_15055# a_9083_13879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17987 a_40858_16488# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X17988 VSS a_3301_26703# a_7113_27253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X17989 VSS a_12901_66959# a_25702_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1799 VSS a_3023_16341# a_2981_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X17990 VSS a_4685_37583# a_7755_38991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17991 a_44474_13508# a_16746_13506# a_44382_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X17992 vcm_commonmode a_16362_10496# a_41462_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17993 a_33857_49007# a_32672_49007# a_33785_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17994 a_18770_11468# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17995 a_41370_8854# a_16362_8488# a_41462_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X17996 a_27406_23548# a_16746_23546# a_27314_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17997 a_11495_18543# a_11049_18543# a_11399_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17998 a_3137_73493# a_2971_73493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X17999 a_11797_66415# a_11710_58487# a_11713_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_20905_32143# a_3339_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X180 VSS a_4674_40277# a_5831_39189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1800 a_35969_28111# a_35550_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18000 a_2107_19631# a_1757_19631# a_2012_19631# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18001 a_2744_46983# a_2952_46805# a_2886_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18002 VDD a_10575_62911# a_10562_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18003 VSS a_10515_22671# a_46786_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18004 a_43774_55166# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18005 VSS a_1929_10651# a_7493_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18006 a_21184_31375# a_5915_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18007 a_17274_8854# a_16362_8488# a_17366_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18008 a_8220_13647# a_8117_12559# a_7623_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X18009 VSS a_32611_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X1801 a_36336_44007# a_35463_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18010 VSS a_12727_67753# a_29718_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18011 a_1757_66415# a_1591_66415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18012 a_26706_65206# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18013 a_49402_61190# a_12981_59343# a_49894_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18014 a_17366_15516# a_16746_15514# a_17274_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18015 a_36612_39655# a_35739_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18016 a_16746_66212# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X18017 a_27406_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18018 a_22786_7452# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18019 VSS a_1799_29556# a_4719_33239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1802 a_14926_31849# a_14747_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X18020 a_33543_41271# a_32611_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18021 a_41462_8488# a_16746_8486# a_41370_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18022 a_1644_71829# a_1591_63151# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18023 a_23694_58178# a_12901_58799# a_23298_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18024 VSS VSS a_20682_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18025 a_37750_71230# a_12947_71576# a_37354_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18026 a_26495_36341# a_12473_36341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18027 VSS a_28980_41831# a_28943_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18028 a_26802_61512# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18029 a_31330_66210# a_16362_66210# a_31422_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1803 a_6473_40277# a_6579_42255# a_6817_42255# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X18030 vcm_commonmode a_16362_11500# a_18370_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18031 VDD a_5795_27497# a_5823_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18032 VDD a_2847_36799# a_2834_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18033 a_1643_72917# a_1846_73195# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18034 VDD a_1929_10651# a_8071_13255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18035 a_17766_19500# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18036 a_11617_72097# a_11399_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X18037 a_48398_67214# a_12983_63151# a_48890_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18038 a_28691_49783# a_27869_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X18039 a_4831_52413# a_1586_51335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1804 a_40366_22910# a_16362_22544# a_40458_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18040 a_3595_37583# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18041 VSS a_2122_20719# a_2228_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18042 a_35742_23914# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18043 a_13241_27497# a_11866_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X18044 a_42770_24918# VSS a_42374_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18045 a_36442_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18046 a_42866_57496# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18047 a_48794_22910# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18048 a_25798_67536# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18049 a_6060_15279# a_5943_15492# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1805 a_8901_15101# a_8857_14709# a_8735_15113# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18050 a_6619_73719# a_5441_72399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18051 a_32730_16886# a_12727_13353# a_32334_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18052 VDD a_3016_60949# a_6929_53725# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X18053 a_9547_49007# a_4298_58951# a_9184_49159# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18054 a_25306_57174# a_16362_57174# a_25398_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18055 a_6059_14165# a_2004_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X18056 VSS a_15959_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X18057 a_8652_17289# a_7571_16917# a_8305_16885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18058 VDD a_26397_51183# a_32134_49159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18059 a_45782_15882# a_12877_14441# a_45386_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1806 a_36487_46859# a_27535_30503# a_36401_46859# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18060 VSS a_12877_16911# a_42770_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18061 a_5825_12265# a_3327_9308# a_5730_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18062 VSS a_4952_68279# a_4211_67655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18063 VSS a_10515_23975# a_25702_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18064 a_11057_25077# a_9669_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18065 a_33830_59504# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18066 a_11491_55535# a_10975_55535# a_11396_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18067 vcm_commonmode VSS a_20378_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18068 a_43537_27497# a_23395_32463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18069 vcm_commonmode a_16362_18528# a_42466_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1807 a_39454_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18070 a_46882_58500# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18071 a_18674_17890# a_12899_11471# a_18278_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18072 a_75794_40594# a_75628_40594# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X18073 a_13047_29575# a_6459_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18074 a_1586_36727# a_4035_33205# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18075 a_9183_72007# a_7925_72399# a_9581_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18076 a_28410_72234# VDD a_28318_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18077 VSS a_10055_58791# a_46786_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18078 a_30418_7484# VDD a_30326_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18079 a_16270_55166# VSS a_16762_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1808 a_36350_12870# a_16362_12504# a_36442_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18080 a_29322_15882# a_12727_13353# a_29814_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18081 VSS a_11067_21583# a_29718_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18082 VSS a_3016_60949# a_6169_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X18083 a_44778_62194# a_12981_62313# a_44382_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18084 a_30326_10862# a_12985_16367# a_30818_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18085 a_12341_3311# a_12171_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18086 a_8128_54223# a_6559_59663# a_7637_53877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18087 a_40366_9858# a_12546_22351# a_40858_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18088 VSS a_13576_42589# a_12677_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X18089 a_18907_48502# a_4482_57863# a_18907_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1809 a_30991_29397# a_31117_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X18090 VSS a_4903_31849# a_9405_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18091 VDD a_12901_58799# a_23298_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18092 a_2847_44629# a_2672_44655# a_3026_44655# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18093 a_11304_71855# a_10969_71631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18094 VSS a_12727_15529# a_19678_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18095 VSS a_14919_37683# a_14425_37981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X18096 a_23694_11866# a_12985_16367# a_23298_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18097 a_32426_17524# a_16746_17522# a_32334_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18098 a_5441_27791# a_5175_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18099 a_2882_56989# a_2124_56891# a_2319_56860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X181 VSS a_1952_60431# a_4600_62069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X1810 VSS a_10010_68021# a_9951_68367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X18100 VSS a_6608_19319# a_5135_19061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18101 a_16969_38365# a_16699_37999# a_16879_37999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18102 a_17300_51183# a_16219_51183# a_16953_51425# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X18103 VSS a_35815_31751# a_37287_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18104 a_43378_70226# a_16362_70226# a_43470_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18105 a_8152_58575# a_7773_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18106 a_26802_9460# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18107 a_1644_70197# a_1591_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18108 a_24302_66210# a_10975_66407# a_24794_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18109 a_11612_26409# a_7571_26151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1811 a_21516_47919# a_19788_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X18110 VSS a_40921_41245# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X18111 a_35742_64202# a_12355_65103# a_35346_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18112 vcm_commonmode a_16362_60186# a_19374_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18113 vcm_commonmode a_16362_19532# a_19374_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18114 a_31726_59182# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18115 vcm_commonmode a_16362_14512# a_20378_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18116 VDD a_12985_7663# a_33338_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18117 VSS a_6243_30662# a_7390_32693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X18118 a_3301_26703# a_2899_27023# a_3137_27023# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X18119 a_2012_51183# a_1867_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1812 a_22690_72234# VDD a_22294_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18120 a_36442_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18121 a_14553_30761# a_8197_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18122 VDD a_11067_67279# a_46390_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18123 vcm_commonmode a_16362_13508# a_33430_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18124 a_16270_72234# VSS a_16362_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18125 a_4149_24527# a_3801_24643# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X18126 a_49494_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18127 a_8191_40303# a_5363_30503# a_8095_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18128 a_20378_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18129 a_46390_61190# a_16362_61190# a_46482_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1813 VSS a_7159_22583# a_7111_22351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18130 VDD a_29513_42333# a_29119_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18131 VDD a_11709_65569# a_11599_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18132 a_3667_60405# a_3870_60563# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18133 a_23593_44007# a_23901_44220# a_23567_44211# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X18134 a_49798_71230# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18135 a_48490_69222# a_16746_69224# a_48398_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18136 VDD a_10055_58791# a_36350_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18137 vcm_commonmode a_16362_66210# a_45478_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18138 a_32589_32143# a_28757_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18139 VDD a_2143_15271# a_10965_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1814 a_2672_66415# a_1591_66415# a_2325_66657# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X18140 a_34434_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18141 VDD a_11067_21583# a_19282_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18142 a_47394_24918# VSS a_47486_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18143 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18144 VSS a_2216_28309# a_3063_34319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18145 VDD a_29055_49525# a_28994_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X18146 a_47486_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18147 VDD a_4052_73865# a_4227_73791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18148 VSS a_22351_47893# a_22285_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18149 VSS a_6637_20407# a_4839_21495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1815 VSS config_1_in[6] a_1591_2767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18150 a_2785_60151# a_1591_59343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X18151 VSS a_12985_19087# a_48794_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18152 VSS a_12981_59343# a_43774_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18153 a_40762_17890# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18154 a_18045_41281# a_17983_41855# a_18915_42089# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18155 VSS a_12901_66665# a_26706_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18156 a_22386_66210# a_16746_66212# a_22294_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18157 VDD a_2689_65103# a_6641_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18158 a_22176_47919# a_21095_47919# a_21829_48161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18159 vcm_commonmode a_16362_65206# a_49494_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1816 VDD a_22132_40865# a_21233_40956# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X18160 a_23303_31171# a_22399_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18161 a_21290_21906# a_16362_21540# a_21382_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18162 a_24394_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18163 a_7841_29423# a_5087_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18164 VDD a_2325_69109# a_2215_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18165 VSS a_1923_73087# a_1881_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18166 a_27271_37455# a_1761_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18167 a_38315_39141# a_36708_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X18168 VSS a_5975_71829# a_5909_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18169 a_27897_32219# a_26505_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X1817 a_8814_16911# a_7737_16917# a_8652_17289# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18170 a_27406_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18171 VSS a_9187_51157# a_6795_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18172 vcm_commonmode a_16362_57174# a_39454_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18173 a_20682_61190# a_12355_15055# a_20286_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18174 a_43470_55166# VDD a_43378_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18175 a_44778_16886# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18176 a_2860_43389# a_2742_42997# a_2788_43389# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X18177 VSS a_37761_44759# a_37706_44135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18178 a_1644_56053# a_1591_54447# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18179 a_42374_10862# a_16362_10496# a_42466_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1818 a_11127_53544# a_6095_44807# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18180 VSS a_32695_43455# a_32641_43777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18181 a_26402_65206# a_16746_65208# a_26310_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18182 a_7311_60975# a_7060_61225# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X18183 VSS a_7189_35015# a_5963_36585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18184 VDD a_1586_69367# a_1591_71317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18185 VSS VSS a_31726_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18186 a_23096_51017# a_22181_50645# a_22749_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18187 a_25306_20902# a_16362_20536# a_25398_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18188 a_28410_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18189 a_36350_69222# a_16362_69222# a_36442_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1819 VSS a_12546_22351# a_41766_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18190 VDD a_12981_62313# a_35346_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18191 a_31330_57174# a_12257_56623# a_31822_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18192 a_40458_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18193 VDD a_9424_60949# a_9649_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18194 VDD a_4993_32929# a_4883_33053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18195 a_6008_69679# a_5682_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X18196 VDD a_9529_28335# a_16060_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18197 a_45386_7850# VDD a_45878_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18198 a_17670_18894# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18199 VDD a_12355_15055# a_48398_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X182 a_32334_19898# a_16362_19532# a_32426_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1820 a_10204_18543# a_5671_21495# a_9983_18870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X18200 VSS a_12899_11471# a_21686_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18201 a_41385_28129# a_30052_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18202 a_17415_29423# a_14926_31849# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X18203 VSS a_34297_35516# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X18204 a_18016_46983# a_3339_32463# a_18158_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X18205 a_18053_28879# a_15851_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18206 a_29414_56170# a_16746_56172# a_29322_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18207 a_39758_7850# VDD a_39362_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18208 VDD a_12895_13967# a_39362_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18209 a_31726_12870# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 a_14076_35077# a_13107_34789# a_14039_34743# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X18210 a_43774_63198# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18211 a_23731_28023# a_9529_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18212 VSS start_conversion_in a_1591_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18213 a_1586_45431# a_7295_43031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18214 a_34222_43439# a_34045_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18215 VSS a_12901_66959# a_33734_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18216 VDD a_6224_73095# a_7571_72512# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X18217 a_27710_7850# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18218 a_22294_59182# a_12901_58799# a_22786_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18219 a_7571_22057# a_4571_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1822 VDD a_2099_59861# a_2695_44119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18220 a_27974_32459# a_27387_32373# a_27890_32459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18221 a_41370_22910# a_10515_23975# a_41862_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18222 a_19780_38341# a_18811_38053# a_19743_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18223 a_34434_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18224 a_9135_22895# a_4798_23759# a_9223_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18225 VDD a_34759_31029# a_37503_31393# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18226 VSS a_12981_62313# a_20682_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18227 a_1908_17141# a_2004_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18228 a_48490_22544# a_16746_22542# a_48398_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18229 a_17366_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1823 a_19374_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18230 a_25461_51183# a_25417_51425# a_25295_51183# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X18231 a_7079_52815# a_6467_53359# a_6985_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X18232 a_34738_65206# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18233 a_47486_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18234 VDD VDD a_32334_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18235 a_34834_17492# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18236 a_34738_23914# a_10515_23975# a_34342_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18237 a_23390_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18238 a_43531_29199# a_12907_27023# a_43362_28879# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X18239 a_47790_64202# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1824 VDD a_12907_56399# a_16362_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X18240 a_45386_21906# a_11067_21583# a_45878_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18241 a_45386_17890# a_16362_17524# a_45478_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18242 VDD a_28446_31375# a_36519_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18243 VDD a_36890_34191# a_37711_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18244 a_34434_70226# a_16746_70228# a_34342_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18245 a_37750_56170# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18246 a_32507_32463# a_31964_30485# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18247 a_38850_16488# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18248 VDD a_13669_35253# a_14081_35606# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18249 a_35346_13874# a_12727_15529# a_35838_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1825 a_30418_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18250 a_11849_12015# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18251 VDD a_9123_57399# a_3714_58345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X18252 a_27710_67214# a_12727_67753# a_27314_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18253 VSS a_11067_13095# a_24698_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18254 VSS a_11764_65845# a_9624_65301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X18255 a_18278_23914# a_12947_23413# a_18770_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18256 a_18278_19898# a_16362_19532# a_18370_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18257 vcm_commonmode a_16362_10496# a_39454_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18258 a_48398_12870# a_12877_16911# a_48890_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18259 a_22786_21508# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1826 a_8998_74575# a_7921_74581# a_8836_74953# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18260 a_22386_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18261 vcm_commonmode a_16362_9492# a_36442_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18262 a_25306_65206# a_16362_65206# a_25398_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18263 a_37446_61190# a_16746_61192# a_37354_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18264 a_17670_59182# a_12727_58255# a_17274_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18265 a_8569_25071# a_8215_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18266 a_35463_36415# a_31847_36893# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X18267 vcm_commonmode VSS a_29414_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18268 a_11311_74005# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18269 a_33830_67536# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1827 a_12901_51017# a_11711_50645# a_12792_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18270 a_40458_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18271 a_30023_41959# a_1761_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18272 VDD a_12877_14441# a_28318_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18273 a_25798_12472# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18274 VSS a_2511_23983# a_2411_19605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18275 a_23298_13874# a_16362_13508# a_23390_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18276 a_43445_28879# a_42709_29199# a_43362_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18277 a_46882_66532# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18278 a_43378_63198# a_12981_62313# a_43870_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18279 a_16362_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1828 a_19678_70226# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18280 vcm_commonmode a_16362_16520# a_38450_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18281 a_8383_27247# a_7939_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18282 a_6607_39991# a_3949_41935# a_6841_40125# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18283 a_42466_14512# a_16746_14510# a_42374_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18284 a_32730_61190# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18285 VSS a_10515_23975# a_33734_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18286 a_23929_47381# a_23763_47381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18287 a_31422_59182# a_16746_59184# a_31330_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18288 a_49402_9858# a_12546_22351# a_49894_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18289 a_25398_24552# VDD a_25306_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1829 a_18370_68218# a_16746_68220# a_18278_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18290 a_29322_66210# a_16362_66210# a_29414_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18291 VDD a_7891_64213# a_7657_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18292 VDD a_8531_70543# a_35061_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18293 a_29814_11468# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18294 a_10865_72719# a_5877_70197# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18295 VDD a_12257_56623# a_40366_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18296 VSS a_3325_69135# a_4075_69143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18297 a_4583_64566# a_1768_13103# a_4124_64391# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18298 a_19774_68540# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18299 VDD a_12983_63151# a_23298_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X183 a_32029_38565# a_32611_39141# a_33484_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X1830 a_16832_42919# a_15959_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X18300 a_20778_63520# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18301 a_47394_62194# a_12355_15055# a_47886_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18302 VSS a_3607_34639# a_7189_35015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18303 a_3417_10927# a_3247_10927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18304 VDD a_2843_71829# a_2601_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X18305 VSS a_1586_36727# a_7295_43031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18306 a_23390_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18307 a_26319_38517# a_24413_39087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18308 vcm_commonmode VSS a_32426_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18309 a_9707_73807# a_9353_72399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1831 VDD a_6260_74031# a_6435_74005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18310 VDD a_7571_29199# a_11711_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18311 a_27411_50069# a_27236_50095# a_27590_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18312 a_21382_9492# a_16746_9490# a_21290_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18313 a_35742_72234# VDD a_35346_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18314 a_2927_39733# a_3663_39991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18315 VDD a_10975_66407# a_27314_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18316 a_24794_62516# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18317 a_7571_31599# a_7695_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18318 a_4433_55581# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18319 a_4949_55357# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1832 a_30908_40743# a_31004_40743# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X18320 VSS a_4803_63669# a_4734_63695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18321 a_48794_71230# a_12947_71576# a_48398_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18322 a_8827_17215# a_8652_17289# a_9006_17277# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18323 a_32509_47081# a_21187_29415# a_28756_55394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18324 VSS a_10665_58487# a_10478_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18325 a_30311_40229# a_29545_40193# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X18326 VSS a_28295_31287# a_28244_31415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X18327 a_17187_31287# a_17459_31145# a_17417_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18328 VDD a_10515_22671# a_17274_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18329 VDD a_76082_39738# a_75824_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1833 a_4499_65327# a_3983_65327# a_4404_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X18330 a_27710_20902# a_11067_67279# a_27314_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18331 a_23540_48981# a_23847_47919# a_23669_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X18332 VDD a_77002_40202# a_76744_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18333 VSS a_20195_49793# a_20156_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18334 a_1887_10749# a_1633_10422# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18335 a_5064_48841# a_3983_48469# a_4717_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18336 a_5135_50069# a_5147_50943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18337 a_22690_69222# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18338 a_9547_13103# a_9227_12015# a_9184_13255# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18339 a_2012_23805# a_1867_23983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1834 a_28607_29673# a_23192_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X18340 VDD a_2473_34293# a_4513_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18341 VSS a_30485_49257# a_30928_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18342 a_46786_23914# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18343 VDD a_24800_43041# a_34909_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X18344 a_17670_12870# a_10055_58791# a_17274_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18345 VDD a_5612_52520# a_5550_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18346 a_47486_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18347 VDD a_17300_51183# a_17475_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18348 VDD a_1643_57685# a_1591_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18349 vcm_commonmode a_16362_23548# a_24394_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1835 a_48490_57174# a_16746_57176# a_48398_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18350 a_2764_52271# a_1849_52271# a_2417_52513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18351 a_7653_72765# a_6224_73095# a_7571_72512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18352 a_23298_58178# a_16362_58178# a_23390_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18353 a_37354_71230# a_16362_71230# a_37446_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18354 VSS a_12895_13967# a_39758_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18355 a_36746_15882# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18356 VDD a_13835_36649# a_16648_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X18357 a_43774_16886# a_12727_13353# a_43378_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18358 VSS a_12727_15529# a_40762_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18359 result_out[14] a_1644_74005# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X1836 a_49798_18894# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18360 a_34342_9858# a_16362_9492# a_34434_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18361 a_4591_18543# a_4241_18543# a_4496_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18362 VSS a_16441_41781# a_16375_41807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18363 a_23298_17890# a_12899_10927# a_23790_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18364 a_11157_53609# a_11303_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18365 a_9063_71553# a_9314_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18366 a_24331_40767# a_22632_41831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X18367 VDD a_12899_10927# a_30326_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18368 a_30663_28585# a_30788_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18369 VDD a_10995_14333# a_10956_14459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1837 a_20682_24918# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18370 VSS a_19004_40413# a_18105_40157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X18371 a_31209_29673# a_28757_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18372 a_44474_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18373 a_4305_16189# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18374 VDD a_7387_64239# a_7758_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18375 a_31422_12504# a_16746_12502# a_31330_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18376 a_11400_26133# a_11251_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18377 a_43470_63198# a_16746_63200# a_43378_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18378 vcm_commonmode a_16362_60186# a_40458_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18379 vcm_commonmode a_16362_19532# a_40458_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1838 a_17274_23914# a_16362_23548# a_17366_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18380 a_44874_59504# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18381 vcm_commonmode a_16362_70226# a_23390_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18382 VSS a_19576_51701# a_19520_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18383 VSS a_4553_64213# a_4487_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18384 VDD a_10873_27497# a_16224_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18385 a_29718_59182# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18386 VSS a_26465_48463# a_27929_48579# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18387 a_29718_17890# a_12899_11471# a_29322_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18388 a_38044_44759# a_38140_44501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18389 VDD a_12901_66665# a_35346_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1839 vcm_commonmode a_16362_64202# a_28410_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18390 a_27314_16886# a_12899_11471# a_27806_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18391 a_4035_33205# a_4191_33449# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X18392 VSS a_10964_25615# a_17020_27253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X18393 a_10865_69679# a_10699_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18394 VDD a_11067_66191# a_12479_8545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18395 a_3487_73865# a_2971_73493# a_3392_73853# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X18396 VDD a_12727_58255# a_21290_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18397 a_18370_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18398 VSS a_12877_14441# a_17670_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18399 vcm_commonmode a_16362_61190# a_26402_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X184 VSS a_12899_11471# a_38754_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1840 VDD a_12546_22351# a_19282_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18400 a_4357_57961# a_4482_57863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18401 a_30418_18528# a_16746_18526# a_30326_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18402 a_12236_25321# a_9751_25071# a_12164_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18403 a_6361_57711# a_5823_57961# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18404 VSS a_7707_70741# a_9225_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18405 a_43538_31375# a_23395_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X18406 a_1952_60431# a_1775_60439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18407 a_22294_67214# a_12983_63151# a_22786_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18408 a_14679_31288# a_10531_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18409 a_33734_65206# a_10975_66407# a_33338_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1841 a_5065_66959# a_4211_67655# a_4983_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X18410 a_36336_42919# a_35463_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18411 a_30005_48463# a_29651_48576# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18412 VDD a_12447_29199# a_29498_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X18413 a_46786_64202# a_12355_65103# a_46390_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18414 a_12473_41781# a_30715_41835# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X18415 a_19877_52245# a_19591_50943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18416 a_37459_51183# a_37423_51335# a_37374_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18417 VDD a_12985_7663# a_44382_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18418 vcm_commonmode a_16362_14512# a_31422_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18419 conversion_finished_out a_1644_77813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X1842 a_34738_58178# a_12901_58799# a_34342_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18420 a_22690_22910# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18421 VSS a_17763_43413# a_17711_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18422 a_47486_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18423 a_19282_21906# a_16362_21540# a_19374_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18424 a_12341_69455# a_12135_69109# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18425 a_24755_42325# a_24931_42657# a_24883_42717# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X18426 VSS a_2497_53903# a_2882_54813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18427 a_42770_9858# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18428 VDD a_12677_36893# a_12283_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18429 VSS a_1586_40455# a_2235_41941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1843 a_27710_9858# a_12985_19087# a_27314_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18430 a_4717_45985# a_4499_45743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18431 a_36746_56170# a_12257_56623# a_36350_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18432 a_47790_7850# VDD a_47394_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18433 a_47790_72234# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18434 a_7101_55535# a_5254_67503# a_6646_54135# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18435 VDD a_12877_16911# a_34342_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18436 VSS a_13643_28327# a_28902_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18437 vcm_commonmode a_16362_67214# a_43470_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18438 a_19678_66210# a_12983_63151# a_19282_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18439 a_15892_51843# a_15261_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1844 a_33734_23914# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18440 a_1823_72381# a_2847_66389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18441 a_12132_51005# a_9240_53877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18442 a_5484_69455# a_4345_69679# a_5393_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X18443 a_9276_12167# a_9484_11989# a_9418_12015# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X18444 a_45478_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18445 VSS a_1586_21959# a_1591_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18446 a_1757_14741# a_1591_14741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18447 VSS a_12546_22351# a_28714_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18448 VSS a_12355_15055# a_41766_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18449 a_7337_42479# a_7293_42721# a_7171_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1845 a_41862_71552# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18450 a_9240_53877# a_11759_51959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18451 a_29322_57174# a_12257_56623# a_29814_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18452 a_38450_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18453 VDD a_6775_53877# a_10503_52828# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X18454 a_8021_53135# a_4339_64521# a_7519_59575# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18455 VSS VDD a_24698_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18456 a_20378_67214# a_16746_67216# a_20286_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18457 VDD a_34482_29941# a_37427_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18458 a_20734_46831# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18459 VSS a_4812_13879# a_5281_11791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1846 a_9821_46831# a_8566_39215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18460 a_39362_7850# VSS a_39454_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18461 a_4803_63669# a_4647_63937# a_4948_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18462 VDD VSS a_42374_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18463 a_21479_38053# a_19780_38341# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X18464 a_29718_12870# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18465 vcm_commonmode a_16362_58178# a_37446_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18466 a_12231_60949# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18467 a_1846_54699# a_2124_54715# a_2080_54813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18468 VSS a_12082_25077# a_12349_25847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18469 a_5731_13647# a_4812_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1847 a_15457_47081# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18470 a_49494_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18471 VSS a_1929_10651# a_5775_12649# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18472 VSS a_3247_20495# a_7153_18038# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18473 VDD a_10883_11177# a_11898_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18474 a_31726_61190# a_12355_15055# a_31330_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18475 VDD a_4443_46607# a_8275_43255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18476 VSS a_2223_28617# a_3801_24643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18477 a_11127_53544# a_11303_53511# a_11513_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18478 a_39362_22910# a_10515_23975# a_39854_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18479 a_43378_71230# a_12901_66665# a_43870_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1848 a_37846_61512# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18480 a_43870_20504# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18481 a_43470_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18482 VSS a_12981_62313# a_18674_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18483 a_25306_8854# a_12985_19087# a_25798_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18484 VDD a_12981_62313# a_46390_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18485 VDD a_5363_30503# a_7910_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18486 a_40218_27247# a_18979_30287# a_40132_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18487 vcm_commonmode a_16362_9492# a_44474_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18488 VDD a_2451_72373# a_8205_75369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18489 a_27406_57174# a_16746_57176# a_27314_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1849 VDD a_26417_47919# a_31186_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.6e+11p ps=5.72e+06u w=1e+06u l=150000u
X18490 a_28714_18894# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18491 a_19678_8854# a_12947_8725# a_19282_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18492 a_5337_23145# a_5211_24759# a_5265_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18493 a_33830_12472# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18494 VSS a_2012_68565# a_1586_69367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18495 VSS a_11619_63151# a_11987_67325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18496 a_31726_8854# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18497 VSS a_12899_11471# a_32730_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18498 a_32273_36161# a_30757_37455# a_32187_36161# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18499 a_38628_47349# a_38805_47081# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X185 a_35742_13874# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1850 a_45478_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18500 a_11067_13095# a_15103_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X18501 a_30418_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18502 a_20778_71552# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18503 a_47394_70226# a_12516_7093# a_47886_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18504 VDD a_11067_67279# a_20286_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18505 VSS a_26417_47919# a_28941_48801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18506 VDD a_12355_65103# a_19282_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18507 VSS a_12663_40871# a_13613_42134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18508 VDD a_7925_72399# a_9075_72737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18509 a_44382_12870# a_16362_12504# a_44474_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1851 a_36607_34191# a_36430_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18510 VDD a_12621_36091# a_36520_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X18511 VSS a_2606_41079# a_5077_46607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X18512 VSS a_1643_56597# a_1591_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18513 a_23390_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18514 a_20286_61190# a_16362_61190# a_20378_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18515 VSS a_12901_66959# a_44778_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18516 a_41766_66210# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18517 a_33430_24552# VDD a_33338_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18518 vcm_commonmode a_16362_63198# a_32426_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18519 a_23447_28853# a_23051_28023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1852 a_7862_34025# a_6372_38279# a_7444_34025# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X18520 a_33338_59182# a_12901_58799# a_33830_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18521 a_39305_48169# a_13643_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18522 a_30125_47919# a_26397_51183# a_30211_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X18523 vcm_commonmode a_16362_20536# a_43470_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18524 a_46482_23548# a_16746_23546# a_46390_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18525 VDD a_8489_74549# a_8379_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18526 a_24794_70548# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18527 a_45478_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18528 a_17274_14878# a_16362_14512# a_17366_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18529 VDD a_1952_60431# a_2635_55329# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1853 vcm_commonmode a_16362_56170# a_18370_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18530 a_21382_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18531 a_13795_39958# a_13613_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18532 a_21686_69222# a_12516_7093# a_21290_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18533 a_24302_60186# a_16362_60186# a_24394_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18534 VSS a_12727_67753# a_48794_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18535 a_12189_46805# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18536 a_45782_65206# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18537 a_29561_49667# a_29055_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18538 a_36442_15516# a_16746_15514# a_36350_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18539 a_11812_30511# a_11183_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X1854 a_38450_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18540 a_45878_17492# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18541 a_6614_74031# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18542 a_29926_30511# a_29942_30663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X18543 a_29987_47375# a_26397_51183# a_29847_48734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18544 a_43378_18894# a_16362_18528# a_43470_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18545 a_3301_16617# a_2283_15797# a_3229_16617# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X18546 a_20378_20536# a_16746_20534# a_20286_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18547 a_35438_8488# a_16746_8486# a_35346_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18548 a_32167_29611# a_33839_28309# a_33797_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18549 a_24800_44129# a_24515_43493# a_25447_43447# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1855 a_24302_71230# a_16362_71230# a_24394_71230# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18550 a_35742_57174# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18551 VDD a_12546_22351# a_27314_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18552 VSS a_27981_37477# a_28115_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18553 a_16902_50639# a_14985_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X18554 a_42770_58178# a_12901_58799# a_42374_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18555 a_7815_49855# a_7640_49929# a_7994_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18556 a_18674_67214# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18557 a_14092_52047# a_5190_59575# a_13925_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.86e+11p ps=2.18e+06u w=650000u l=150000u
X18558 a_45478_70226# a_16746_70228# a_45386_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18559 a_25702_68218# a_12901_66959# a_25306_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1856 a_26447_39141# a_25300_39655# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X18560 a_48794_56170# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18561 a_23141_52521# a_4891_47388# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X18562 VSS a_12355_65103# a_22690_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18563 vcm_commonmode a_16362_11500# a_37446_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18564 a_49894_16488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18565 a_46390_13874# a_12727_15529# a_46882_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18566 a_20378_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18567 a_36842_19500# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18568 a_40858_68540# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18569 a_35438_62194# a_16746_62196# a_35346_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1857 a_23694_15882# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18570 vcm_commonmode a_16362_8488# a_33430_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18571 VSS a_7377_18012# a_12713_20495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18572 VSS a_11067_13095# a_12710_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X18573 a_28361_51701# a_28143_52105# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18574 a_39758_14878# a_12727_15529# a_39362_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18575 a_18770_63520# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18576 VDD a_7862_34025# a_25299_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18577 a_28714_59182# a_12727_58255# a_28318_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18578 VSS a_12947_56817# a_25702_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18579 VDD a_12355_15055# a_22294_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1858 VSS a_12895_13967# a_26706_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18580 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18581 a_20378_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18582 VSS a_6752_29941# a_9019_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18583 VDD a_12727_13353# a_26310_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18584 VDD a_35615_30199# a_33839_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X18585 a_7171_42479# a_6725_42479# a_7075_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18586 a_44874_67536# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18587 a_41370_64202# a_11067_13095# a_41862_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18588 a_27406_10496# a_16746_10494# a_27314_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18589 a_2284_31287# a_1915_35015# a_2426_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1859 a_7755_70543# a_7289_70767# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=0p ps=0u w=650000u l=150000u M=4
X18590 a_32370_50871# a_2959_47113# a_32584_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=0p ps=0u w=1e+06u l=150000u
X18591 a_77285_39738# a_77381_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18592 a_44382_57174# a_16362_57174# a_44474_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18593 a_30722_62194# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18594 a_6739_59049# a_6361_57711# a_6521_58773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18595 a_27314_67214# a_16362_67214# a_27406_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18596 VSS VSS a_29718_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18597 VDD a_10391_49855# a_10378_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18598 a_24883_42717# a_12641_43124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18599 VDD a_1923_59583# a_4948_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X186 a_16746_21538# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X1860 a_35132_47695# a_34906_47491# a_34763_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18600 VSS a_10515_23975# a_44778_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18601 a_6807_36611# a_5631_38127# a_6735_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18602 a_17766_69544# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18603 a_2913_54991# a_2635_55329# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X18604 VSS a_35033_37692# a_34725_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18605 VDD a_12727_67753# a_21290_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18606 VSS a_8071_13255# a_7901_13077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18607 a_17274_59182# a_16362_59182# a_17366_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18608 a_31822_24520# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18609 a_7749_37903# a_3305_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1861 a_30722_16886# a_12727_13353# a_30326_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18610 a_21382_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18611 VSS a_3049_14343# a_2926_15253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18612 a_37750_17890# a_12899_11471# a_37354_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18613 a_12970_34191# a_12793_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18614 a_35346_55166# VSS a_35838_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18615 a_26748_7638# a_30891_28309# a_30663_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X18616 a_21686_22910# a_11067_21583# a_21290_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18617 VSS a_11067_21583# a_48794_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18618 VSS a_1586_51335# a_3891_50645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18619 a_18278_65206# a_12355_65103# a_18770_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1862 a_11619_56615# a_11067_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X18620 a_4161_37961# a_2971_37589# a_4052_37961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18621 vcm_commonmode a_16362_61190# a_34434_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18622 a_15207_30511# a_14361_29967# a_16494_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X18623 a_46786_72234# VDD a_46390_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18624 a_32334_20902# a_12985_7663# a_32826_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18625 a_32334_16886# a_16362_16520# a_32426_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18626 VSS a_20897_42917# a_22411_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X18627 VDD a_9989_46831# a_12489_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X18628 VDD a_12901_58799# a_42374_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18629 a_7201_56399# a_7169_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1863 VSS a_17039_51157# a_17365_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18630 vcm_commonmode a_16362_71230# a_17366_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18631 VSS a_12727_15529# a_38754_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18632 a_35742_10862# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18633 a_37888_43983# a_37711_43983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18634 a_30745_28111# a_18703_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18635 VDD a_23567_44211# a_23593_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X18636 a_42770_11866# a_12985_16367# a_42374_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18637 a_18674_20902# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18638 a_16228_28335# a_15599_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X18639 VSS a_8531_70543# a_34895_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1864 VDD a_7571_68047# a_4307_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.63335e+12p ps=2.328e+07u w=1e+06u l=150000u M=4
X18640 a_22294_12870# a_12877_16911# a_22786_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18641 a_25702_21906# a_12985_7663# a_25306_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18642 VSS a_3019_13621# a_4866_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18643 a_29791_52436# a_25419_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18644 VDD a_10515_22671# a_28318_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18645 a_16746_16518# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X18646 a_33825_32143# a_33694_30761# a_33741_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18647 a_33734_69222# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18648 a_17927_31573# a_4443_46607# a_18358_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X18649 vcm_commonmode VSS a_22386_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1865 VDD a_23901_35516# a_23507_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18650 VDD a_4351_26703# a_9135_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18651 a_6782_29967# a_7019_30511# a_6625_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18652 a_43319_31029# a_12907_27023# a_43538_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18653 a_28714_12870# a_10055_58791# a_28318_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18654 a_35346_72234# VSS a_35438_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18655 VSS a_12727_58255# a_37750_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18656 VSS a_11067_67279# a_37750_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18657 VSS a_32795_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X18658 VDD a_3325_18543# a_4627_27613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18659 a_26319_37429# a_13097_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1866 VDD a_14926_31849# a_23626_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18660 a_4298_58951# a_7815_49855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18661 a_25321_29673# a_2235_30503# a_25321_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18662 VDD a_33264_37601# a_32365_37692# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X18663 a_48398_71230# a_16362_71230# a_48490_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18664 result_out[0] a_1644_53877# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X18665 a_21290_18894# a_12895_13967# a_21782_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18666 VSS a_8201_62839# a_7619_62581# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18667 VSS a_22151_29941# a_22243_30491# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18668 a_18501_50645# a_18335_50645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18669 a_28410_18528# a_16746_18526# a_28318_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1867 a_2405_19087# a_2228_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18670 VDD a_11067_21583# a_38358_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18671 a_11987_67325# a_10379_66389# a_11881_67325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18672 vcm_commonmode a_16362_15516# a_25398_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18673 a_5691_36727# a_4685_37583# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X18674 VSS a_11400_26133# a_11430_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X18675 a_7461_27247# a_7113_27253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X18676 a_42466_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18677 a_8822_48829# a_2595_47653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18678 VDD a_15607_46805# a_35458_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18679 a_9408_25071# a_6559_22671# a_9218_25321# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1868 a_49494_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18680 a_25398_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18681 VSS a_10515_22671# a_31726_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18682 VSS a_26397_51183# a_32509_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X18683 a_14097_31375# a_8753_31055# a_14109_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X18684 a_41462_66210# a_16746_66212# a_41370_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18685 VDD a_16244_34973# a_16648_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X18686 a_34943_51335# a_35495_51157# a_35412_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X18687 a_3215_68351# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18688 a_43470_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18689 a_7010_39465# a_4941_35727# a_6927_39215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1869 a_42770_69222# a_12516_7093# a_42374_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18690 a_40366_21906# a_16362_21540# a_40458_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18691 vcm_commonmode a_16362_14512# a_29414_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18692 VDD a_19576_51701# a_22015_51840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18693 VSS a_10515_63143# a_14902_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18694 VDD a_12901_66665# a_46390_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18695 a_39454_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18696 a_36350_11866# a_16362_11500# a_36442_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18697 VSS a_3983_10927# a_1689_10396# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X18698 VDD a_9370_69831# a_9319_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18699 a_25306_19898# a_11067_67279# a_25798_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X187 a_2834_18909# a_1757_18543# a_2672_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1870 a_17462_51549# a_16385_51183# a_17300_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18700 a_46482_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18701 a_8215_31055# a_7460_31055# a_8297_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18702 a_10590_21263# a_10151_21379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X18703 a_6393_34837# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18704 a_2672_71689# a_1757_71317# a_2325_71285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18705 VSS a_6435_74005# a_6369_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18706 a_29414_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18707 a_22690_71230# a_12947_71576# a_22294_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18708 a_2672_9839# a_1591_9839# a_2325_10081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X18709 a_8133_52047# a_7933_51433# a_8051_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1871 VDD a_24800_35425# a_23901_35516# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X18710 VDD VDD a_19282_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18711 a_44382_20902# a_16362_20536# a_44474_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18712 VDD a_12947_8725# a_45386_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18713 VSS a_12985_19087# a_41766_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18714 a_19374_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18715 VSS a_10103_48682# a_9392_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X18716 a_33338_67214# a_12983_63151# a_33830_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18717 a_44778_65206# a_10975_66407# a_44382_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18718 a_9577_60437# a_9411_60437# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18719 a_27183_43493# a_23567_43123# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X1872 a_14293_39631# a_13867_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X18720 a_28747_37503# a_27981_37477# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X18721 a_18370_67214# a_16746_67216# a_18278_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18722 a_17187_31287# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18723 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18724 a_4906_60431# a_4148_60547# a_4343_60405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18725 a_48490_56170# a_16746_56172# a_48398_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18726 a_49798_17890# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18727 a_20682_23914# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18728 a_17274_22910# a_16362_22544# a_17366_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18729 VSS a_2873_13879# a_3049_14343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1873 a_31822_59504# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18730 VDD a_20713_36929# a_21800_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X18731 a_21382_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18732 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X18733 a_34738_57174# a_10515_22671# a_34342_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18734 a_27710_8854# a_12947_8725# a_27314_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18735 a_33734_22910# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18736 vcm_commonmode a_16362_68218# a_41462_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18737 VDD a_21057_30669# a_21012_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18738 VDD a_14983_51157# a_14859_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18739 VSS a_2235_30503# a_25368_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1874 a_27710_14878# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18740 a_10515_63143# a_12489_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X18741 VDD a_12907_27023# a_32867_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18742 VSS a_12899_10927# a_26706_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18743 a_4856_54991# a_4642_54991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18744 a_30722_15882# a_12877_14441# a_30326_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18745 a_43378_8854# a_16362_8488# a_43470_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18746 a_36442_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18747 VSS a_75162_39738# a_75111_39506# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18748 VDD a_7841_12167# a_7815_19319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18749 a_49494_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1875 vcm_commonmode a_16362_22544# a_37446_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18750 VSS a_21479_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X18751 a_10957_57711# a_10791_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18752 a_19282_8854# a_16362_8488# a_19374_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18753 VSS a_3607_34639# a_5547_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18754 VSS a_12381_43957# a_12325_44310# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18755 a_34062_47607# a_27535_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18756 VDD a_12516_7093# a_39362_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18757 a_31822_58500# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18758 a_27710_13874# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18759 a_2672_44655# a_1591_44655# a_2325_44897# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1876 a_46390_24918# VSS a_46882_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18760 VSS a_10055_58791# a_31726_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18761 a_29414_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18762 a_28410_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18763 a_18770_71552# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18764 a_39454_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18765 a_38499_37503# a_37733_37477# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X18766 a_36350_56170# a_16362_56170# a_36442_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18767 a_24794_7452# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18768 a_20682_7850# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18769 a_6619_16341# a_6444_16367# a_6798_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1877 a_18770_72556# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18770 vcm_commonmode a_16362_58178# a_48490_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18771 a_32649_28853# a_32038_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18772 a_2291_47753# a_1775_47381# a_2196_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X18773 a_43470_8488# a_16746_8486# a_43378_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18774 a_39758_66210# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18775 a_32802_32463# a_31691_32143# a_32507_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18776 a_27175_47375# a_22989_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18777 VSS a_11067_13095# a_43774_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18778 a_6882_15645# a_5805_15279# a_6720_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18779 VSS VDD a_30722_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1878 a_41462_20536# a_16746_20534# a_41370_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18780 a_37354_23914# a_12947_23413# a_37846_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18781 VSS a_2004_42453# a_2776_41167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18782 a_41370_72234# VDD a_41862_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18783 a_37354_19898# a_16362_19532# a_37446_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18784 a_41862_21508# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18785 a_31186_48169# a_26514_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18786 a_17774_28111# a_9529_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X18787 a_8123_34319# a_4685_37583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X18788 a_41462_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18789 a_29545_35841# a_29207_36415# a_30139_36649# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1879 a_36350_57174# a_16362_57174# a_36442_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18790 a_44382_65206# a_16362_65206# a_44474_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18791 VSS a_33641_29967# a_35049_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18792 VDD a_1586_21959# a_1591_21807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X18793 a_13180_29423# a_13143_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18794 VSS a_12947_56817# a_33734_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18795 VSS a_12981_62313# a_29718_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18796 a_26706_60186# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18797 a_25398_58178# a_16746_58180# a_25306_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18798 a_39454_71230# a_16746_71232# a_39362_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18799 a_26706_19898# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X188 a_2215_19997# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X1880 a_24794_8456# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18800 a_6007_23145# a_5991_21263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18801 a_16746_61192# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X18802 a_20682_64202# a_12355_65103# a_20286_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18803 VDD a_8295_47388# a_34342_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18804 VDD a_12877_14441# a_47394_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18805 a_40402_28111# a_18979_30287# a_40316_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18806 a_44874_12472# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18807 a_9576_32259# a_5346_33775# a_9355_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X18808 VSS a_10472_52423# a_9271_52789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18809 a_42374_13874# a_16362_13508# a_42466_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1881 VSS a_5599_74549# a_5557_74895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X18810 a_18370_20536# a_16746_20534# a_18278_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18811 a_21382_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18812 a_27806_22512# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18813 a_6825_29673# a_6649_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18814 a_21948_34973# a_21479_34239# a_22411_34473# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18815 a_17366_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18816 VDD a_11067_67279# a_31330_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18817 VDD a_8461_32937# a_13357_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X18818 a_17020_27253# a_12349_25847# a_16948_27253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18819 a_14482_27497# a_12349_25847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1882 a_20682_8854# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18820 a_7903_48841# a_7553_48469# a_7808_48829# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18821 a_31330_61190# a_16362_61190# a_31422_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18822 a_34738_10862# a_12546_22351# a_34342_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18823 a_9693_63695# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X18824 a_44474_24552# VDD a_44382_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18825 vcm_commonmode a_16362_21540# a_41462_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18826 a_17766_14480# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18827 a_5600_47919# a_4240_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18828 VDD a_10055_58791# a_21290_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18829 a_18370_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1883 a_36336_42919# a_36432_42919# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X18830 vcm_commonmode a_16362_66210# a_30418_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18831 VSS a_1923_54591# a_9425_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X18832 a_6093_67503# a_3143_66972# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18833 a_48890_11468# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18834 a_10964_25615# a_10521_25731# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18835 a_38850_68540# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18836 a_2215_45199# a_1591_45205# a_2107_45577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18837 VDD a_30052_32117# a_41141_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18838 a_32334_24918# VSS a_32426_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18839 a_1899_53387# a_1823_54973# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1884 VDD a_6795_51157# a_6671_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18840 a_12911_53609# a_12818_52521# a_12815_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18841 VDD a_12983_63151# a_42374_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18842 VDD a_2339_38129# a_2691_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18843 a_6141_16367# a_6097_16609# a_5975_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18844 a_28318_14878# a_16362_14512# a_28410_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18845 a_34434_16520# a_16746_16518# a_34342_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18846 a_20794_28335# a_15661_29199# a_20685_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18847 a_5612_52520# a_6985_52815# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X18848 a_2369_69501# a_2325_69109# a_2203_69513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18849 a_32426_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1885 VDD a_12901_66665# a_22294_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18850 a_7097_40303# a_6671_40630# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18851 a_6791_70455# a_7063_70313# a_7021_70339# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X18852 VSS a_16244_34973# a_15345_34717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X18853 vcm_commonmode VSS a_22386_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18854 VDD a_3295_62083# a_7963_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18855 a_47486_15516# a_16746_15514# a_47394_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18856 a_11885_67503# a_11053_69135# a_11803_67503# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18857 a_18278_10862# a_12985_16367# a_18770_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18858 VDD a_12985_16367# a_25306_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18859 a_32426_7484# VDD a_32334_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1886 a_40458_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18860 VSS a_34763_47349# a_34711_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18861 VSS a_8643_48767# a_8577_48841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18862 a_39362_64202# a_11067_13095# a_39854_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18863 a_46786_57174# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18864 VSS a_30311_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X18865 a_43870_62516# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18866 a_41059_29199# a_33641_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18867 a_10295_47919# a_9945_47919# a_10200_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X18868 a_42374_9858# a_12546_22351# a_42866_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18869 a_16648_37253# a_15775_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1887 a_7171_62313# a_7097_63151# a_7077_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X18870 vcm_commonmode a_16362_57174# a_24394_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18871 a_7189_35015# a_3607_34639# a_7352_35113# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18872 vcm_commonmode a_16362_11500# a_48490_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18873 a_47886_19500# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18874 a_31243_40183# a_30311_40229# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18875 a_27890_32459# a_5363_30503# a_27897_32219# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18876 a_15193_42917# a_15775_42405# a_16648_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X18877 a_21290_69222# a_16362_69222# a_21382_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18878 VDD a_12981_62313# a_20286_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18879 a_28810_9460# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1888 VDD a_12981_59343# a_18278_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18880 a_7571_20291# a_4792_20443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18881 a_29814_63520# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18882 a_2375_49172# a_2467_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X18883 VDD a_12139_71829# a_5877_70197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X18884 a_2012_18543# a_1895_18756# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18885 a_25398_11500# a_16746_11498# a_25306_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18886 a_13795_38870# a_13613_38870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18887 a_4274_60431# a_4148_60547# a_3870_60563# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X18888 VDD a_33385_46805# a_29760_55394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X18889 VSS a_5877_70197# a_5208_70063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1889 a_43470_9492# a_16746_9490# a_43378_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X18890 VDD a_12895_13967# a_24302_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18891 a_42374_58178# a_16362_58178# a_42466_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18892 a_17274_60186# a_12727_58255# a_17766_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18893 a_25306_68218# a_16362_68218# a_25398_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18894 a_11674_16367# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18895 a_37446_64202# a_16746_64204# a_37354_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X18896 a_42374_17890# a_12899_10927# a_42866_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18897 VSS a_12947_23413# a_42770_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18898 a_39454_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18899 a_27509_47695# a_22989_48437# a_27425_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X189 a_2672_45577# a_1591_45205# a_2325_45173# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X1890 a_39758_67214# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X18900 a_5021_70561# a_2952_66139# a_4935_70561# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X18901 VDD a_6559_22671# a_7431_22441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18902 a_8338_20969# a_7377_18012# a_8256_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X18903 a_33430_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18904 a_35742_18894# a_12899_10927# a_35346_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18905 a_3387_22390# a_2315_24540# a_2928_22583# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X18906 a_28318_59182# a_16362_59182# a_28410_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18907 vcm_commonmode a_16362_70226# a_42466_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18908 a_32426_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18909 a_48794_17890# a_12899_11471# a_48398_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1891 VSS a_12355_65103# a_43774_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18910 a_36324_34191# a_36147_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18911 VSS a_22259_48981# a_22193_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18912 a_2319_64476# a_2124_64507# a_2629_64239# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X18913 a_5173_44655# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18914 a_32730_64202# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18915 a_46390_55166# VSS a_46882_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18916 a_30326_21906# a_11067_21583# a_30818_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18917 a_29127_35561# a_28195_35327# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18918 a_2847_30271# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18919 a_30326_17890# a_16362_17524# a_30418_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1892 VSS a_12985_19087# a_30722_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X18920 VDD a_12727_58255# a_40366_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18921 VSS a_12877_14441# a_36746_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18922 vcm_commonmode a_16362_61190# a_45478_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18923 a_40491_27247# a_40218_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X18924 a_22690_56170# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18925 a_19282_18894# a_12895_13967# a_19774_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18926 VSS VSS a_19678_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18927 VSS a_34923_32375# a_17599_52263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18928 vcm_commonmode a_16362_71230# a_28410_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18929 a_2122_19087# a_1945_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1893 a_2325_19873# a_2107_19631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X18930 a_7553_69679# a_6921_72943# a_7469_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X18931 a_23790_16488# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18932 VSS a_12727_15529# a_49798_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18933 a_6467_55527# a_37534_51701# a_37478_52047# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X18934 a_20286_13874# a_12727_15529# a_20778_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18935 a_46786_10862# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18936 a_1915_35015# a_3983_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18937 a_1887_10422# a_1761_9295# a_1815_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X18938 VDD a_13047_29575# a_12999_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.85e+11p ps=2.57e+06u w=1e+06u l=150000u
X18939 VSS a_17039_51157# a_21781_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1894 a_23850_48463# a_23579_48463# a_23767_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18940 a_1644_71829# a_1591_63151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X18941 a_3705_40079# a_3663_39991# a_2927_39733# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X18942 vcm_commonmode a_16362_10496# a_24394_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18943 a_13143_29575# a_13241_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X18944 a_41697_27497# a_41334_29575# a_9135_27239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X18945 a_33338_12870# a_12877_16911# a_33830_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18946 a_32795_42943# a_31648_43781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X18947 a_38327_44759# a_34222_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18948 a_15828_38695# a_12889_39889# a_15970_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18949 a_22386_61190# a_16746_61192# a_22294_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1895 VDD a_12899_11471# a_43378_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18950 a_32003_35307# a_30757_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18951 vcm_commonmode a_16362_60186# a_49494_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18952 a_47394_7850# VDD a_47886_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18953 vcm_commonmode a_16362_19532# a_49494_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18954 VDD a_16510_8760# a_16746_8486# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X18955 a_26706_13874# a_12877_16911# a_26310_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18956 a_23450_51005# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18957 a_36746_9858# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18958 VDD a_5156_18543# a_5331_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18959 VDD a_9307_30663# a_10597_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1896 a_40858_14480# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18960 vcm_commonmode VSS a_33430_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18961 a_18753_27275# a_10873_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X18962 a_2629_72943# a_2250_73309# a_2557_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18963 a_46390_72234# VSS a_46482_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18964 a_27314_68218# a_12727_67753# a_27806_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18965 a_4717_20961# a_4499_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X18966 a_38754_66210# a_12983_63151# a_38358_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18967 a_12967_50943# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18968 a_31822_66532# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18969 a_26402_60186# a_16746_60188# a_26310_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1897 a_10667_74031# a_10221_74031# a_10571_74031# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X18970 a_29718_7850# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18971 a_24773_48463# a_24743_48437# a_24683_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X18972 vcm_commonmode a_16362_16520# a_23390_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18973 a_26402_19532# a_16746_19530# a_26310_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18974 VDD a_10515_23975# a_36350_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18975 a_36350_64202# a_16362_64202# a_36442_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18976 VDD a_11067_21583# a_49402_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18977 a_40458_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18978 a_34923_32375# a_18979_30287# a_35069_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X18979 vcm_commonmode a_16362_69222# a_35438_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1898 VSS a_7037_19385# a_6971_19453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18980 VSS VDD a_43774_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18981 VDD a_2589_62839# a_2099_64757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X18982 VDD a_7841_12167# a_8220_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18983 VSS a_1689_10396# a_2108_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18984 a_2518_23222# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18985 VSS a_75162_40202# a_75111_40050# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18986 a_15505_52521# a_15557_52245# a_8132_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X18987 a_32334_62194# a_12355_15055# a_32826_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X18988 VDD a_12727_15529# a_39362_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X18989 a_37446_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1899 a_41462_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18990 VSS a_1775_60663# a_2944_59893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X18991 a_2872_44111# a_2695_44119# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X18992 a_2325_51425# a_2107_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18993 a_16928_36391# a_15959_36415# a_16891_36649# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X18994 a_40762_7850# VDD a_40366_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18995 VSS a_5964_67655# a_5167_68060# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X18996 a_8015_21807# a_7571_22057# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X18997 a_6978_58487# a_7107_58487# a_7115_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18998 a_21879_30663# a_22243_30491# a_22178_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18999 a_12369_42693# a_12677_42333# a_12343_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X19 a_28703_29423# a_23928_28585# a_28513_29673# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X190 a_21382_72234# VDD a_21290_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1900 VSS a_29943_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X19000 a_7075_45577# a_6725_45205# a_6980_45565# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X19001 vcm_commonmode a_16362_68218# a_39454_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19002 a_20682_72234# VDD a_20286_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19003 a_2461_31599# a_2417_31841# a_2295_31599# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19004 VDD a_1923_59583# a_2464_63517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19005 a_14117_38341# a_14425_37981# a_13909_37571# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X19006 VSS a_3295_62083# a_3108_62043# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X19007 a_12831_39997# a_12651_39997# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19008 VSS a_12546_22351# a_21686_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19009 a_17366_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1901 a_8197_15279# a_7987_15431# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X19010 VSS a_2959_47113# a_30928_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19011 a_34738_60186# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19012 a_11711_32143# a_10515_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X19013 a_33430_58178# a_16746_58180# a_33338_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19014 a_34738_19898# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19015 vcm_commonmode a_16362_9492# a_38450_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19016 a_26118_51183# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19017 a_17670_70226# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19018 a_31726_9858# a_12985_19087# a_31330_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19019 VDD a_22995_30663# a_22151_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X1902 VSS a_19807_28111# a_32135_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X19020 a_38454_34191# a_38277_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19021 a_1849_33237# a_1683_33237# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19022 VDD a_15812_31029# a_7598_36103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X19023 a_46482_57174# a_16746_57176# a_46390_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19024 a_47790_18894# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19025 a_24331_39679# a_22448_39429# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X19026 a_29414_67214# a_16746_67216# a_29322_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19027 vcm_commonmode a_16362_64202# a_26402_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19028 a_10589_12879# a_10317_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19029 a_31726_23914# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1903 VDD a_1586_40455# a_5179_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19030 a_42466_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19031 a_28318_22910# a_16362_22544# a_28410_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19032 a_15683_40767# a_12343_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X19033 VDD a_28883_52031# a_28870_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19034 a_19594_35823# a_19417_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19035 VDD a_12355_65103# a_38358_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19036 a_35838_61512# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19037 VDD a_41636_37601# a_40737_37692# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X19038 a_32401_46831# a_20359_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19039 a_32426_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1904 VDD a_8273_42479# a_10730_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19040 a_36097_31375# a_33694_30761# a_35907_31055# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X19041 VSS a_4629_13647# a_6829_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19042 a_9481_24847# a_5449_25071# a_9043_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19043 a_19374_59182# a_16746_59184# a_19282_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19044 a_18370_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19045 a_22294_71230# a_16362_71230# a_22386_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19046 a_27710_62194# a_12981_62313# a_27314_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19047 VSS a_20543_46831# a_20661_47713# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19048 VSS a_12895_13967# a_24698_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19049 a_21686_15882# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1905 VSS a_12257_56623# a_33734_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19050 a_8539_47414# a_6559_22671# a_8080_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19051 a_5595_12167# a_5867_11995# a_5825_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19052 a_39362_72234# VDD a_39854_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19053 a_7805_69679# a_6921_72943# a_7721_69679# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X19054 a_23303_28335# a_14926_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19055 a_43870_70548# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19056 VDD a_27239_36341# a_13576_37149# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19057 a_16735_51183# a_16219_51183# a_16640_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X19058 a_39854_60508# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19059 a_9485_62613# a_9319_62613# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1906 a_12877_16911# a_11067_13095# a_12723_17231# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X19060 a_47486_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19061 a_40762_69222# a_12516_7093# a_40366_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19062 a_11096_10205# a_10659_9813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19063 a_32611_41317# a_31004_40743# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X19064 a_25702_14878# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19065 vcm_commonmode a_16362_22544# a_35438_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19066 a_16762_72556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19067 a_15397_39631# a_15131_39997# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19068 a_7539_63695# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19069 VDD a_12901_66665# a_20286_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1907 a_39454_72234# VDD a_39362_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19070 VDD a_2216_16885# a_2126_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.89e+11p ps=1.74e+06u w=420000u l=150000u
X19071 a_23390_9492# a_16746_9490# a_23298_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19072 a_29814_71552# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19073 a_37750_67214# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19074 VSS a_12875_31751# a_12215_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X19075 a_38837_46983# a_7295_44647# a_39000_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19076 a_17210_50639# a_14983_51157# a_16902_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19077 VSS a_12355_65103# a_41766_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19078 VDD a_2872_44111# a_19439_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X19079 a_21267_52047# a_20535_51727# a_21095_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X1908 VDD a_1823_67668# a_1775_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X19080 VDD a_12899_11471# a_41370_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19081 a_29322_61190# a_16362_61190# a_29414_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19082 VDD a_13975_44527# a_14081_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19083 VSS a_3325_69135# a_4906_67509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19084 a_33727_43177# a_32795_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19085 vcm_commonmode a_16362_21540# a_39454_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19086 a_48398_23914# a_12947_23413# a_48890_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19087 a_48398_19898# a_16362_19532# a_48490_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19088 a_28959_49783# a_28855_48801# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X19089 a_2781_66415# a_1591_66415# a_2672_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1909 a_4734_63695# a_4608_63811# a_4330_63827# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X19090 a_37446_72234# VDD a_37354_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19091 VSS a_2099_59861# a_2695_44119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19092 a_47790_59182# a_12727_58255# a_47394_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19093 VSS a_12947_56817# a_44778_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19094 a_38358_15882# a_12727_13353# a_38850_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19095 a_33430_11500# a_16746_11498# a_33338_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19096 VDD a_12727_13353# a_45386_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19097 a_42866_13476# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19098 VSS a_21021_46805# a_20955_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19099 VDD config_2_in[7] a_1591_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X191 a_42770_14878# a_12727_15529# a_42374_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1910 a_4345_32259# a_4157_32259# a_4263_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19100 VSS a_10975_66407# a_27710_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19101 VDD a_12895_13967# a_32334_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19102 a_31726_64202# a_12355_65103# a_31330_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19103 a_25798_23516# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19104 a_25398_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19105 a_6895_15253# a_6720_15279# a_7074_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19106 a_46482_10496# a_16746_10494# a_46390_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19107 a_29414_20536# a_16746_20534# a_29322_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19108 a_32426_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19109 a_2571_72040# a_2747_72007# a_2957_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1911 a_26267_34473# a_13484_39325# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X19110 VSS a_4075_64239# a_4167_64783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X19111 a_5670_22467# a_3339_43023# a_5588_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19112 a_21686_56170# a_12257_56623# a_21290_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19113 VDD a_12899_10927# a_18278_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19114 a_32730_72234# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19115 VSS a_11019_59575# a_10969_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19116 a_36842_69544# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19117 a_4440_57711# a_3016_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19118 a_19374_12504# a_16746_12502# a_19282_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19119 VDD a_7841_12167# a_9865_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1912 a_16746_62196# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X19120 VDD a_12727_67753# a_40366_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19121 a_26310_15882# a_16362_15516# a_26402_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19122 a_29414_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19123 VDD a_3143_22364# a_4165_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19124 a_30418_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19125 a_49894_68540# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19126 a_46482_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19127 a_19282_69222# a_16362_69222# a_19374_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19128 a_45478_16520# a_16746_16518# a_45386_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19129 a_20705_27791# a_15681_27497# a_20359_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1913 VSS a_12947_56817# a_46786_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19130 a_23390_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19131 a_25702_55166# VSS a_25306_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19132 a_4607_65693# a_3983_65327# a_4499_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19133 a_20713_39105# a_21387_38591# a_22260_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19134 a_23784_42583# a_23880_42325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19135 a_40762_22910# a_11067_21583# a_40366_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19136 VSS a_16744_40517# a_16265_39868# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X19137 a_37354_65206# a_12355_65103# a_37846_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19138 a_6655_46261# a_7090_46419# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19139 VDD a_12901_66959# a_26310_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1914 a_20682_65206# a_10975_66407# a_20286_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19140 vcm_commonmode a_16362_58178# a_22386_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19141 a_24591_31599# a_24716_31757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19142 VSS a_2292_43291# a_2860_43389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19143 a_10981_71311# a_2451_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19144 VDD a_6515_62037# a_7657_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19145 a_37750_20902# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19146 VSS a_1923_54591# a_1881_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19147 a_2375_13268# a_2313_12015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19148 VDD a_2325_10081# a_2215_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19149 a_35357_32463# a_35299_32375# a_34923_32375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1915 VDD a_12727_13353# a_47394_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19150 VDD a_10515_22671# a_47394_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19151 VSS a_12901_66665# a_35742_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19152 a_24302_22910# a_10515_23975# a_24794_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19153 a_7761_68047# a_5024_67885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19154 a_27806_64524# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19155 a_31871_51433# a_2775_46025# a_31669_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19156 VDD a_12981_62313# a_31330_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19157 a_22352_42693# a_21479_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19158 a_17670_23914# a_10515_23975# a_17274_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19159 a_16648_34215# a_15775_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1916 a_44874_13476# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19160 a_47790_12870# a_10055_58791# a_47394_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19161 a_17766_56492# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19162 a_9204_30663# a_8733_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X19163 VSS a_12516_7093# a_39758_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19164 a_5599_74549# a_6435_74005# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19165 a_35438_65206# a_16746_65208# a_35346_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19166 a_32334_70226# a_12516_7093# a_32826_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19167 a_44778_9858# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19168 a_11049_18543# a_10883_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19169 a_40366_18894# a_12895_13967# a_40858_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1917 a_41370_10862# a_12985_16367# a_41862_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19170 a_28318_60186# a_12727_58255# a_28810_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19171 VSS VSS a_40762_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19172 a_3856_70223# a_3588_70589# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19173 a_37446_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19174 a_2467_29397# a_2347_28918# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19175 VDD a_2497_53903# a_2882_54813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19176 vcm_commonmode a_16362_15516# a_44474_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19177 a_4615_40303# a_4578_40455# a_4446_40553# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19178 a_18487_28487# a_9529_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19179 a_33734_60186# a_12981_59343# a_33338_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1918 a_9135_27023# a_3607_34639# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=150000u
X19180 a_33734_19898# a_12895_13967# a_33338_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19181 a_35969_28111# a_35550_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19182 a_31422_23548# a_16746_23546# a_31330_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19183 VSS a_17039_51157# a_25461_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19184 a_44474_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19185 a_30418_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19186 a_14675_35831# a_15069_35805# a_14735_35805# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X19187 a_46786_18894# a_12899_10927# a_46390_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19188 a_19743_34743# a_18811_34789# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19189 vcm_commonmode a_16362_17524# a_17366_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1919 a_29667_31055# a_29416_31171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X19190 a_15775_41317# a_13097_40719# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X19191 a_30722_65206# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19192 a_21663_42943# a_20897_42917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X19193 VDD a_35815_31751# a_37287_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19194 a_21382_15516# a_16746_15514# a_21290_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19195 a_33101_36161# a_30757_37455# a_33015_36161# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X19196 a_30818_17492# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19197 a_44382_19898# a_11067_67279# a_44874_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19198 VDD a_2325_44897# a_2215_45021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19199 vcm_commonmode a_16362_62194# a_43470_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X192 a_36442_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1920 VSS a_10975_66407# a_29718_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19200 a_19678_61190# a_12355_15055# a_19282_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19201 a_6377_67503# a_6094_67825# a_5964_67655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19202 a_20682_57174# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19203 VSS a_8383_27247# a_9217_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19204 a_48490_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19205 vcm_commonmode VSS a_26402_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19206 a_76648_39738# a_76744_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19207 VSS a_12877_14441# a_47790_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19208 a_30418_70226# a_16746_70228# a_30326_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19209 VSS a_2292_17179# a_7493_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X1921 a_18370_21540# a_16746_21538# a_18278_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19210 VSS a_1803_20719# a_1945_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19211 VDD VDD a_38358_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19212 a_33734_56170# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19213 VDD a_9307_30663# a_10825_29688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19214 VDD a_12947_8725# a_39362_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19215 VSS a_12985_19087# a_35742_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19216 vcm_commonmode a_16362_11500# a_22386_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19217 a_31330_13874# a_12727_15529# a_31822_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19218 VDD a_5535_18012# a_8539_18231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19219 a_38450_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1922 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19220 a_21782_19500# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19221 a_8999_41974# a_8491_41383# a_8540_42167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19222 a_8853_61839# a_8999_61493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19223 a_16297_31849# a_2235_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19224 a_11507_18909# a_10883_18543# a_11399_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19225 a_20914_49551# a_20156_49667# a_20351_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19226 a_20378_62194# a_16746_62196# a_20286_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19227 a_27314_8854# a_12985_19087# a_27806_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19228 a_5725_21379# a_5671_21495# a_5629_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19229 vcm_commonmode a_16362_64202# a_34434_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1923 a_27806_23516# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19230 VSS a_6236_54421# a_6180_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19231 a_24698_14878# a_12727_15529# a_24302_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19232 a_17669_32509# a_17191_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19233 VSS a_10515_63143# a_12723_17231# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19234 a_33734_8854# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19235 a_7989_19425# a_5825_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19236 a_25306_69222# a_12901_66959# a_25798_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19237 a_49402_21906# a_16362_21540# a_49494_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19238 a_5695_47919# a_5179_47919# a_5600_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X19239 a_36746_67214# a_12727_67753# a_36350_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1924 a_4437_34639# a_2473_34293# a_4219_34551# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19240 a_13005_43983# a_12579_44310# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19241 a_2319_63388# a_2124_63419# a_2629_63151# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X19242 a_27333_32509# a_25953_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19243 a_6641_63401# a_6831_63303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19244 a_49798_66210# a_12983_63151# a_49402_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19245 a_3025_64783# a_1768_13103# a_2689_65103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X19246 a_12895_13967# a_11067_13095# a_12723_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X19247 a_20955_46831# a_12869_2741# a_20592_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X19248 VSS a_4792_20443# a_5825_20495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19249 VDD a_4553_64213# a_4583_64566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1925 VSS a_75445_40202# a_75258_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19250 a_26402_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19251 a_3229_26703# a_2223_28617# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19252 a_5909_51433# a_5135_50069# a_5909_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19253 a_3026_39037# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19254 VSS a_20964_31029# a_20911_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X19255 a_40585_42369# a_41167_42943# a_42099_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X19256 vcm_commonmode a_16362_69222# a_46482_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19257 a_10865_69679# a_10699_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19258 VSS a_4987_58229# a_4918_58255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19259 a_22690_17890# a_12899_11471# a_22294_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1926 a_48490_10496# a_16746_10494# a_48398_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19260 a_2122_20719# a_1945_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19261 VSS a_37888_43983# a_37994_43983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19262 a_20682_8854# a_12947_8725# a_20286_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19263 a_6752_29941# a_4248_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X19264 a_2101_10422# a_1929_10651# a_1887_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X19265 a_20286_55166# VSS a_20778_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19266 a_29718_23914# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19267 VDD a_1923_54591# a_2464_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19268 a_37446_8488# a_16746_8486# a_37354_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19269 a_41766_61190# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1927 a_27406_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19270 a_40458_59182# a_16746_59184# a_40366_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19271 a_27393_47919# a_26917_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.34e+11p pd=2.02e+06u as=0p ps=0u w=650000u l=150000u
X19272 a_38358_66210# a_16362_66210# a_38450_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19273 a_2656_42301# a_2539_42106# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19274 a_31726_72234# VDD a_31330_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19275 a_19678_15882# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19276 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19277 VSS a_12727_15529# a_23694_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19278 a_20682_10862# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19279 VSS a_13975_34191# a_14081_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1928 a_2751_42313# a_2401_41941# a_2656_42301# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X19280 a_6743_20969# a_3339_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19281 a_5729_36611# a_5691_36727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19282 a_75199_40594# a_75111_40050# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19283 VDD a_12447_29199# a_40387_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19284 a_7213_62215# a_7107_65871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19285 a_10289_55862# a_8132_53511# a_10075_55862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19286 VSS a_12981_62313# a_48794_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19287 a_45782_60186# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19288 a_4491_52854# a_4240_53083# a_4032_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19289 a_44474_58178# a_16746_58180# a_44382_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1929 a_6818_50959# a_4298_58951# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.46e+11p pd=5.58e+06u as=0p ps=0u w=650000u l=150000u M=2
X19290 vcm_commonmode VSS a_41462_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19291 a_45782_19898# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19292 a_28714_70226# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19293 a_27406_68218# a_16746_68220# a_27314_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19294 a_40133_48463# a_38067_47349# a_40050_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X19295 VSS a_9529_28335# a_14287_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19296 a_2830_15431# a_3019_13621# a_2965_13967# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19297 a_33830_23516# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19298 a_33430_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19299 VSS a_26345_40871# a_19919_38695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X193 a_23694_9858# a_12985_19087# a_23298_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1930 VDD a_12901_58799# a_34342_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19300 a_22386_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19301 a_26310_23914# a_16362_23548# a_26402_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19302 a_8475_44343# a_8143_44982# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19303 VDD a_10975_66407# a_36350_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19304 VSS a_7387_46831# a_7387_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X19305 VDD a_35602_34191# a_36147_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19306 VSS a_10339_14735# a_10673_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19307 a_16746_19530# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X19308 a_46882_22512# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19309 a_18674_62194# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1931 VDD a_12985_7663# a_31330_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19310 a_36442_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19311 VDD a_12355_65103# a_49402_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19312 a_20286_72234# VSS a_20378_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19313 a_25702_63198# a_15439_49525# a_25306_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19314 VSS a_12727_58255# a_22690_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19315 VSS a_11067_67279# a_22690_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19316 a_3693_68047# a_3215_68351# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19317 VDD a_4831_52413# a_4792_52539# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19318 VDD a_11611_12252# a_11542_12381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19319 a_16928_35303# a_15959_35327# a_16891_35561# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1932 a_11157_53609# a_11127_53544# a_10680_54171# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X19320 a_33338_71230# a_16362_71230# a_33430_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19321 a_36842_14480# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19322 a_36746_20902# a_11067_67279# a_36350_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19323 a_34342_15882# a_16362_15516# a_34434_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19324 VSS a_7071_62581# a_5428_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19325 VDD a_10055_58791# a_40366_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19326 VDD a_12257_56623# a_39362_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19327 a_36519_28879# a_32823_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19328 a_19774_24520# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19329 VDD a_11067_21583# a_23298_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1933 a_5064_45743# a_4149_45743# a_4717_45985# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X19330 VDD a_2847_40277# a_2834_40669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19331 a_10147_65984# a_9513_65301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19332 a_47394_14878# a_16362_14512# a_47486_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19333 a_4377_16189# a_3998_15823# a_4305_16189# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X19334 vcm_commonmode VSS a_16362_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19335 VSS a_30912_39429# a_30875_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19336 VSS a_4037_58773# a_3618_58487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19337 a_6929_53725# a_6666_53359# a_6516_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19338 a_34780_56398# a_34987_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19339 VSS a_10680_54171# a_8199_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X1934 a_4104_60431# a_3667_60405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19340 a_37354_10862# a_12985_16367# a_37846_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19341 a_6619_73719# a_5599_74549# a_6793_73825# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19342 vcm_commonmode a_16362_22544# a_46482_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19343 a_31280_36165# a_30311_35877# a_31184_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19344 a_27806_72556# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19345 a_35742_68218# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19346 VDD a_12985_7663# a_27314_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19347 a_36350_9858# a_12546_22351# a_36842_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19348 VDD a_12901_66665# a_31330_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19349 a_24394_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1935 VDD a_35676_49525# a_37307_51339# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19350 a_21290_11866# a_16362_11500# a_21382_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19351 a_12591_31029# a_7695_31573# a_12989_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19352 a_8143_44982# a_2787_32679# a_8143_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19353 a_10472_54135# a_10680_54171# a_10614_54269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19354 a_10379_66389# a_10391_67477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19355 a_27314_62194# a_16362_62194# a_27406_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19356 a_48794_67214# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19357 VSS a_11803_64239# a_11801_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19358 a_39454_17524# a_16746_17522# a_39362_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19359 a_4149_20719# a_3983_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1936 a_31330_62194# a_16362_62194# a_31422_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19360 a_31422_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19361 VDD a_2764_52271# a_2939_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19362 a_40458_12504# a_16746_12502# a_40366_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19363 VSS a_11145_60431# a_11341_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19364 VDD a_12877_16911# a_17274_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19365 VDD a_28841_29575# a_28607_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19366 a_3983_70767# a_2686_70223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19367 a_38754_59182# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19368 a_40366_69222# a_16362_69222# a_40458_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19369 VSS a_12257_56623# a_42770_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1937 a_34738_11866# a_12985_16367# a_34342_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19370 a_36350_16886# a_12899_11471# a_36842_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19371 a_28410_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19372 a_1945_16911# a_1908_17141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19373 VSS a_12983_63151# a_25702_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19374 a_48890_63520# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19375 a_8566_39215# a_8127_39465# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X19376 a_9914_68279# a_9513_65301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19377 VDD a_8468_48841# a_8643_48767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19378 a_44474_11500# a_16746_11498# a_44382_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19379 a_30716_51701# a_29361_51727# a_30939_52047# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X1938 VDD a_6795_51157# a_9963_50959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19380 a_11943_63125# a_12231_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19381 VSS a_7295_44647# a_39035_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X19382 VDD a_12895_13967# a_43378_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19383 a_27406_21540# a_16746_21538# a_27314_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19384 VDD a_43319_31029# a_43267_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19385 a_5259_39367# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19386 a_44382_68218# a_16362_68218# a_44474_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19387 VDD a_15439_49525# a_25306_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19388 VDD a_3983_12015# a_3983_12879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19389 a_17366_13508# a_16746_13506# a_17274_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1939 a_23694_56170# a_12257_56623# a_23298_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19390 a_12757_9295# a_12479_9633# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X19391 VDD a_12899_10927# a_29322_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19392 a_16746_64204# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X19393 a_47886_69544# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19394 a_9551_23145# a_7187_23439# a_9443_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19395 VDD a_32765_31287# a_31964_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X19396 VSS a_10515_22671# a_19678_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19397 a_16746_11498# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X19398 a_21782_9460# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19399 a_16666_55166# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 VSS a_12801_38517# a_24382_41629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1940 a_36629_27791# a_36459_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19400 a_11964_71855# a_10883_71855# a_11617_72097# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19401 a_11212_57711# a_6417_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19402 a_12815_19319# a_12672_18115# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19403 a_21382_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19404 a_47394_59182# a_16362_59182# a_47486_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19405 a_28789_50613# a_28968_50871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19406 a_11574_22869# a_12349_25847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X19407 VDD a_10860_47919# a_11035_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19408 VDD a_12985_19087# a_31330_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19409 VDD a_28524_47919# a_30735_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1941 VDD a_8772_63927# a_9649_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X19410 VDD a_12516_7093# a_24302_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19411 a_48398_65206# a_12355_65103# a_48890_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19412 VSS a_2847_38975# a_2781_39049# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X19413 VSS a_26550_40871# a_26345_40871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19414 a_18959_50639# a_18335_50645# a_18851_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19415 a_4918_52637# a_4792_52539# a_4514_52523# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X19416 vcm_commonmode VSS a_34434_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19417 a_24394_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19418 a_21290_56170# a_16362_56170# a_21382_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19419 VDD a_25300_39655# a_25204_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X1942 a_17766_15484# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19420 a_4227_73791# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19421 VSS VSS a_38754_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19422 a_35742_21906# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19423 vcm_commonmode a_16362_58178# a_33430_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19424 vcm_commonmode a_16362_71230# a_47486_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19425 VDD a_2685_59933# a_2785_60151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19426 VSS a_8273_42479# a_9367_29397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19427 a_24698_66210# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19428 a_38358_57174# a_12257_56623# a_38850_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19429 a_12161_31849# a_3339_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1943 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19430 a_42866_55488# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19431 a_48794_20902# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19432 a_22294_23914# a_12947_23413# a_22786_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19433 VDD a_17039_51157# a_17787_47349# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19434 a_22294_19898# a_16362_19532# a_22386_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19435 a_19333_48463# a_18907_48502# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19436 a_25798_65528# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19437 a_4187_60673# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19438 VDD a_12947_8725# a_47394_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19439 VSS a_12985_19087# a_43774_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1944 vcm_commonmode a_16362_67214# a_30418_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19440 a_32730_14878# a_12727_15529# a_32334_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19441 a_41462_61190# a_16746_61192# a_41370_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19442 a_28410_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19443 a_25306_55166# VSS a_25398_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19444 a_34579_50613# a_35403_50069# a_35349_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19445 a_8060_58799# a_7773_63927# a_7969_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19446 a_38754_12870# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19447 VDD a_26413_31055# a_28063_32193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19448 a_24394_71230# a_16746_71232# a_24302_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19449 a_3107_66237# a_1768_16367# a_2744_66103# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X1945 VDD a_12877_16911# a_21290_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19450 VSS a_9187_10901# a_8556_10357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19451 a_45782_13874# a_12877_16911# a_45386_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19452 VSS a_12985_16367# a_42770_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19453 a_4052_37961# a_3137_37589# a_3705_37557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X19454 a_2437_28309# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19455 a_28810_17492# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19456 a_25306_14878# a_12877_14441# a_25798_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19457 VSS a_12985_7663# a_25702_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19458 a_28714_23914# a_10515_23975# a_28318_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19459 a_36107_36965# a_34699_37683# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X1946 a_38850_69544# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19460 VDD a_3280_70501# a_3372_70197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19461 a_2375_76372# a_2361_74575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X19462 a_37553_46831# a_27535_30503# a_37427_47893# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19463 VDD a_7803_11703# a_7755_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X19464 VDD a_5363_30503# a_27387_32373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X19465 vcm_commonmode a_16362_16520# a_42466_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19466 a_1761_43567# a_1591_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19467 a_18674_15882# a_12877_14441# a_18278_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19468 a_7807_69455# a_7755_68591# a_7449_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X19469 a_28410_70226# a_16746_70228# a_28318_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1947 a_35346_66210# a_10975_66407# a_35838_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19470 VDD a_13909_37571# a_14117_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X19471 a_24209_48463# a_23767_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19472 VDD a_2235_30503# a_17415_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19473 a_29322_13874# a_12727_15529# a_29814_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19474 a_27345_50095# a_26155_50095# a_27236_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X19475 a_2426_36278# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X19476 a_42466_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19477 a_44778_60186# a_12981_59343# a_44382_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19478 a_45386_8854# a_16362_8488# a_45478_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19479 a_44778_19898# a_12895_13967# a_44382_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1948 VDD a_12727_67753# a_42374_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19480 a_23790_68540# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19481 a_40366_7850# VDD a_40858_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19482 a_18370_62194# a_16746_62196# a_18278_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19483 VDD a_22448_38341# a_22521_37692# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X19484 a_13867_39958# a_13837_39860# a_13795_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X19485 a_19774_58500# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19486 VDD a_5411_12791# a_5227_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X19487 VSS a_10055_58791# a_19678_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19488 a_34738_7850# VDD a_34342_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19489 a_41243_30080# a_32823_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1949 a_28318_15882# a_16362_15516# a_28410_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19490 a_16471_42134# a_15193_41781# a_16012_41959# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19491 vcm_commonmode a_16362_17524# a_28410_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19492 VSS a_7187_20719# a_7571_22057# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19493 a_11145_60431# a_10667_60735# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19494 a_32426_15516# a_16746_15514# a_32334_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19495 vcm_commonmode a_16362_63198# a_41462_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19496 a_16953_51425# a_16735_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X19497 a_6607_42167# a_6559_27907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X19498 a_37503_31393# a_32970_31145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19499 VDD a_33203_34191# a_33309_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X195 a_18674_23914# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1950 VSS a_3484_61493# a_2944_63400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X19500 a_26802_7452# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19501 a_22690_7850# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19502 a_24302_64202# a_11067_13095# a_24794_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19503 a_31726_57174# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19504 a_3162_53942# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X19505 VDD a_75728_39738# a_75541_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19506 VSS VDD a_32730_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19507 a_36442_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19508 VDD VDD a_49402_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19509 vcm_commonmode a_16362_11500# a_33430_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1951 a_21387_38591# a_19780_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X19510 VDD a_2713_31353# a_2743_31094# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19511 VSS a_18811_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X19512 a_49494_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19513 a_32826_19500# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19514 VSS a_9314_69367# a_10883_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19515 a_34342_23914# a_16362_23548# a_34434_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19516 VDD a_30599_28023# a_19720_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19517 a_48490_67214# a_16746_67216# a_48398_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19518 vcm_commonmode a_16362_64202# a_45478_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19519 VDD a_12546_22351# a_36350_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1952 a_32426_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19520 VDD a_2787_32679# a_5767_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19521 a_47394_22910# a_16362_22544# a_47486_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19522 a_7761_55785# a_7213_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X19523 VDD a_11067_67279# a_19282_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19524 a_34738_68218# a_12901_66959# a_34342_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19525 VSS a_30155_32375# a_23736_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19526 a_39758_61190# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19527 a_38450_59182# a_16746_59184# a_38358_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19528 vcm_commonmode a_16362_56170# a_35438_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19529 a_2437_28309# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1953 a_28115_43447# a_13835_43177# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X19530 a_22293_31171# a_15548_30761# a_22197_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19531 a_40762_15882# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19532 VSS a_12895_13967# a_43774_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19533 VSS a_4308_45431# a_4259_45199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19534 vcm_commonmode a_16362_66210# a_18370_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19535 a_14293_39631# a_13867_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19536 a_1761_31055# a_1591_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19537 a_22386_64202# a_16746_64204# a_22294_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19538 VDD a_2163_54589# a_2124_54715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19539 VDD a_2847_12863# a_2834_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1954 vcm_commonmode a_16362_8488# a_22386_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19540 VDD a_1689_10396# a_2101_10422# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19541 a_24394_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19542 a_30939_52047# a_2959_47113# a_30845_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X19543 VSS a_15775_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X19544 a_37761_44759# a_37857_44501# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19545 vcm_commonmode VSS a_39454_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19546 a_41059_32143# a_31659_31751# a_41141_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19547 a_20682_18894# a_12899_10927# a_20286_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19548 VDD a_7640_45577# a_7815_45503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19549 a_44778_14878# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1955 vcm_commonmode a_16362_59182# a_20378_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19550 vcm_commonmode VSS a_24394_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19551 a_27710_24918# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19552 a_17366_9492# a_16746_9490# a_17274_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19553 a_32217_28585# a_19807_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X19554 a_4263_32259# a_4157_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19555 a_36350_67214# a_16362_67214# a_36442_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19556 VDD a_12981_59343# a_35346_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19557 a_26447_38543# a_24413_39087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19558 a_48890_71552# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19559 a_31330_55166# VSS a_31822_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1956 VDD a_3143_66972# a_6927_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19560 VDD a_34759_31029# a_41243_30080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19561 a_1948_42479# a_1689_10396# a_1645_42453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X19562 a_16362_55166# VDD a_16270_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19563 a_17670_16886# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19564 VSS a_12877_14441# a_21686_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19565 a_44382_9858# a_12546_22351# a_44874_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19566 a_4522_34319# a_1915_35015# a_4219_34551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19567 vcm_commonmode a_16362_61190# a_30418_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19568 a_2601_72105# a_2747_72007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19569 a_40858_24520# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1957 a_47486_16520# a_16746_16518# a_47394_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19570 VSS a_8815_13879# a_8026_13885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X19571 a_15548_30761# a_10531_31055# a_16158_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19572 a_32611_39141# a_30912_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X19573 a_4365_64061# a_4330_63827# a_4127_63669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19574 a_13445_50639# a_12967_50943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19575 a_31726_10862# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19576 a_2375_34102# a_2011_34837# a_1916_33927# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19577 a_29207_36415# a_28441_36389# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X19578 a_1969_34863# a_1915_35015# a_1887_34863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19579 a_7257_73193# a_5599_74549# a_6835_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X1958 VDD a_35196_35425# a_36336_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X19580 VDD a_12947_71576# a_25306_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19581 VSS a_12983_63151# a_33734_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19582 a_20821_30511# a_20946_30669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19583 a_3173_46805# a_2656_45895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19584 VDD a_2529_24825# a_2559_24566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X19585 a_8569_24527# a_8031_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19586 a_4676_47607# a_4891_47388# a_4818_47414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19587 VSS a_10975_66407# a_46786_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19588 a_9187_51157# a_9390_51435# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19589 VDD a_4351_67279# a_15974_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1959 a_27710_55166# VSS a_27314_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19590 a_41370_20902# a_12985_7663# a_41862_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19591 a_44874_23516# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19592 a_7473_32259# a_6243_30662# a_7377_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19593 a_44474_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19594 a_41370_16886# a_16362_16520# a_41462_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19595 VDD a_7461_27247# a_9413_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19596 a_48490_20536# a_16746_20534# a_48398_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19597 a_4803_63669# a_4608_63811# a_5113_64061# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X19598 a_47486_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19599 a_19282_11866# a_16362_11500# a_19374_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X196 a_11067_21583# a_12516_7093# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X1960 a_8373_26409# a_7461_27247# a_8205_26159# VSS sky130_fd_pr__nfet_01v8 ad=2.21e+11p pd=1.98e+06u as=0p ps=0u w=650000u l=150000u
X19600 a_7925_72399# a_7571_72512# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19601 a_40762_56170# a_12257_56623# a_40366_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19602 VDD a_12899_10927# a_37354_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19603 a_31330_72234# VSS a_31422_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19604 a_1954_61677# a_4307_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19605 a_34834_15484# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19606 a_34738_21906# a_12985_7663# a_34342_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19607 a_24667_31055# a_24223_31171# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19608 VDD a_11067_46823# a_40783_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19609 a_23694_66210# a_12983_63151# a_23298_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1961 a_2325_29941# a_2107_30345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X19610 VSS a_37307_51339# a_37545_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19611 a_38450_12504# a_16746_12502# a_38358_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19612 a_47886_14480# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19613 a_11120_69679# a_8958_65961# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X19614 VDD a_10515_23975# a_21290_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19615 a_22595_35561# a_21663_35327# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19616 a_48490_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19617 a_45386_15882# a_16362_15516# a_45478_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19618 a_4591_18543# a_4075_18543# a_4496_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19619 a_26417_40193# a_25987_41317# a_26919_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X1962 a_18278_11866# a_10055_58791# a_18770_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19620 a_3026_49917# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19621 a_21290_64202# a_16362_64202# a_21382_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19622 a_40895_36919# a_41289_36893# a_25133_37571# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X19623 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19624 VDD a_12663_40871# a_13613_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X19625 vcm_commonmode a_16362_69222# a_20378_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19626 a_35346_11866# a_10055_58791# a_35838_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19627 a_3301_16617# a_2899_16367# a_3137_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X19628 a_27710_65206# a_10975_66407# a_27314_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19629 VDD a_12516_7093# a_32334_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1963 VDD a_14365_46805# a_11251_59879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u M=2
X19630 a_18278_21906# a_11067_21583# a_18770_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19631 a_18278_17890# a_16362_17524# a_18370_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19632 VDD a_12727_15529# a_24302_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19633 a_38883_29217# a_38210_30199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19634 a_12064_30287# a_12024_30199# a_11803_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19635 a_48398_10862# a_12985_16367# a_48890_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19636 a_22386_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19637 a_16287_38870# a_12889_39889# a_15828_38695# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19638 VDD a_12901_66959# a_45386_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19639 a_25306_63198# a_16362_63198# a_25398_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1964 a_38837_46983# a_8491_41383# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19640 a_46786_68218# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19641 a_37446_18528# a_16746_18526# a_37354_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19642 a_17670_57174# a_10515_22671# a_17274_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19643 a_2319_64476# a_2163_64381# a_2464_64605# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X19644 a_29733_48829# a_14831_50095# a_29651_48576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19645 VSS a_10286_26311# a_11400_26133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19646 vcm_commonmode a_16362_68218# a_24394_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19647 a_4341_62109# a_3295_62083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19648 a_10717_53113# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19649 VSS a_12447_29199# a_28113_29217# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1965 a_3854_29977# a_2216_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19650 VDD a_23565_38565# a_23685_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X19651 a_7837_68591# a_7707_70741# a_7755_68591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19652 a_4563_32900# a_5595_33205# a_5553_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19653 a_10570_67503# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19654 a_33830_65528# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19655 VDD a_12877_16911# a_28318_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19656 a_25019_37782# a_24837_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19657 a_25798_10464# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19658 VSS a_10515_22671# a_40762_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19659 a_1761_4399# a_1591_4399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1966 a_36520_38341# a_35647_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X19660 a_46882_64524# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19661 VDD a_7078_36103# a_7102_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19662 VSS a_7773_63927# a_7731_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19663 a_43378_61190# a_12981_59343# a_43870_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19664 VSS a_1586_9991# a_5179_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19665 vcm_commonmode a_16362_14512# a_38450_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19666 VDD a_1586_21959# a_10239_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19667 vcm_commonmode a_16362_59182# a_27406_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19668 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19669 VSS a_12985_7663# a_33734_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1967 a_32426_8488# a_16746_8486# a_32334_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19670 a_8251_39367# a_7910_38671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19671 a_31422_57174# a_16746_57176# a_31330_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19672 a_49402_7850# VDD a_49894_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19673 a_32730_18894# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19674 a_36842_56492# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19675 a_38754_9858# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19676 a_19774_66532# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19677 VDD a_12355_65103# a_23298_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19678 a_20778_61512# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19679 a_47394_60186# a_12727_58255# a_47886_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1968 a_42770_22910# a_11067_21583# a_42374_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X19680 a_19282_56170# a_16362_56170# a_19374_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19681 a_8994_63927# a_9643_63125# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19682 a_4149_20719# a_3983_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19683 a_2939_52245# a_2764_52271# a_3118_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19684 VDD a_24937_39306# a_12801_38517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X19685 a_13837_39860# a_13867_38870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19686 a_10138_26159# a_8373_26409# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19687 a_7458_10515# a_7775_10625# a_7733_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19688 a_24302_72234# VDD a_24794_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19689 a_16494_30511# a_10531_31055# a_15548_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1969 VSS a_28757_27247# a_30665_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.085e+11p ps=7.38e+06u w=650000u l=150000u M=2
X19690 VSS a_2656_70197# a_2686_70223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X19691 a_35742_70226# a_12901_66665# a_35346_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19692 VSS a_33939_43439# a_34045_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19693 VSS a_28963_28853# a_18611_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19694 VSS a_12135_69109# a_11985_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19695 VDD a_40581_31599# a_42941_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19696 a_24794_60508# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19697 a_32426_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19698 a_3870_60563# a_4187_60673# a_4145_60797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19699 a_2325_18785# a_2107_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X197 vcm_commonmode VSS a_47486_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1970 a_39362_65206# a_12355_65103# a_39854_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19700 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X19701 a_4883_33053# a_4259_32687# a_4775_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19702 vcm_commonmode a_16362_22544# a_20378_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19703 VDD VSS a_17274_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19704 a_38754_61190# a_12355_15055# a_38358_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19705 a_42770_7850# VDD a_42374_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19706 VSS a_12899_10927# a_35742_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19707 VSS a_1586_40455# a_1591_43029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19708 vcm_commonmode VSS a_45478_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19709 VDD a_6831_63303# a_28699_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1971 VSS a_9989_46831# a_11067_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X19710 a_13097_39631# a_12831_39997# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19711 a_22690_67214# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19712 VDD a_1586_9991# a_1591_12565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19713 VDD a_5913_48161# a_5803_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19714 VSS a_16257_38517# a_16191_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19715 a_49402_18894# a_12895_13967# a_49894_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19716 a_46786_21906# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19717 VSS VSS a_49798_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19718 a_17670_10862# a_12546_22351# a_17274_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19719 a_17774_27791# a_12631_28585# a_17774_28111# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X1972 a_40366_60186# a_12727_58255# a_40858_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19720 VSS a_12546_22351# a_23694_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19721 a_7203_71017# a_2843_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19722 vcm_commonmode a_16362_21540# a_24394_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19723 a_33338_23914# a_12947_23413# a_33830_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19724 a_5993_37039# a_5455_37039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19725 a_33338_19898# a_16362_19532# a_33430_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19726 a_40858_58500# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19727 VSS a_12899_11471# a_39758_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19728 a_36746_13874# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19729 a_22386_72234# VDD a_22294_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1973 a_46786_58178# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19730 VDD a_20359_29199# a_43353_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19731 a_43774_14878# a_12727_15529# a_43378_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19732 VSS a_10055_58791# a_40762_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19733 a_37446_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19734 a_6417_15279# a_6373_15521# a_6251_15279# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19735 a_7203_24527# a_7111_22351# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19736 a_34342_7850# VSS a_34434_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19737 VDD a_7571_31599# a_8197_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X19738 a_26802_18496# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19739 a_26706_24918# VSS a_26310_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1974 a_8856_64015# a_8772_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X19740 a_23298_15882# a_12727_13353# a_23790_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19741 VDD a_12727_13353# a_30326_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19742 a_27901_52513# a_27683_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19743 VDD a_9367_29397# a_9576_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19744 a_8275_43255# a_8383_43255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19745 a_44382_69222# a_12901_66959# a_44874_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19746 a_1644_66933# a_1823_66941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19747 vcm_commonmode a_16362_12504# a_27406_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19748 vcm_commonmode a_16362_63198# a_39454_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19749 a_44474_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1975 VDD a_12901_66959# a_28318_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19750 a_2284_36103# a_2216_28309# a_2426_36278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19751 a_42375_42089# a_41443_41855# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19752 a_31422_10496# a_16746_10494# a_31330_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19753 a_2012_21807# a_1867_21263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19754 VDD a_2840_66103# a_35224_49871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19755 a_2126_43023# a_1591_43029# a_2040_43401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19756 a_7676_61493# a_9735_63669# a_9693_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19757 a_29718_57174# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19758 a_3118_31599# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19759 a_29718_15882# a_12877_14441# a_29322_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1976 a_5147_50943# a_4972_51017# a_5326_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19760 a_25269_27791# a_24991_28129# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X19761 VDD a_24892_38237# a_23993_37981# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X19762 a_8497_56873# a_8123_56399# a_8082_56775# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X19763 a_52778_39198# a_52590_39198# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.66e+06u as=0p ps=0u w=500000u l=150000u M=2
X19764 a_5905_44655# a_5715_44343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19765 a_21782_69544# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19766 a_20286_8854# a_12985_19087# a_20778_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19767 a_12680_53511# a_12953_53339# a_12911_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19768 a_17766_59504# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19769 a_10961_19087# a_10791_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1977 VSS a_7925_72399# a_9225_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X19770 VDD a_9405_31599# a_10423_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19771 a_39431_43177# a_38499_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19772 a_5077_46607# a_4443_46607# a_4500_45289# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19773 a_29414_62194# a_16746_62196# a_29322_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19774 vcm_commonmode a_16362_18528# a_26402_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19775 a_12441_26409# a_9751_25071# a_12345_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19776 a_30818_8456# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19777 a_27239_36341# a_27415_36341# a_27367_36367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X19778 a_3020_54135# a_2913_54991# a_3162_53942# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19779 a_30418_16520# a_16746_16518# a_30326_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1978 a_6743_20969# a_4792_20443# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X19780 a_4214_37583# a_3137_37589# a_4052_37961# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19781 a_11957_67503# a_11710_58487# a_11885_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19782 VSS a_2847_49855# a_2781_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X19783 a_8357_44982# a_2787_32679# a_8143_44982# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19784 a_4242_35407# a_3803_35523# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X19785 a_22294_65206# a_12355_65103# a_22786_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19786 a_4789_58621# a_4311_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19787 a_43774_71230# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19788 a_42466_69222# a_16746_69224# a_42374_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19789 a_2781_39049# a_1591_38677# a_2672_39049# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1979 a_9361_28335# a_7281_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X19790 a_5813_39759# a_3949_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X19791 a_41370_24918# VSS a_41462_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19792 a_3031_47679# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19793 a_12231_55509# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19794 VSS a_8197_31599# a_11372_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19795 a_3203_17620# a_3063_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19796 a_22690_20902# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19797 a_47486_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19798 a_25306_56170# a_12947_56817# a_25798_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19799 a_34434_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X198 a_3280_70501# a_1586_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1980 vcm_commonmode a_16362_58178# a_24394_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19800 a_8367_44343# a_4443_46607# a_8541_44449# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19801 VSS a_12901_66665# a_20682_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19802 a_47790_70226# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19803 a_46482_68218# a_16746_68220# a_46390_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19804 a_6365_62063# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19805 VDD a_12985_16367# a_34342_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19806 vcm_commonmode a_16362_65206# a_43470_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19807 a_19678_64202# a_12355_65103# a_19282_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19808 a_8923_30287# a_8273_42479# a_8733_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19809 a_15162_32463# a_12412_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X1981 a_36708_39655# a_35739_39679# a_36612_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X19810 a_45386_23914# a_16362_23548# a_45478_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19811 a_2843_71829# a_2847_71615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X19812 a_13867_38870# a_13837_38772# a_13795_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X19813 a_37750_62194# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19814 VSS a_12727_58255# a_41766_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19815 VSS a_11067_67279# a_41766_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19816 a_29322_55166# VSS a_29814_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19817 a_14081_39958# a_13909_39747# a_13867_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X19818 VSS a_12516_7093# a_24698_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19819 a_49494_59182# a_16746_59184# a_49402_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1982 VSS a_1952_60431# a_3680_57527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X19820 vcm_commonmode a_16362_56170# a_46482_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19821 a_20378_65206# a_16746_65208# a_20286_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19822 a_22386_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19823 VDD a_7841_22895# a_11339_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19824 a_75728_40202# a_75824_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19825 a_38850_24520# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19826 VSS a_6095_44807# a_12289_54475# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19827 VSS a_4629_13647# a_5869_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19828 VDD a_11067_21583# a_42374_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19829 a_29718_10862# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1983 a_33830_55488# a_12869_2741# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19830 VSS a_3339_43023# a_3983_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19831 VDD a_3357_22649# a_3387_22390# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19832 a_48490_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19833 VSS a_12981_59343# a_27710_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19834 a_3668_10749# a_3417_10927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19835 VSS a_3693_68047# a_4906_67509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19836 VDD a_12727_15529# a_32334_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X19837 VDD a_9314_69367# a_10883_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19838 a_6737_60751# a_5024_67885# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19839 a_31726_18894# a_12899_10927# a_31330_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1984 a_2529_24825# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19840 VSS a_18811_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X19841 a_31031_47919# a_27869_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19842 VDD a_20359_29199# a_42801_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19843 a_39362_20902# a_12985_7663# a_39854_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19844 a_46882_72556# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19845 a_39362_16886# a_16362_16520# a_39454_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19846 a_10378_49551# a_9301_49557# a_10216_49929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19847 a_43470_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19848 a_40366_11866# a_16362_11500# a_40458_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19849 a_9325_29673# a_8383_27247# a_9135_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1985 a_11372_30511# a_10595_30511# a_11281_30511# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X19850 VDD a_12981_59343# a_46390_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19851 a_29322_72234# VSS a_29414_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19852 a_27406_55166# VDD a_27314_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19853 a_28714_16886# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19854 VDD a_6451_22895# a_7113_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19855 a_33830_10464# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19856 VSS a_12877_14441# a_32730_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19857 VSS a_13067_38517# a_12879_38517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19858 VDD a_2007_39978# a_1778_42631# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X19859 a_6750_19453# a_3247_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1986 a_39758_20902# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X19860 a_26310_10862# a_16362_10496# a_26402_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19861 a_42466_22544# a_16746_22542# a_42374_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19862 VDD VDD a_23298_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19863 a_2369_71677# a_2325_71285# a_2203_71689# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19864 VDD a_12981_62313# a_19282_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19865 a_19282_64202# a_16362_64202# a_19374_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19866 a_53260_40156# a_7841_12167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19867 a_23390_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19868 a_40861_30511# a_32970_31145# a_40773_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=0p ps=0u w=420000u l=150000u
X19869 VSS a_12983_63151# a_44778_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1987 VDD a_11619_3303# a_12171_3311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X19870 a_41766_64202# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19871 a_4607_46109# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19872 a_6671_40630# a_6559_39759# a_6599_40630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19873 a_6782_29967# a_5993_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19874 a_41141_32143# a_11067_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19875 a_46482_21540# a_16746_21538# a_46390_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19876 VSS a_27600_36165# a_27563_35831# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19877 VSS a_12901_58799# a_34738_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19878 a_1824_61127# a_1768_13103# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19879 a_17274_12870# a_16362_12504# a_17366_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1988 VSS a_15345_34717# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X19880 VSS a_12901_66959# a_17670_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19881 a_1761_41935# a_1591_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X19882 VSS a_8539_71829# a_8485_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19883 a_21686_67214# a_12727_67753# a_21290_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19884 a_13867_38543# a_13613_38870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19885 a_1757_19631# a_1591_19631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19886 VSS a_1586_45431# a_3983_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19887 a_36442_13508# a_16746_13506# a_36350_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19888 VSS a_9751_25071# a_11711_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19889 VDD a_12899_10927# a_48398_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1989 a_32029_41829# a_32611_41317# a_33543_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X19890 a_45878_15484# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19891 a_2672_66415# a_1757_66415# a_2325_66657# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19892 a_19374_23548# a_16746_23546# a_19282_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19893 a_10965_11177# a_10661_10383# a_10883_11177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X19894 a_2629_56623# a_2250_56989# a_2557_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19895 a_49494_12504# a_16746_12502# a_49402_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19896 a_5975_71829# a_5800_71855# a_6154_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X19897 VSS a_10515_22671# a_38754_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19898 a_35742_55166# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19899 a_35581_31599# a_29927_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X199 a_22294_15882# a_12727_13353# a_22786_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1990 a_5541_53609# a_1823_63677# a_5541_53359# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X19900 a_18674_65206# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19901 a_49402_69222# a_16362_69222# a_49494_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19902 vcm_commonmode a_16362_69222# a_31422_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19903 VSS a_17039_51157# a_26933_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19904 a_46390_11866# a_10055_58791# a_46882_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19905 a_36350_68218# a_12727_67753# a_36842_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19906 a_5213_70223# a_4935_70561# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X19907 VDD a_12516_7093# a_43378_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19908 a_40858_66532# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19909 VDD a_4215_51157# a_18335_50645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1991 VSS a_12901_66665# a_37750_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19910 a_35438_60186# a_16746_60188# a_35346_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19911 VDD a_12727_58255# a_39362_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19912 a_35438_19532# a_16746_19530# a_35346_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X19913 VSS a_3325_29967# a_3983_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19914 a_43470_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19915 a_40366_56170# a_16362_56170# a_40458_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19916 VSS a_23395_32463# a_28757_30539# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19917 a_27367_36367# a_12641_37684# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19918 a_19096_44129# a_18627_44581# a_19559_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X19919 VDD a_4298_58951# a_8051_52047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1992 a_30326_71230# a_12901_66665# a_30818_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19920 VDD a_11053_69135# a_11801_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19921 a_18770_61512# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19922 a_33656_43439# a_33479_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X19923 a_26402_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19924 a_23298_66210# a_16362_66210# a_23390_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19925 a_28714_57174# a_10515_22671# a_28318_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19926 a_3911_16065# a_1586_9991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19927 VSS a_2411_26133# a_2461_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19928 a_20195_49793# a_4191_33449# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X19929 VDD a_3339_30503# a_12591_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1993 a_23915_39126# a_23733_39126# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19930 a_7067_19126# a_6816_19355# a_6608_19319# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19931 VSS a_3949_41935# a_7948_38377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19932 VSS a_12985_19087# a_37750_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19933 a_40691_30511# a_34759_31029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19934 VSS a_22448_37253# a_22411_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X19935 a_44874_65528# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19936 a_41370_62194# a_12355_15055# a_41862_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19937 VDD config_1_in[15] a_1591_25071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X19938 a_2620_17277# a_2040_17289# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X19939 a_44382_55166# VSS a_44474_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1994 a_29814_64524# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19940 a_30722_60186# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19941 a_29322_8854# a_12985_19087# a_29814_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19942 a_30722_19898# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19943 a_43470_71230# a_16746_71232# a_43378_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19944 a_6641_67279# a_5682_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19945 a_34834_57496# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19946 a_7623_13621# a_8026_13885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19947 a_3881_15055# a_3023_16341# a_2873_13879# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19948 VSS a_11759_59575# a_11019_59575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19949 a_44382_14878# a_12877_14441# a_44874_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1995 a_26310_61190# a_12981_59343# a_26802_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19950 a_47790_23914# a_10515_23975# a_47394_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19951 VSS a_12985_7663# a_44778_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19952 a_17766_67536# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19953 VDD a_10975_66407# a_21290_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19954 a_47886_56492# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19955 a_6671_40303# a_6417_40630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19956 a_27314_24918# VSS a_27806_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19957 a_17274_57174# a_16362_57174# a_17366_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19958 a_31822_22512# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19959 a_2012_69501# a_1775_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1996 a_35438_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19960 a_21382_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19961 a_37750_15882# a_12877_14441# a_37354_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19962 VSS a_12877_16911# a_34738_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19963 a_39141_39655# a_39449_39868# a_13909_39747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X19964 VSS a_10515_23975# a_17670_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19965 a_23447_28853# a_23195_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19966 a_3629_16189# a_3594_15955# a_3391_15797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19967 a_21782_14480# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19968 a_21686_20902# a_11067_67279# a_21290_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19969 VSS a_2411_26133# a_2369_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1997 a_24746_31849# a_24716_31757# a_24674_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=5.72e+06u as=0p ps=0u w=1e+06u l=150000u
X19970 VDD a_12947_8725# a_40366_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19971 a_2479_50899# a_2419_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X19972 a_6909_51183# a_6795_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19973 VDD a_12257_56623# a_24302_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19974 a_27945_52271# a_27901_52513# a_27779_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19975 VSS a_21233_40956# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X19976 a_46786_70226# a_12901_66665# a_46390_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19977 vcm_commonmode a_16362_18528# a_34434_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19978 VSS a_13669_35253# a_13613_35606# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19979 VSS a_22632_42919# a_22595_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X1998 VSS a_12985_16367# a_33734_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X19980 a_38850_58500# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19981 a_32334_14878# a_16362_14512# a_32426_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19982 VSS a_6516_53511# a_6467_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X19983 a_20905_32143# a_7862_34025# a_20905_32463# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X19984 VDD a_1586_9991# a_5179_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X19985 a_3887_30083# a_3854_29977# a_3805_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X19986 VSS a_10055_58791# a_38754_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19987 a_14859_51183# a_13925_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19988 vcm_commonmode a_16362_17524# a_47486_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19989 a_26147_31171# a_13357_32143# a_26065_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1999 inn_analog a_8583_33551# ctopn VDD sky130_fd_pr__pfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7075e+12p ps=2.185e+07u w=1.9e+06u l=220000u M=4
X19990 a_2325_45173# a_2107_45577# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19991 a_36746_62194# a_12981_62313# a_36350_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19992 a_22690_8854# a_12947_8725# a_22294_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19993 a_22294_10862# a_12985_16367# a_22786_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19994 a_5924_69135# a_5295_69135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X19995 a_8969_42233# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19996 vcm_commonmode a_16362_22544# a_31422_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19997 VDD VSS a_28318_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X19998 a_19678_72234# VDD a_19282_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19999 a_20682_68218# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_26495_37429# a_13669_37429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20 a_2127_4943# a_1683_5059# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X200 a_48794_12870# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2000 a_4404_48829# a_4287_48634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X20000 a_39454_8488# a_16746_8486# a_39362_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20001 a_3070_66998# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20002 a_49798_61190# a_12355_15055# a_49402_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20003 a_13762_43222# a_13716_43047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20004 VSS a_30788_28487# a_32951_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20005 VSS a_5085_23047# a_7203_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20006 a_33734_67214# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20007 a_23749_36929# a_24055_36415# a_24928_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20008 a_24394_17524# a_16746_17522# a_24302_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20009 VSS a_4123_37013# a_2952_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2001 a_11981_57711# a_10791_57711# a_11872_57711# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20010 a_8065_59049# a_7773_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20011 a_28714_10862# a_12546_22351# a_28318_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20012 a_2529_24825# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X20013 a_35346_70226# a_16362_70226# a_35438_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20014 VDD a_34699_38771# a_34725_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20015 VSS a_14131_44135# a_13944_43957# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20016 a_32626_30083# a_26523_29199# a_32544_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20017 a_2835_62215# a_1952_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20018 VDD a_27600_36165# a_27504_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20019 a_23694_59182# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2002 a_19774_56492# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20020 VDD a_18579_27399# a_17278_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X20021 a_8195_16911# a_7571_16917# a_8087_17289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20022 a_21290_16886# a_12899_11471# a_21782_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20023 VSS a_31959_34751# a_31905_35073# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20024 a_8379_74575# a_7755_74581# a_8271_74953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20025 a_28410_16520# a_16746_16518# a_28318_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20026 VDD a_11067_67279# a_38358_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20027 a_19127_43439# a_18950_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20028 vcm_commonmode a_16362_13508# a_25398_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20029 VSS a_20715_41245# a_20655_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X2003 VSS a_4215_51157# a_22015_50645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20030 a_24394_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20031 a_38358_61190# a_16362_61190# a_38450_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20032 a_25971_52263# a_32038_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X20033 VDD a_2339_38129# a_5670_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20034 a_27710_58178# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20035 vcm_commonmode a_16362_66210# a_37446_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20036 VDD a_13143_29575# a_14289_29687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20037 a_41462_64202# a_16746_64204# a_41370_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20038 a_39362_24918# VSS a_39454_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20039 VDD a_4887_36495# a_5455_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2004 a_7188_39215# a_7078_36103# a_6927_39215# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X20040 a_43470_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20041 VSS a_2284_31287# a_2235_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20042 VDD a_27411_50069# a_27398_50461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20043 a_39454_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20044 a_3751_72373# a_4227_73791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X20045 a_39758_69222# a_12516_7093# a_39362_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20046 a_32826_69544# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20047 a_27406_63198# a_16746_63200# a_27314_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20048 vcm_commonmode VSS a_18370_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20049 a_40961_31375# a_32970_31145# a_40743_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2005 a_30125_47919# a_26514_47375# a_30039_47919# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X20050 VSS a_12901_66665# a_18674_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20051 VDD a_3143_66972# a_6737_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20052 VDD a_20747_27765# a_20705_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20053 a_32334_59182# a_16362_59182# a_32426_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X20054 a_10681_12559# a_9491_12297# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20055 a_16362_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20056 a_27247_43047# a_27271_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20057 VDD a_12901_66665# a_19282_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20058 a_41766_72234# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20059 a_10654_60431# a_9577_60437# a_10492_60809# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2006 a_4918_52637# a_4831_52413# a_4514_52523# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20060 a_19374_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20061 VDD a_3247_20495# a_6743_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X20062 a_14088_41807# a_12889_40977# a_13867_42134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X20063 a_33338_65206# a_12355_65103# a_33830_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20064 a_38358_9858# a_12546_22351# a_38850_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20065 VDD a_30835_38695# a_13669_38517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X20066 VDD a_13837_39860# a_16879_37999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20067 VDD clk_vcm a_77972_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20068 a_18370_65206# a_16746_65208# a_18278_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20069 a_34342_10862# a_16362_10496# a_34434_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2007 a_37446_65206# a_16746_65208# a_37354_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20070 VSS a_5671_21495# a_11887_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20071 VSS a_35932_41953# a_35033_42044# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X20072 VDD a_11067_67279# a_12901_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20073 a_7072_56053# a_3295_62083# a_7295_56399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20074 VSS a_2411_18517# a_10897_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20075 a_4918_58255# a_4831_58497# a_4514_58387# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20076 a_49798_15882# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20077 VSS VSS a_23694_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20078 a_5239_65301# a_5064_65327# a_5418_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X20079 a_20682_21906# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2008 a_8117_27497# a_5085_23047# a_8021_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20080 a_17274_20902# a_16362_20536# a_17366_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20081 vcm_commonmode a_16362_71230# a_32426_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20082 VDD a_2143_15271# a_9729_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20083 a_5140_71855# a_5023_72068# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20084 a_23298_57174# a_12257_56623# a_23790_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20085 a_2325_22049# a_2107_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20086 a_34738_55166# a_8295_47388# a_34342_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20087 VSS a_75475_38962# a_76180_38962# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20088 a_33734_20902# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20089 a_19684_42693# a_18811_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2009 a_42374_18894# a_12895_13967# a_42866_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20090 VSS a_1950_59887# a_2511_60431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20091 a_45478_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20092 VDD a_13669_39605# a_14081_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20093 VDD a_9705_11989# a_9735_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20094 a_75162_39738# a_75258_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20095 VDD a_1643_59317# a_1591_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20096 VSS a_12727_13353# a_26706_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20097 a_23694_12870# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20098 a_35742_63198# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20099 a_24573_41263# a_14293_41807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X201 VSS a_11067_21583# a_22690_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2010 VSS VSS a_42770_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20100 a_30722_13874# a_12877_16911# a_30326_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20101 VSS a_34711_47375# a_34987_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X20102 a_19131_39958# a_18949_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20103 a_13173_29673# a_13143_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20104 a_48794_62194# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20105 VDD a_6649_25615# a_8485_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20106 a_2199_33609# a_1849_33237# a_2104_33597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20107 a_33819_41001# a_32887_40767# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20108 a_31691_32143# a_31440_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X20109 a_6929_53725# a_7050_53333# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2011 a_39454_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20110 a_42770_66210# a_12983_63151# a_42374_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20111 a_6269_43567# a_5791_43541# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20112 a_27314_58178# a_10515_22671# a_27806_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20113 a_10789_74273# a_10571_74031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X20114 VDD a_10515_23975# a_40366_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20115 VDD a_12727_67753# a_39362_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20116 VSS a_6816_19355# a_7571_20291# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20117 a_27710_11866# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20118 a_3162_54269# a_2840_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20119 a_33591_32375# a_30788_28487# a_33741_32463# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2012 a_12369_40517# a_12249_43457# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X20120 a_40366_64202# a_16362_64202# a_40458_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20121 a_49894_24520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20122 a_8021_39221# a_7187_37583# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20123 a_39454_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20124 a_3026_30333# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20125 VSS a_2100_24759# a_2007_23957# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20126 a_4647_63937# a_1586_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20127 VSS a_12355_15055# a_25702_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20128 VDD a_9219_71285# a_9150_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20129 a_23790_9460# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2013 VDD a_12445_50613# a_12335_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X20130 a_12066_20175# a_5671_21495# a_11763_20407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20131 a_39758_64202# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20132 a_39758_22910# a_11067_21583# a_39362_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20133 a_37354_21906# a_11067_21583# a_37846_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20134 a_37354_17890# a_16362_17524# a_37446_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20135 a_41370_70226# a_12516_7093# a_41862_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20136 VDD a_12727_15529# a_43378_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20137 VSS a_30679_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X20138 a_41462_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20139 VSS a_33313_51157# a_33071_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X2014 a_36350_20902# a_16362_20536# a_36442_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20140 VDD VSS a_26310_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20141 VSS a_2595_47653# a_7337_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20142 a_44382_63198# a_16362_63198# a_44474_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20143 a_11461_14191# a_11082_14557# a_11389_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20144 a_2781_49929# a_1591_49557# a_2672_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20145 a_19203_39631# a_18949_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20146 a_40458_23548# a_16746_23546# a_40366_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20147 a_5685_56623# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20148 VSS a_11611_12252# a_11542_12381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20149 VDD a_12877_16911# a_47394_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2015 VDD a_12473_41781# a_12885_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20150 a_44874_10464# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20151 a_17274_65206# a_16362_65206# a_17366_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20152 a_14081_38870# a_13909_38659# a_13867_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20153 a_2672_71689# a_1591_71317# a_2325_71285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20154 a_21382_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20155 a_27806_20504# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20156 VSS a_12727_67753# a_42770_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20157 a_27406_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20158 a_10401_21379# a_7377_18012# a_10328_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20159 a_2847_21781# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2016 VSS a_12901_66959# a_31726_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20160 VSS a_2143_15271# a_9729_18870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20161 VSS a_11667_63303# a_11619_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20162 a_5797_21379# a_4792_20443# a_5725_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20163 a_19283_37737# a_18351_37503# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20164 vcm_commonmode a_16362_69222# a_29414_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20165 a_17766_12472# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20166 VSS a_2143_15271# a_10791_15529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20167 a_31330_9858# a_16362_9492# a_31422_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20168 vcm_commonmode a_16362_64202# a_30418_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20169 VDD a_12546_22351# a_21290_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2017 VSS a_11619_56615# a_12672_18115# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20170 a_3137_28111# a_2473_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20171 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20172 a_8739_28879# a_8206_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X20173 VDD a_7841_12167# a_53714_40254# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20174 a_7469_69679# a_7289_70767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20175 a_38850_66532# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20176 a_35346_63198# a_12981_62313# a_35838_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20177 VDD a_3668_56311# a_7871_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20178 a_32334_22910# a_16362_22544# a_32426_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20179 VSS a_25971_29967# a_25971_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2018 VDD a_7097_67655# a_5160_68315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X20180 VSS a_12901_58799# a_45782_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20181 VDD a_12355_65103# a_42374_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20182 a_28318_12870# a_16362_12504# a_28410_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20183 a_40581_31599# a_40233_31605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X20184 a_34434_14512# a_16746_14510# a_34342_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20185 a_24698_61190# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20186 a_23390_59182# a_16746_59184# a_23298_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20187 vcm_commonmode a_16362_56170# a_20378_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20188 VDD a_17187_31287# a_16087_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X20189 a_17366_24552# VDD a_17274_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2019 a_6816_19355# a_8827_17215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X20190 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20191 VSS a_15069_35805# a_14761_36165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20192 a_2571_68425# a_2125_68053# a_2475_68425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20193 a_47486_13508# a_16746_13506# a_47394_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20194 VDD a_12257_56623# a_32334_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20195 a_38784_42589# a_38499_42943# a_39431_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20196 a_7963_58255# a_8199_58229# a_8157_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20197 a_39362_62194# a_12355_15055# a_39854_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20198 VSS a_10515_22671# a_49798_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20199 a_43870_60508# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X202 a_25702_24918# VSS a_25306_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2020 a_17493_50639# a_16902_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20200 a_46786_55166# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20201 VSS a_20881_28111# a_24223_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20202 a_47394_8854# a_16362_8488# a_47486_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20203 a_42374_7850# VDD a_42866_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20204 vcm_commonmode VSS a_24394_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20205 VSS a_43680_29941# a_43624_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20206 VSS a_2606_41079# a_18653_48502# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20207 a_7725_31599# a_7695_31573# a_7653_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20208 a_36746_7850# VDD a_36350_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20209 VSS a_18627_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X2021 a_33430_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20210 VDD a_15851_27791# a_15941_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X20211 a_21290_67214# a_16362_67214# a_21382_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20212 a_26706_58178# a_12901_58799# a_26310_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20213 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20214 VDD a_12981_59343# a_20286_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20215 VDD a_76082_40202# a_75824_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20216 a_28810_7452# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20217 a_24698_7850# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20218 a_35069_32143# a_35299_32375# a_34923_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20219 a_29814_61512# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2022 a_35742_60186# a_12981_59343# a_35346_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20220 a_35438_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20221 a_15009_47919# a_14655_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20222 a_25263_44535# a_24331_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20223 VSS a_12546_22351# a_17670_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20224 VDD a_22749_50613# a_22639_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20225 a_17964_28111# a_10873_27497# a_17774_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20226 a_41418_29673# a_41334_29575# a_41335_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X20227 VDD a_4461_53113# a_4491_52854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20228 a_41462_72234# VDD a_41370_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20229 VSS a_10575_69439# a_10509_69513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2023 a_35742_19898# a_12895_13967# a_35346_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20230 a_38754_23914# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20231 a_42374_15882# a_12727_13353# a_42866_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20232 VSS a_11067_21583# a_42770_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20233 a_45782_24918# VSS a_45386_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20234 a_5169_13353# a_4429_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20235 a_39454_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20236 a_4514_52523# a_4831_52413# a_4789_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20237 VSS a_10975_66407# a_31726_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20238 a_45878_57496# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20239 a_7293_49525# a_7075_49929# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2024 a_6224_73095# a_9011_74879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X20240 vcm_commonmode a_16362_22544# a_29414_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20241 a_35742_16886# a_12727_13353# a_35346_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20242 a_2215_66781# a_1591_66415# a_2107_66415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20243 a_28318_57174# a_16362_57174# a_28410_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20244 a_32426_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20245 a_48794_15882# a_12877_14441# a_48398_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20246 VDD a_12899_10927# a_22294_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20247 VSS a_12877_16911# a_45782_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20248 a_16699_37999# a_13669_39605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20249 a_4717_20961# a_4499_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X2025 vcm_commonmode a_16362_20536# a_30418_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20250 a_23390_12504# a_16746_12502# a_23298_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20251 a_2417_33205# a_2199_33609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20252 a_32826_14480# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20253 a_11886_29967# a_6459_30511# a_11803_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X20254 VSS a_7067_30663# a_7019_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20255 a_28056_37253# a_27183_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20256 a_36842_59504# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20257 a_30326_15882# a_16362_15516# a_30418_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20258 a_2928_67191# a_3143_66972# a_3070_66998# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20259 a_13620_43047# a_13835_43177# a_13762_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2026 a_18674_70226# a_12901_66665# a_18278_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20260 a_48490_62194# a_16746_62196# a_48398_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20261 a_34613_31375# a_34759_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20262 vcm_commonmode a_16362_18528# a_45478_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20263 a_49894_58500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20264 a_6169_57711# a_4891_47388# a_5823_57961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20265 a_19282_16886# a_12899_11471# a_19774_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20266 a_35517_34954# a_4443_46607# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20267 a_34738_63198# a_15439_49525# a_34342_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20268 a_7115_58575# a_6417_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20269 a_12805_14441# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2027 a_32426_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20270 VSS a_10055_58791# a_49798_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20271 a_20286_11866# a_10055_58791# a_20778_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20272 a_4240_53083# a_6646_54135# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20273 a_13762_36694# a_13123_38231# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20274 VSS a_41842_27221# a_43003_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20275 VSS a_13669_37429# a_26495_37429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20276 VSS a_2847_30271# a_2781_30345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X20277 a_19374_9492# a_16746_9490# a_19282_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20278 a_11245_25321# a_11057_25077# a_11163_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20279 a_25296_40517# a_24423_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2028 a_11760_46983# a_11067_47695# a_11902_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X20280 a_33338_10862# a_12985_16367# a_33830_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20281 a_4073_50095# a_4031_50247# a_3983_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X20282 VDD a_32371_32117# a_23395_52047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20283 vcm_commonmode a_16362_61190# a_18370_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20284 VDD a_12901_66959# a_30326_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20285 a_31726_68218# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20286 a_22386_18528# a_16746_18526# a_22294_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20287 VDD a_12901_58799# a_26310_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20288 a_37594_50755# a_36821_50095# a_37512_50755# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20289 VSS a_29269_44545# a_30323_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X2029 a_46482_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20290 a_27236_50095# a_26321_50095# a_26889_50337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20291 a_26706_11866# a_12985_16367# a_26310_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20292 a_1915_24148# a_2007_23957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X20293 a_10045_50959# a_4298_58951# a_9963_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20294 VDD a_1586_69367# a_5179_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X20295 VSS a_19311_35823# a_19417_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20296 a_12231_65301# a_1950_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20297 a_44382_56170# a_12947_56817# a_44874_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20298 a_46390_70226# a_16362_70226# a_46482_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20299 a_11942_70045# a_10865_69679# a_11780_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X203 a_19374_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2030 VDD a_21041_37429# a_21071_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20300 a_27314_66210# a_10975_66407# a_27806_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20301 a_38754_64202# a_12355_65103# a_38358_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20302 a_31822_64524# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20303 VDD a_12985_7663# a_36350_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20304 vcm_commonmode a_16362_14512# a_23390_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20305 a_10521_25731# a_10570_25625# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20306 a_13975_44527# a_13798_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20307 VSS a_9271_52789# a_9217_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X20308 VDD a_5135_50069# a_4127_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20309 a_39454_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2031 a_10509_69513# a_9319_69141# a_10400_69513# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20310 a_36350_62194# a_16362_62194# a_36442_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20311 a_3877_57167# a_3521_57283# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20312 a_27509_47695# a_27175_47375# a_27425_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=0p ps=0u w=1e+06u l=150000u
X20313 VDD a_1642_18231# a_1591_17999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20314 a_40458_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20315 VDD a_11067_67279# a_49402_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20316 a_21782_56492# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20317 a_39758_72234# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20318 vcm_commonmode a_16362_67214# a_35438_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20319 VDD a_20881_28111# a_23553_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2032 a_48794_18894# a_12899_10927# a_48398_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20320 VSS a_12516_7093# a_43774_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20321 a_8082_56775# a_7773_63927# a_8219_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20322 a_12473_37429# a_30991_35307# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X20323 a_32334_60186# a_12727_58255# a_32826_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20324 VDD a_10055_58791# a_39362_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20325 a_41462_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20326 vcm_commonmode a_16362_66210# a_48490_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20327 VDD a_6269_43567# a_6579_42255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X20328 a_10761_29745# a_10825_29688# a_10607_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20329 VDD a_5239_45717# a_5226_46109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2033 VSS a_12727_13353# a_45782_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20330 a_37446_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20331 VDD a_5963_20149# a_8999_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X20332 VSS a_12355_15055# a_33734_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20333 a_8017_36495# a_7479_36495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20334 a_30007_38695# a_26433_39631# a_30181_38571# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X20335 a_2275_28918# a_2093_28918# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20336 a_20103_30287# a_14625_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20337 a_20682_70226# a_12901_66665# a_20286_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20338 VSS a_12981_59343# a_46786_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20339 a_42466_56170# a_16746_56172# a_42374_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2034 vcm_commonmode a_16362_17524# a_19374_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20340 a_43774_17890# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20341 a_4514_52523# a_4792_52539# a_4748_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20342 VSS a_12901_66665# a_29718_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20343 a_25398_66210# a_16746_66212# a_25306_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20344 a_35959_30485# a_35815_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20345 a_27406_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20346 a_19500_34215# a_18627_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20347 a_12713_41923# a_15683_40767# a_16615_41001# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20348 VDD a_15439_49525# a_34342_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20349 a_4425_29673# a_2216_28309# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2035 a_32730_65206# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20350 a_10833_74031# a_10789_74273# a_10667_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20351 VDD a_7917_13885# a_7623_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20352 VDD a_2292_17179# a_4212_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20353 VDD a_17039_51157# a_20496_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20354 a_13762_36367# a_13123_38231# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20355 a_23694_61190# a_12355_15055# a_23298_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20356 VSS a_12899_10927# a_20682_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20357 a_46482_55166# VDD a_46390_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20358 a_47790_16886# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20359 a_1757_51183# a_1591_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2036 VDD a_12985_19087# a_19282_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20360 vcm_commonmode VSS a_30418_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20361 VDD a_10382_58487# a_10331_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20362 a_45386_10862# a_16362_10496# a_45478_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20363 a_35346_71230# a_12901_66665# a_35838_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20364 a_29414_65206# a_16746_65208# a_29322_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20365 VDD VDD a_42374_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20366 a_31726_21906# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20367 a_28318_20902# a_16362_20536# a_28410_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20368 VDD a_12981_62313# a_38358_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20369 a_2107_30345# a_1757_29973# a_2012_30333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2037 a_23390_15516# a_16746_15514# a_23298_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20370 a_41462_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20371 a_3417_31599# a_2939_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20372 a_19374_57174# a_16746_57176# a_19282_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20373 a_27710_60186# a_12981_59343# a_27314_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20374 a_27710_19898# a_12895_13967# a_27314_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20375 VSS a_12899_11471# a_24698_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20376 a_21686_13874# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20377 a_22386_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20378 a_39362_70226# a_12516_7093# a_39854_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20379 a_7657_64489# a_7567_64391# a_7439_64213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2038 VSS a_5775_12649# a_5411_12791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X20380 a_46786_63198# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20381 a_5173_20719# a_3983_20719# a_5064_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20382 a_4702_32143# a_4263_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X20383 VSS a_12901_66959# a_36746_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20384 VSS a_2163_54589# a_2124_54715# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20385 a_8815_13879# a_9083_13879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20386 a_40762_67214# a_12727_67753# a_40366_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20387 vcm_commonmode a_16362_63198# a_24394_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20388 VDD a_18126_28023# a_17691_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20389 VSS a_9123_55223# a_3780_56347# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2039 vcm_commonmode a_16362_12504# a_20378_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20390 a_25306_59182# a_12901_58799# a_25798_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20391 a_49402_11866# a_16362_11500# a_49494_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20392 a_12713_36483# a_24515_34789# a_25388_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20393 VSS a_18197_44220# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X20394 VDD a_2672_36873# a_2847_36799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20395 VSS a_23487_49007# a_23579_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X20396 a_2080_73309# a_1643_72917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20397 a_38450_23548# a_16746_23546# a_38358_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20398 vcm_commonmode a_16362_20536# a_35438_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20399 a_37446_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X204 VSS a_1824_61127# a_1775_60663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2040 a_31330_9858# a_12546_22351# a_31822_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20400 a_30908_44869# a_30035_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20401 a_37750_65206# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20402 a_4503_51017# a_4057_50645# a_4407_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20403 a_2944_64488# a_5274_62313# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X20404 a_37846_17492# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20405 a_26402_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20406 VDD a_12877_14441# a_41370_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20407 a_35346_18894# a_16362_18528# a_35438_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20408 a_8113_24847# a_6162_28487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20409 VDD a_8399_49159# a_8399_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2041 a_2215_22173# a_1591_21807# a_2107_21807# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X20410 a_8540_42167# a_8491_41383# a_8682_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20411 VDD a_16441_41781# a_16471_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20412 a_48398_21906# a_11067_21583# a_48890_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20413 a_48398_17890# a_16362_17524# a_48490_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20414 VDD a_13669_38517# a_14081_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20415 a_37446_70226# a_16746_70228# a_37354_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20416 a_17670_68218# a_12901_66959# a_17274_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20417 a_42374_66210# a_16362_66210# a_42466_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20418 a_47790_57174# a_10515_22671# a_47394_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20419 a_38358_13874# a_12727_15529# a_38850_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2042 a_32826_17492# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20420 a_42866_11468# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20421 VSS a_11067_13095# a_27710_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20422 a_7815_42453# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20423 VDD a_12215_31573# a_14747_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X20424 VDD a_16152_43677# a_15253_43421# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X20425 a_25798_21508# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20426 a_25398_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20427 a_28318_65206# a_16362_65206# a_28410_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20428 VDD a_8123_56399# a_9557_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20429 a_21021_46805# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2043 a_11587_55535# a_11141_55535# a_11491_55535# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X20430 a_32426_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20431 a_12541_20719# a_7377_18012# a_12263_20969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X20432 VDD a_10901_54201# a_10931_53942# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20433 VSS a_12947_56817# a_17670_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20434 a_8569_49007# a_8399_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X20435 VDD a_12727_13353# a_18278_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20436 a_32730_70226# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20437 a_31422_68218# a_16746_68220# a_31330_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20438 a_9217_29423# a_7841_29673# a_9135_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20439 a_36842_67536# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2044 a_20925_44007# a_21233_44220# a_20899_44211# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X20440 a_19374_10496# a_16746_10494# a_19282_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20441 a_25517_37455# a_25091_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20442 a_30326_23914# a_16362_23548# a_30418_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20443 a_7749_55535# a_7803_55509# a_7761_55785# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20444 VDD a_10975_66407# a_40366_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20445 a_26310_13874# a_16362_13508# a_26402_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20446 a_2215_38671# a_1591_38677# a_2107_39049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20447 VDD a_14963_39783# a_14951_39997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20448 a_49894_66532# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20449 a_46390_63198# a_12981_62313# a_46882_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2045 a_30326_18894# a_16362_18528# a_30418_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20450 a_22690_62194# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20451 a_46482_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20452 a_22365_31171# a_2787_30503# a_22293_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20453 a_19282_67214# a_16362_67214# a_19374_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20454 VDD a_4584_20407# a_3799_20407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20455 a_9468_55311# a_8123_56399# a_9278_55311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20456 a_45478_14512# a_16746_14510# a_45386_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20457 a_49402_56170# a_16362_56170# a_49494_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20458 VSS a_10515_23975# a_36746_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20459 VSS a_4351_67279# a_15892_51843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2046 a_35036_34191# a_34859_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20460 VDD a_12947_8725# a_34342_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20461 vcm_commonmode a_16362_56170# a_31422_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20462 a_10244_26159# a_10286_26311# a_10055_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X20463 a_23628_35823# a_23451_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20464 a_22632_41831# a_21663_41855# a_22595_42089# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X20465 a_40762_20902# a_11067_67279# a_40366_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20466 VSS a_7281_29423# a_7725_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20467 VDD a_12257_56623# a_43378_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20468 a_23790_24520# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20469 VDD a_12983_63151# a_26310_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2047 a_24375_47753# a_23929_47381# a_24279_47753# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X20470 a_22294_8854# a_12985_19087# a_22786_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20471 a_10472_52423# a_10680_52245# a_10614_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20472 a_11753_55535# a_11709_55777# a_11587_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20473 VSS a_11311_74005# a_8003_72917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20474 VSS a_11711_12559# a_12174_12381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20475 VSS a_18487_28487# a_18126_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X20476 a_26402_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20477 a_4499_20719# a_4149_20719# a_4404_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20478 VSS a_6775_53877# a_8021_53135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20479 a_75475_40594# a_75199_40594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2048 VDD a_8305_16885# a_8195_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X20480 VSS a_27195_32375# a_27167_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20481 a_32826_8456# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20482 a_10239_74575# a_10109_73487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20483 a_41599_28335# a_20635_29415# a_41261_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20484 a_28756_7638# a_22291_29415# a_32217_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20485 a_8999_22351# a_8933_22583# a_8891_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20486 a_38754_72234# VDD a_38358_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20487 VDD VSS a_47394_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20488 a_24302_20902# a_12985_7663# a_24794_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20489 a_31822_72556# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2049 a_14079_43222# a_13005_43983# a_13620_43047# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X20490 a_24302_16886# a_16362_16520# a_24394_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20491 VDD a_2040_17289# a_2216_16885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20492 VDD a_11151_14428# a_11082_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20493 a_25091_37782# a_25133_37571# a_25091_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20494 a_27806_62516# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20495 VSS a_13669_38517# a_14088_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20496 a_5909_51183# a_3325_49551# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20497 VDD a_12981_59343# a_31330_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20498 a_43470_17524# a_16746_17522# a_43378_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20499 a_17670_21906# a_12985_7663# a_17274_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 a_4238_55123# a_4555_55233# a_4513_55357# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X2050 vcm_commonmode a_16362_62194# a_45478_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20500 a_42721_28879# a_11067_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20501 a_9643_49334# a_9392_48981# a_9184_49159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20502 a_47790_10862# a_12546_22351# a_47394_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20503 VSS a_2021_17973# a_27359_43985# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20504 VSS a_1586_21959# a_10239_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20505 VDD a_2345_33749# a_2375_34102# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20506 VDD a_8275_43255# a_8171_43541# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X20507 a_15959_35327# a_14735_35805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X20508 a_42770_59182# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20509 a_36746_24918# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2051 a_46390_58178# a_10515_22671# a_46882_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20510 a_1823_67668# a_1915_67477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X20511 VSS a_34411_50613# a_33360_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X20512 a_40366_16886# a_12899_11471# a_40858_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20513 a_19697_29423# a_19442_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20514 a_25702_69222# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20515 VSS a_7407_46529# a_7368_46403# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20516 VDD a_13357_32143# a_22230_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20517 VDD a_13445_51335# a_12755_51562# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X20518 VSS a_32920_34191# a_33026_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20519 vcm_commonmode a_16362_13508# a_44474_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2052 a_22690_57174# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20520 VSS a_3805_30083# a_4248_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20521 a_7545_32259# a_6883_37019# a_7473_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20522 vcm_commonmode a_16362_23548# a_27406_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20523 VSS a_24800_41953# a_25263_41001# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20524 a_9645_60214# a_6559_59879# a_9431_60214# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20525 a_31422_21540# a_16746_21538# a_31330_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20526 a_26310_58178# a_16362_58178# a_26402_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20527 a_1757_16917# a_1591_16917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20528 a_46786_16886# a_12727_13353# a_46390_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20529 a_5333_59343# a_5411_59317# a_5179_59663# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2053 a_2121_54447# a_1643_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20530 a_29718_68218# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20531 a_6989_24233# a_7059_24135# a_6835_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20532 vcm_commonmode a_16362_15516# a_17366_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20533 a_26310_17890# a_12899_10927# a_26802_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20534 VDD a_12947_71576# a_34342_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20535 a_5497_71855# a_5453_72097# a_5331_71855# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20536 a_21382_13508# a_16746_13506# a_21290_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20537 a_30818_15484# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20538 a_17763_35797# a_14293_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20539 a_33641_29967# a_33363_30305# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X2054 VDD a_12907_27023# a_43445_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X20540 a_13620_36519# a_13835_36649# a_13762_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20541 a_2319_57948# a_2124_57979# a_2629_57711# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X20542 a_11155_30663# a_10761_29745# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20543 a_34434_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20544 vcm_commonmode a_16362_8488# a_30418_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20545 a_4443_36611# a_4242_35407# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20546 a_19217_51701# a_4758_45369# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20547 a_46482_63198# a_16746_63200# a_46390_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20548 vcm_commonmode a_16362_60186# a_43470_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20549 a_17366_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2055 vcm_commonmode VSS a_28410_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20550 vcm_commonmode a_16362_19532# a_43470_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20551 a_47886_59504# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20552 a_19678_18894# a_12899_10927# a_19282_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20553 VSS a_10515_22671# a_23694_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20554 VSS a_5336_54965# a_5274_54991# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20555 a_20682_55166# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20556 a_33430_66210# a_16746_66212# a_33338_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20557 vcm_commonmode a_16362_70226# a_26402_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20558 VSS a_7377_18012# a_12323_20904# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X20559 a_7021_70339# a_5877_70197# a_6926_70339# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2056 VSS a_12877_14441# a_49798_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20560 VSS a_32181_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X20561 VDD a_12901_66665# a_38358_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20562 a_31330_11866# a_10055_58791# a_31822_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20563 a_17274_19898# a_11067_67279# a_17766_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20564 a_18627_42943# a_17711_43439# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X20565 a_21290_68218# a_12727_67753# a_21782_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20566 VDD a_12473_42869# a_12417_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20567 a_38450_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20568 VDD a_16257_38517# a_16287_38870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20569 a_3217_34319# a_3187_34293# a_3145_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2057 a_46786_11866# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20570 a_20378_60186# a_16746_60188# a_20286_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20571 a_25199_51183# a_24849_51183# a_25104_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20572 VDD a_12727_58255# a_24302_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20573 a_20378_19532# a_16746_19530# a_20286_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20574 VDD a_37527_29397# a_37747_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20575 VDD a_2840_66103# a_10147_65984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20576 VDD config_1_in[9] a_1591_7119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X20577 a_13431_27247# a_11430_26159# a_13241_27497# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X20578 a_42374_57174# a_12257_56623# a_42866_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20579 a_17777_49007# a_16587_49007# a_17668_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2058 a_2672_39049# a_1591_38677# a_2325_38645# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X20580 a_25306_67214# a_12983_63151# a_25798_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20581 a_36746_65206# a_10975_66407# a_36350_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20582 VDD a_2325_71285# a_2215_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20583 VSS a_9613_48981# a_9547_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20584 VDD a_23993_37981# a_23599_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20585 a_38606_28585# a_36904_28879# a_38524_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20586 a_49798_64202# a_12355_65103# a_49402_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20587 a_33712_51183# a_4482_57863# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X20588 a_42770_12870# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20589 a_30845_52047# a_28881_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2059 VSS a_14735_35805# a_14675_35831# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X20590 a_3985_22901# a_3325_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20591 a_2939_52245# a_1923_54591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20592 VSS a_2292_17179# a_2860_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.66e+10p ps=1.3e+06u w=420000u l=150000u
X20593 a_25702_22910# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20594 a_2672_39049# a_1757_38677# a_2325_38645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20595 VDD a_26417_47919# a_29956_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20596 VDD a_1586_21959# a_1591_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X20597 a_7376_60137# a_6559_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20598 a_9747_49929# a_9301_49557# a_9651_49929# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X20599 a_39758_56170# a_12257_56623# a_39362_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 a_15660_49257# a_10515_63143# a_15566_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X2060 a_32426_70226# a_16746_70228# a_32334_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20600 a_32826_56492# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20601 vcm_commonmode a_16362_67214# a_46482_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20602 VSS a_13576_37149# a_12677_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X20603 VSS a_12899_10927# a_18674_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20604 a_22690_15882# a_12877_14441# a_22294_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20605 a_17766_9460# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20606 a_29718_21906# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20607 vcm_commonmode a_16362_59182# a_36442_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20608 VSS a_12355_15055# a_44778_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20609 a_40458_57174# a_16746_57176# a_40366_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2061 a_12066_57167# a_11710_58487# a_11763_57399# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X20610 a_41766_18894# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20611 VSS VDD a_27710_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20612 a_31726_70226# a_12901_66665# a_31330_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20613 a_23790_58500# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20614 a_30091_35253# a_13097_36367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20615 a_19678_13874# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20616 a_2107_36873# a_1591_36501# a_2012_36861# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X20617 VSS a_10055_58791# a_23694_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20618 VSS a_10515_63143# a_12539_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20619 a_28115_43447# a_27183_43493# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2062 vcm_commonmode a_16362_11500# a_24394_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X20620 VDD VSS a_45386_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20621 vcm_commonmode a_16362_17524# a_32426_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20622 a_6971_19453# a_4792_20443# a_6608_19319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20623 a_4057_50645# a_3891_50645# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20624 a_24959_30503# a_34895_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20625 a_21686_62194# a_12981_62313# a_21290_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20626 a_7457_62927# a_2840_53511# a_7373_62927# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X20627 a_2781_30345# a_1591_29973# a_2672_30345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X20628 a_5136_34551# a_2473_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20629 a_7837_26703# a_3301_26703# a_7755_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2063 VSS a_33515_30511# a_33694_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X20630 VDD a_4343_60405# a_4274_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20631 a_33830_21508# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20632 a_33430_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20633 a_9560_58575# a_9424_60949# a_9370_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20634 a_16746_17522# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X20635 a_46390_71230# a_12901_66665# a_46882_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20636 a_36280_50639# a_35568_49525# a_35683_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20637 a_46882_20504# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20638 a_46482_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20639 VSS a_12985_19087# a_39758_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2064 a_10288_17143# a_5671_21495# a_10430_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X20640 a_18674_60186# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20641 a_17366_58178# a_16746_58180# a_17274_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20642 a_18674_19898# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20643 a_49402_64202# a_16362_64202# a_49494_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20644 VDD a_12981_62313# a_49402_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20645 a_20286_70226# a_16362_70226# a_20378_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20646 a_26345_40871# a_24561_41583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20647 a_7009_56623# a_1823_66941# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20648 a_15037_35077# a_15345_34717# a_15011_34717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X20649 a_49798_8854# a_12947_8725# a_49402_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2065 a_33338_13874# a_12727_15529# a_33830_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X20650 VSS a_2292_17179# a_6417_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20651 a_36842_12472# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20652 VDD a_12659_54965# a_12605_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20653 a_34342_13874# a_16362_13508# a_34434_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20654 VDD a_12546_22351# a_40366_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20655 a_19774_22512# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20656 a_37471_27497# a_20635_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20657 a_3063_34319# a_3187_34293# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20658 VDD a_11067_67279# a_23298_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20659 a_47394_12870# a_16362_12504# a_47486_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2066 a_34434_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20660 a_26402_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20661 a_23298_61190# a_16362_61190# a_23390_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20662 VSS a_12901_66959# a_47790_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20663 a_36442_24552# VDD a_36350_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20664 VDD a_17222_27247# a_18977_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20665 a_30835_39783# a_12725_44527# a_31009_39659# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20666 vcm_commonmode a_16362_66210# a_22386_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20667 a_35349_50095# a_35224_49871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20668 vcm_commonmode a_16362_20536# a_46482_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20669 a_49494_23548# a_16746_23546# a_49402_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2067 a_21479_40229# a_20713_40193# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X20670 VDD a_6515_62037# a_8497_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20671 a_24302_24918# VSS a_24394_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20672 VSS a_14646_29423# a_23303_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20673 a_27806_70548# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20674 a_41766_59182# a_12727_58255# a_41370_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20675 VDD a_12947_8725# a_42374_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20676 a_36350_7850# VDD a_36842_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20677 a_35838_18496# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20678 a_24394_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20679 a_21719_48285# a_21095_47919# a_21611_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2068 a_8740_64783# a_7803_55509# a_8638_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=150000u
X20680 VSS a_10286_26311# a_10244_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20681 VSS a_28963_28853# a_29545_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20682 a_39459_44527# a_39282_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20683 a_24698_69222# a_12516_7093# a_24302_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20684 a_33668_38567# a_32795_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20685 a_27314_60186# a_16362_60186# a_27406_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20686 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X20687 a_48794_65206# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20688 a_5791_43541# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20689 a_39454_15516# a_16746_15514# a_39362_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2069 a_23790_19500# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20690 vcm_commonmode a_16362_12504# a_36442_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20691 VSS a_1586_36727# a_2971_37589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20692 a_40458_10496# a_16746_10494# a_40366_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20693 a_46390_18894# a_16362_18528# a_46482_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20694 a_35647_38053# a_32031_37683# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X20695 VDD a_12985_16367# a_17274_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20696 a_19913_49917# a_19878_49683# a_19675_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20697 a_7815_49855# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20698 a_9775_64783# a_9280_65327# a_9557_64757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20699 a_3714_56118# a_3668_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X207 a_25798_57496# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2070 a_22386_62194# a_16746_62196# a_22294_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20700 a_26239_31849# a_13357_32143# a_26157_31605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20701 VDD a_6521_58773# a_5612_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20702 a_38754_57174# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20703 a_18674_7850# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20704 a_40366_67214# a_16362_67214# a_40458_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20705 a_45782_58178# a_12901_58799# a_45386_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20706 VSS VSS a_42770_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20707 VDD a_23628_35823# a_23734_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20708 VDD a_1923_59583# a_1643_59317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20709 a_5531_22895# a_5087_23145# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X2071 a_17798_32143# a_17711_32385# a_17394_32275# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20710 a_13925_51727# a_13735_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20711 a_2886_65910# a_2840_66103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20712 a_32167_29611# a_4811_34855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20713 a_5885_39759# a_4314_40821# a_5813_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20714 VSS a_21233_40956# a_20925_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20715 a_28714_68218# a_12901_66959# a_28318_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20716 VSS a_12355_65103# a_25702_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20717 a_48890_61512# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20718 a_36275_47695# a_22291_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20719 vcm_commonmode a_16362_56170# a_29414_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2072 a_13097_39631# a_12831_39997# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20720 a_39854_19500# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20721 VSS a_32795_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X20722 a_40366_8854# a_16362_8488# a_40458_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20723 VSS a_17709_48761# a_17643_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20724 a_6892_40303# a_6559_39759# a_6671_40630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20725 VDD a_12355_15055# a_25306_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20726 VSS a_2467_67668# a_2263_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X20727 a_30418_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20728 a_17366_11500# a_16746_11498# a_17274_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20729 VDD a_12727_13353# a_29322_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2073 a_47394_8854# a_12985_19087# a_47886_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20730 a_8021_27497# a_3301_26703# a_7939_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20731 a_33515_48576# a_32856_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20732 VDD a_4482_57863# a_30561_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20733 VDD a_10873_27497# a_20027_27221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X20734 a_12404_34191# a_12227_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20735 a_34342_58178# a_16362_58178# a_34434_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20736 a_47886_67536# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20737 VDD a_14471_28585# a_16101_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X20738 a_14095_30083# a_6459_30511# a_14013_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20739 a_20682_63198# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2074 a_12793_44310# a_12621_44099# a_12579_44310# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X20740 a_26402_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20741 a_17274_68218# a_16362_68218# a_17366_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20742 a_21782_7452# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20743 VDD a_2840_53511# a_7079_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20744 VDD a_3143_66972# a_7155_55509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X20745 a_47394_57174# a_16362_57174# a_47486_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20746 a_33734_62194# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20747 a_34342_17890# a_12899_10927# a_34834_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20748 VSS a_12947_23413# a_34738_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20749 a_4055_30083# a_3325_29967# a_3983_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2075 a_26706_14878# a_12727_15529# a_26310_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20750 a_7183_42845# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20751 VDD VDD a_31330_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20752 a_8205_26159# a_4528_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20753 VDD a_10515_22671# a_41370_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20754 VSS a_10515_23975# a_47790_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20755 VSS a_6515_67477# a_7197_66237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X20756 a_12024_30199# a_11710_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20757 a_32187_36161# a_30757_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20758 VDD a_12727_67753# a_24302_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20759 VSS a_43495_28487# a_43445_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2076 VDD a_11764_65845# a_9624_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X20760 a_10045_29967# a_3339_32463# a_9963_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20761 VDD a_2606_41079# a_18653_48502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20762 VDD a_1761_35407# a_32143_35281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X20763 vcm_commonmode a_16362_70226# a_34434_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20764 a_6793_47713# a_6727_47607# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20765 a_24394_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20766 a_4866_13647# a_4812_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20767 a_5962_72221# a_4885_71855# a_5800_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20768 a_11947_68279# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20769 a_6641_67279# a_6224_73095# a_6156_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2077 a_9775_64783# a_9735_63669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X20770 a_2467_67668# a_2559_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20771 a_41766_12870# a_10055_58791# a_41370_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20772 a_2215_45199# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20773 a_9290_57167# a_8491_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20774 a_24698_64202# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20775 a_38358_55166# VSS a_38850_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20776 a_10713_14191# a_10678_14443# a_10475_14165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20777 a_24698_22910# a_11067_21583# a_24302_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20778 a_22294_21906# a_11067_21583# a_22786_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20779 a_22294_17890# a_16362_17524# a_22386_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2078 a_28108_48463# a_27509_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20780 VSS a_3295_54421# a_10791_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20781 VDD a_12727_58255# a_32334_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20782 a_9643_13430# a_7841_12167# a_9184_13255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20783 vcm_commonmode a_16362_61190# a_37446_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20784 a_49798_72234# VDD a_49402_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20785 VDD a_9367_29397# a_9325_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20786 VDD a_12901_58799# a_45386_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20787 a_41462_18528# a_16746_18526# a_41370_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20788 a_39000_47081# a_8491_41383# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20789 a_38754_10862# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2079 a_2981_27023# a_2315_24540# a_2899_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20790 a_45782_11866# a_12985_16367# a_45386_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20791 a_28810_15484# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20792 a_25306_12870# a_12877_16911# a_25798_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20793 a_28714_21906# a_12985_7663# a_28318_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20794 VSS a_23467_41237# a_23415_41263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20795 VDD a_4339_64521# a_9645_60214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20796 a_3707_25731# a_2315_24540# a_3611_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X20797 a_18358_31599# a_18328_31573# a_18063_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20798 a_8958_65961# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20799 vcm_commonmode a_16362_14512# a_42466_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X208 a_15221_39631# a_14951_39997# a_15131_39997# VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2080 VDD a_2928_22583# a_2007_20149# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20800 VSS a_24800_35425# a_25263_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X20801 a_18674_13874# a_12877_16911# a_18278_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20802 a_21611_47919# a_21095_47919# a_21516_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20803 vcm_commonmode VSS a_25398_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20804 VSS a_12703_38517# a_12341_41281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20805 VSS a_22015_28111# a_33597_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20806 a_38358_72234# VSS a_38450_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20807 a_29322_11866# a_10055_58791# a_29814_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20808 a_42466_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20809 a_19282_68218# a_12727_67753# a_19774_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2081 a_5993_37039# a_5455_37039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20810 a_16158_30511# a_14361_29967# a_15207_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20811 VSS a_36890_34191# a_37711_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20812 a_23790_66532# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20813 a_20286_63198# a_12981_62313# a_20778_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20814 a_18370_60186# a_16746_60188# a_18278_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20815 a_18370_19532# a_16746_19530# a_18278_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20816 a_37374_51183# a_37307_51339# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20817 VSS a_12901_58799# a_30722_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20818 VSS a_7755_26703# a_8516_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20819 VDD a_36324_34191# a_36430_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2082 a_2882_54813# a_2163_54589# a_2319_54684# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X20820 VDD a_20027_27221# a_19889_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X20821 a_10870_31599# a_9307_30663# a_10701_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20822 vcm_commonmode a_16362_15516# a_28410_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20823 a_32426_13508# a_16746_13506# a_32334_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20824 a_29956_48169# a_26514_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20825 a_9031_54135# a_2840_53511# a_9376_54223# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X20826 a_28902_28335# a_23928_28585# a_28816_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20827 VDD a_21737_49249# a_21627_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20828 a_1761_25615# a_1591_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X20829 a_45478_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2083 VSS a_9669_26703# a_11251_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20830 a_3813_39759# a_3759_39991# a_2927_39733# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20831 VDD a_1952_60431# a_1899_53387# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20832 a_24302_62194# a_12355_15055# a_24794_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20833 a_8215_25071# a_6162_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20834 a_12981_59343# a_12712_59343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X20835 a_10901_52245# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X20836 a_10109_73487# a_9707_73807# a_9945_73807# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X20837 VSS a_12901_66665# a_48794_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20838 a_31726_55166# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20839 a_44474_66210# a_16746_66212# a_44382_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2084 a_27314_69222# a_12901_66959# a_27806_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20840 VSS a_30052_32117# a_30743_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20841 VDD a_12473_36341# a_12417_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X20842 a_46482_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20843 VDD a_24194_35823# a_24703_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20844 a_43378_21906# a_16362_21540# a_43470_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20845 a_18811_38053# a_18045_38017# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X20846 VDD a_12901_66665# a_49402_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20847 a_14859_43447# a_15253_43421# a_14919_43421# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X20848 a_8935_27791# a_8662_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X20849 a_11829_63151# a_11145_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2085 a_38754_67214# a_12727_67753# a_38358_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20850 a_28318_19898# a_11067_67279# a_28810_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20851 a_9637_30511# a_9161_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X20852 a_49494_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20853 a_42770_61190# a_12355_15055# a_42374_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20854 a_1887_10422# a_1929_10651# a_1887_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20855 VDD a_5903_13967# a_6362_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X20856 a_37527_29397# a_38378_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20857 VDD a_2847_51157# a_2834_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20858 a_25702_71230# a_12947_71576# a_25306_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20859 VDD a_4035_11989# a_3983_12015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2086 a_27891_41495# a_12725_44527# a_28065_41601# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20860 VSS a_9613_13077# a_9547_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20861 a_48490_65206# a_16746_65208# a_48398_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20862 a_40457_27765# a_40086_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20863 a_20378_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20864 a_35438_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20865 VDD a_4555_55233# a_4516_55107# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X20866 VDD a_7037_19385# a_7067_19126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20867 a_47394_20902# a_16362_20536# a_47486_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20868 a_4043_44343# a_3987_19623# a_4217_44449# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20869 a_4607_48463# a_3983_48469# a_4499_48841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2087 VDD a_10680_52245# a_8491_57487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X20870 a_12985_16367# a_12815_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X20871 a_2058_33775# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20872 a_38450_57174# a_16746_57176# a_38358_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20873 a_39758_18894# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20874 a_2596_16911# a_1757_16917# a_2620_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20875 VSS a_12899_11471# a_43774_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20876 a_40762_13874# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20877 vcm_commonmode a_16362_64202# a_18370_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20878 a_41462_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20879 VSS a_9484_11989# a_10341_10703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2088 VSS a_11067_13095# a_35742_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X20880 a_23694_23914# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20881 a_40743_31287# a_32970_31145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X20882 a_30722_24918# VSS a_30326_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20883 a_24394_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20884 a_33338_9858# a_16362_9492# a_33430_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20885 a_35438_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20886 a_2693_68021# a_2475_68425# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X20887 a_3383_54269# a_2913_54991# a_3020_54135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20888 a_30818_57496# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20889 a_44382_59182# a_12901_58799# a_44874_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2089 a_31822_67536# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20890 VSS a_2775_46025# a_30530_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20891 a_20682_16886# a_12727_13353# a_20286_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20892 VSS a_12899_10927# a_29718_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20893 a_26341_47491# a_25015_48437# a_26259_47491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20894 VSS a_12877_16911# a_30722_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20895 VSS a_12981_62313# a_42770_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20896 a_39454_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20897 a_1644_58229# a_1591_56623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20898 VSS a_43495_28487# a_43531_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20899 VSS a_2686_70223# a_5021_70561# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X209 a_33689_29423# a_30788_28487# a_33008_28853# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2090 a_29718_8854# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20900 a_32730_69222# a_12516_7093# a_32334_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20901 VDD config_1_in[8] a_1591_6031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X20902 a_9669_26703# a_9289_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20903 VDD a_15271_41781# a_15095_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20904 a_2012_9839# a_1867_10927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20905 a_16648_40517# a_15775_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20906 a_3583_73865# a_3137_73493# a_3487_73865# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20907 a_21782_59504# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20908 a_11455_12157# a_1586_18695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20909 a_17670_14878# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2091 a_2743_31094# a_1915_35015# a_2284_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X20910 a_7197_66237# a_6927_65871# a_7107_65871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20911 a_49402_8854# a_16362_8488# a_49494_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20912 a_36350_24918# VSS a_36842_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20913 a_19424_39631# a_15189_39889# a_19203_39958# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20914 a_44382_7850# VDD a_44874_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20915 a_40858_22512# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20916 vcm_commonmode a_16362_18528# a_30418_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20917 a_9223_23145# a_5531_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20918 a_2663_43541# a_2872_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X20919 VDD a_7571_26151# a_12236_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2092 a_9731_22895# a_9223_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.35e+11p pd=2.67e+06u as=0p ps=0u w=1e+06u l=150000u
X20920 VSS a_3024_67191# a_8994_63927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20921 a_25305_37782# a_25133_37571# a_25091_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X20922 a_38754_7850# VDD a_38358_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20923 VSS a_12473_36341# a_12417_36694# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20924 a_8509_47673# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X20925 VSS a_12355_65103# a_33734_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20926 a_36432_42919# a_35463_42943# a_36336_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20927 VDD a_12899_11471# a_33338_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20928 VSS a_13484_39325# a_12585_39069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X20929 a_16746_70228# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X2093 VSS a_10883_18007# a_1586_18695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X20930 a_12202_54019# a_6095_44807# a_12120_54019# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X20931 VSS a_11067_13095# a_46786_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20932 a_18611_52047# a_28817_29111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20933 a_5600_10927# a_5483_11140# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20934 a_44874_21508# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20935 a_28108_48463# a_27929_48579# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20936 a_44474_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20937 a_41370_14878# a_16362_14512# a_41462_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20938 VSS a_12546_22351# a_19678_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20939 a_7159_50260# a_7251_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2094 VDD a_9361_28335# a_9529_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=6
X20940 a_7871_59049# a_7107_58487# a_8065_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20941 a_35458_28879# a_32823_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20942 a_47394_65206# a_16362_65206# a_47486_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20943 a_13239_29575# a_12965_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X20944 VDD a_19626_31751# a_32626_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20945 VSS a_12947_56817# a_36746_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20946 a_14008_51727# a_12683_51329# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20947 a_29718_9858# a_12985_19087# a_29322_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20948 a_31330_70226# a_16362_70226# a_31422_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20949 VDD a_12727_13353# a_37354_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2095 a_36350_65206# a_16362_65206# a_36442_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20950 a_34834_13476# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20951 a_11163_25321# a_9955_20969# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20952 VSS a_10975_66407# a_19678_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20953 a_23694_64202# a_12355_65103# a_23298_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20954 a_17766_23516# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20955 a_39836_38567# a_38867_38591# a_39740_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X20956 a_17366_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20957 a_7229_30511# a_5441_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20958 a_38450_10496# a_16746_10494# a_38358_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20959 a_2672_49929# a_1757_49557# a_2325_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2096 a_10873_15529# a_10673_15055# a_10791_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20960 a_12710_63151# a_10515_63143# a_12624_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20961 a_47886_12472# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20962 VDD a_12985_7663# a_21290_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20963 a_45386_13874# a_16362_13508# a_45478_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20964 a_22181_50645# a_22015_50645# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20965 a_1915_24148# a_2007_23957# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20966 VDD a_14831_50095# a_32494_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20967 a_24394_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20968 a_21290_62194# a_16362_62194# a_21382_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20969 a_24698_72234# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2097 VDD a_3339_43023# a_8583_33551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u M=6
X20970 VSS a_2473_40821# a_1895_40516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X20971 vcm_commonmode a_16362_67214# a_20378_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20972 a_4797_62063# a_4441_62327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20973 a_2012_44655# a_1778_42631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20974 a_20592_46983# a_7571_29199# a_20734_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20975 a_47486_24552# VDD a_47394_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20976 VDD a_12727_67753# a_32334_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20977 a_18278_15882# a_16362_15516# a_18370_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20978 vcm_commonmode a_16362_66210# a_33430_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20979 VDD a_10055_58791# a_24302_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2098 VDD a_10515_23975# a_49402_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X20980 a_2824_70197# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20981 a_22386_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20982 a_3572_56311# a_3005_56079# a_3714_56118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20983 a_31022_31375# a_29926_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20984 VDD a_12983_63151# a_45386_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X20985 a_42866_63520# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20986 vcm_commonmode a_16362_9492# a_35438_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20987 a_37446_16520# a_16746_16518# a_37354_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X20988 VSS a_2292_43291# a_2369_45565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20989 a_17670_55166# VSS a_17274_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2099 a_40458_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X20990 a_2744_66103# a_1768_16367# a_2886_65910# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X20991 VSS a_21663_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X20992 VSS a_35647_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X20993 a_10753_12559# a_10317_13647# a_10681_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20994 a_32730_22910# a_11067_21583# a_32334_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20995 VSS a_10391_49855# a_10325_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20996 VSS a_12981_59343# a_31726_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20997 a_10912_14557# a_10475_14165# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20998 VDD a_33694_30761# a_41046_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X20999 a_28410_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u M=564
X210 a_11433_69921# a_11215_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X2100 VDD a_43003_30761# a_23395_32463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21000 VDD a_2689_65103# a_6457_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21001 a_45478_9492# a_16746_9490# a_45386_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21002 a_36746_58178# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21003 VSS a_9963_29967# a_10506_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21004 VDD a_12985_16367# a_28318_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21005 VDD a_12901_66959# a_18278_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21006 a_13527_27247# a_12349_25847# a_13431_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21007 a_16615_41001# a_12713_41923# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21008 a_7821_20291# a_4792_20443# a_7749_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21009 a_16615_39095# a_15683_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2101 VSS a_40737_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21010 a_46882_62516# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21011 a_36579_40183# a_35647_40229# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21012 a_7159_22583# a_7431_22441# a_7389_22467# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21013 vcm_commonmode a_16362_57174# a_27406_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21014 VDD a_2317_28892# a_5337_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21015 VSS a_18197_36604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21016 a_31422_55166# VDD a_31330_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21017 a_32730_16886# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21018 a_10299_47607# a_10407_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21019 a_30326_10862# a_16362_10496# a_30418_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2102 a_13867_39631# a_13613_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21020 a_13888_43781# a_13015_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21021 a_20286_71230# a_12901_66665# a_20778_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21022 a_41370_59182# a_16362_59182# a_41462_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21023 a_19774_64524# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21024 a_30835_38695# a_26433_39631# a_31009_38571# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X21025 a_12663_35431# a_32187_36161# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X21026 VDD a_12981_62313# a_23298_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21027 a_9123_57399# a_9135_56623# a_9468_57487# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X21028 a_39188_39429# a_38315_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21029 a_44778_69222# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2103 VSS a_10515_23975# a_31726_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21030 a_77664_40024# clk_vcm a_77922_40050# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21031 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X21032 a_7183_49551# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21033 VSS a_6099_23983# a_5085_23047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21034 a_24561_41583# a_24382_41629# a_24573_41263# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21035 a_12161_62973# a_11943_63125# a_12055_62973# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.596e+11p ps=1.6e+06u w=420000u l=150000u
X21036 a_34395_31287# a_32970_31145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21037 a_24302_70226# a_12516_7093# a_24794_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21038 a_45386_58178# a_16362_58178# a_45478_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21039 a_31726_63198# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2104 a_40762_70226# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21040 vcm_commonmode a_16362_71230# a_41462_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21041 VSS a_9187_56597# a_9135_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21042 VDD a_32971_35281# a_32831_35307# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21043 a_28318_68218# a_16362_68218# a_28410_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21044 a_9490_11177# a_9455_11079# a_9187_10901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21045 VSS a_12901_66959# a_21686_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21046 a_12713_53181# a_12202_54599# a_12631_52928# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21047 a_45386_17890# a_12899_10927# a_45878_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21048 VSS a_12947_23413# a_45782_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21049 a_30908_40743# a_30035_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2105 a_28410_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21050 vcm_commonmode a_16362_20536# a_20378_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21051 a_23390_23548# a_16746_23546# a_23298_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21052 VDD a_32370_50871# a_32091_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X21053 a_22386_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21054 VSS a_38076_31573# a_30788_28487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21055 a_36442_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21056 a_38754_18894# a_12899_10927# a_38358_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21057 VSS a_12727_13353# a_35742_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21058 VSS a_41842_27221# a_41783_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21059 a_1941_47381# a_1775_47381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2106 VDD a_20715_34717# a_20741_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X21060 vcm_commonmode a_16362_70226# a_45478_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21061 VSS a_32795_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21062 a_14634_47349# a_5039_42167# a_15017_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X21063 a_22690_65206# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21064 a_29708_27907# a_16863_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21065 a_37799_43777# a_12357_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21066 a_22786_17492# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21067 a_49402_16886# a_12899_11471# a_49894_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21068 a_20286_18894# a_16362_18528# a_20378_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21069 a_11763_62581# a_11521_66567# a_12161_62973# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2107 VDD a_9963_50959# a_12993_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X21070 VSS a_3247_20495# a_5353_43343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21071 a_40366_68218# a_12727_67753# a_40858_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21072 a_39431_37737# a_38499_37503# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21073 vcm_commonmode a_16362_62194# a_35438_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21074 a_33338_21906# a_11067_21583# a_33830_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21075 a_36350_58178# a_10515_22671# a_36842_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21076 a_12713_20495# a_4792_20443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21077 a_33338_17890# a_16362_17524# a_33430_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21078 a_4607_65693# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21079 a_12289_54475# a_12202_54599# a_12203_54475# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2108 a_4340_58799# a_4298_58951# a_4037_58773# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X21080 a_5869_15055# a_5755_14709# a_5052_14709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21081 VSS a_75199_38962# a_75628_38962# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21082 VDD a_12727_58255# a_43378_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21083 VSS a_1761_47919# a_28099_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21084 vcm_commonmode VSS a_18370_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21085 VSS a_12877_14441# a_39758_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21086 a_36746_11866# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21087 VDD a_2847_23743# a_2834_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21088 vcm_commonmode a_16362_61190# a_48490_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21089 a_3254_19126# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2109 VDD a_12877_14441# a_39362_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21090 a_5781_44449# a_5715_44343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21091 a_22386_70226# a_16746_70228# a_22294_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21092 VSS a_12901_58799# a_28714_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21093 a_25702_56170# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21094 a_1757_18543# a_1591_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21095 VSS a_4571_26677# a_7939_27497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21096 a_26802_16488# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21097 a_23298_13874# a_12727_15529# a_23790_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21098 a_5757_56623# a_5378_56989# a_5685_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21099 a_44382_67214# a_12983_63151# a_44874_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X211 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u M=394
X2110 vcm_commonmode a_16362_69222# a_48490_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21100 a_18627_44581# a_16928_44007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X21101 vcm_commonmode a_16362_10496# a_27406_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21102 a_23195_29967# a_22922_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21103 a_14830_48463# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21104 a_43470_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21105 a_15775_40229# a_15009_40193# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X21106 a_25398_61190# a_16746_61192# a_25306_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21107 a_7653_22057# a_5085_23047# a_7571_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21108 a_2319_57948# a_2163_57853# a_2464_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21109 a_29718_55166# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2111 a_27688_42693# a_27245_41829# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X21110 a_29718_13874# a_12877_16911# a_29322_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21111 a_7467_61751# a_7676_61493# a_7634_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21112 a_38077_29941# a_38210_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21113 a_44778_22910# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21114 VDD a_4685_37583# a_6807_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21115 a_17274_69222# a_12901_66959# a_17766_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21116 a_21782_67536# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21117 VSS a_49876_41198# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.84e+07u l=3.9e+06u
X21118 a_7942_31849# a_5993_32687# a_7828_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21119 a_31330_63198# a_12981_62313# a_31822_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2112 VDD a_10935_11989# a_9491_12297# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21120 a_29414_60186# a_16746_60188# a_29322_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21121 a_16746_68220# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X21122 vcm_commonmode a_16362_16520# a_26402_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21123 a_29414_19532# a_16746_19530# a_29322_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21124 VDD a_10515_23975# a_39362_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21125 a_11780_69679# a_10865_69679# a_11433_69921# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21126 a_30418_14512# a_16746_14510# a_30326_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21127 VSS a_10515_23975# a_21686_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21128 VDD a_1925_22583# a_1738_22325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21129 a_18370_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2113 a_2629_57711# a_2250_58077# a_2557_57711# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X21130 a_11793_12559# a_10753_12559# a_11711_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21131 a_2464_64605# a_2250_64605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21132 VDD a_7571_29199# a_12513_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21133 VSS a_1803_20719# a_32327_40191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21134 vcm_commonmode a_16362_69222# a_38450_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21135 VSS VDD a_46786_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21136 a_42466_67214# a_16746_67216# a_42374_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21137 a_8102_11587# a_7203_10383# a_8029_11587# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21138 VDD a_7695_31573# a_12875_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21139 a_11617_72097# a_11399_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2114 VSS a_3972_25615# a_6835_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21140 a_4866_13967# a_4057_13647# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21141 a_41370_22910# a_16362_22544# a_41462_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21142 a_13983_36367# a_13835_36649# a_13620_36519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21143 a_3421_57167# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21144 VDD a_3339_43023# a_12227_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21145 a_23734_29941# a_15548_30761# a_24042_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21146 a_40762_62194# a_12981_62313# a_40366_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21147 a_3137_73493# a_2971_73493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21148 VDD a_20351_49525# a_20282_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21149 a_28810_57496# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2115 VDD a_3295_62083# a_3108_62043# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X21150 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X21151 a_23694_72234# VDD a_23298_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21152 VDD a_30788_28487# a_22843_29415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X21153 a_7757_21379# a_2339_38129# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21154 VSS a_13848_44135# a_13661_43957# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21155 a_33591_32375# a_29927_29199# a_33825_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21156 a_12445_50613# a_12227_51017# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21157 a_30625_52245# a_28881_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21158 a_7473_24527# a_4571_26677# a_7367_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
X21159 a_5269_43809# a_5051_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2116 a_40762_8854# a_12947_8725# a_40366_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21160 a_7959_15279# a_7987_15431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21161 a_2244_22583# config_1_in[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21162 VSS a_12877_16911# a_28714_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21163 VDD a_6177_61127# a_5653_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X21164 a_37750_60186# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21165 a_36442_58178# a_16746_58180# a_36350_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21166 a_37750_19898# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21167 a_34909_44869# a_35217_44509# a_24800_43041# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21168 a_27791_52637# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21169 a_19374_68218# a_16746_68220# a_19282_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2117 VDD a_1923_54591# a_4311_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21170 a_10791_27247# a_7369_24233# a_10873_27497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21171 a_49494_57174# a_16746_57176# a_49402_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21172 a_21686_24918# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21173 a_77568_40202# a_77664_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21174 a_18278_23914# a_16362_23548# a_18370_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21175 a_28757_30539# a_28670_30663# a_28671_30539# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X21176 a_12757_8207# a_12479_8545# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21177 a_11507_18909# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21178 a_38850_22512# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21179 a_4404_45743# a_4259_45199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2118 VDD a_14679_31288# a_5915_30287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X21180 a_16953_51425# a_16735_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21181 a_42866_71552# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21182 VDD a_11067_67279# a_42374_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21183 a_5340_32687# a_4425_32687# a_4993_32929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21184 VSS a_13620_36519# a_12889_35537# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21185 a_17670_63198# a_15439_49525# a_17274_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21186 a_42374_61190# a_16362_61190# a_42466_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21187 a_25306_71230# a_16362_71230# a_25398_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21188 a_48490_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21189 VSS a_12895_13967# a_27710_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2119 a_22294_55166# VSS a_22786_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21190 VDD a_10055_58791# a_32334_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21191 a_31726_16886# a_12727_13353# a_31330_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21192 a_8165_48829# a_8121_48437# a_7999_48841# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X21193 VDD a_12947_8725# a_36350_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21194 VSS a_8969_42233# a_8903_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21195 a_46882_70548# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21196 a_39362_14878# a_16362_14512# a_39454_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21197 VDD a_24893_37429# a_25305_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21198 a_43470_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21199 a_43774_69222# a_12516_7093# a_43378_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X212 a_34434_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2120 VDD a_17927_31573# a_17488_48731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21200 VSS a_10975_66407# a_40762_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21201 a_24302_8854# a_12985_19087# a_24794_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21202 a_2847_66389# a_2672_66415# a_3026_66415# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21203 a_31422_63198# a_16746_63200# a_31330_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21204 a_29322_70226# a_16362_70226# a_29414_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21205 a_32826_59504# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21206 a_31994_30511# a_31964_30485# a_31904_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21207 a_28714_14878# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21208 a_5064_20719# a_4149_20719# a_4717_20961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21209 a_3325_29967# a_2847_30271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2121 a_43774_61190# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21210 vcm_commonmode a_16362_22544# a_38450_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21211 a_12877_14441# a_11067_63143# a_12805_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21212 a_18674_8854# a_12947_8725# a_18278_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21213 a_42466_20536# a_16746_20534# a_42374_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21214 a_19774_72556# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21215 VSS a_14471_28585# a_16824_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21216 a_2691_40847# a_2606_41079# a_2473_40821# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21217 a_30722_8854# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21218 VDD a_10288_53047# a_9507_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21219 VDD a_12901_66665# a_23298_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2122 a_10506_30511# a_9405_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X21220 VDD a_12981_59343# a_19282_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21221 a_19282_62194# a_16362_62194# a_19374_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21222 VDD a_11335_10076# a_11266_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21223 a_9353_72399# a_9075_72737# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21224 a_26445_38341# a_26753_37981# a_13909_38659# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21225 a_23390_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21226 a_47790_68218# a_12901_66959# a_47394_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21227 VSS a_12355_65103# a_44778_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21228 VDD a_12899_11471# a_44382_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21229 a_42466_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2123 a_42466_59182# a_16746_59184# a_42374_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21230 VDD a_35676_49525# a_37594_50755# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21231 a_42040_42919# a_41167_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21232 VDD a_9484_11989# a_9497_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21233 VDD a_5885_39759# a_6927_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21234 VSS a_12257_56623# a_34738_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21235 a_30657_29967# a_30565_30199# a_30440_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21236 a_7523_62581# a_9544_61635# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21237 a_27333_52271# a_27167_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21238 VSS a_12983_63151# a_17670_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21239 a_21686_65206# a_10975_66407# a_21290_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2124 a_26706_71230# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21240 VSS a_12947_56817# a_47790_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21241 a_5451_14735# a_5465_14967# a_5052_14709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21242 VSS a_23901_43132# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21243 VDD a_16953_51425# a_16843_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21244 a_36442_11500# a_16746_11498# a_36350_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21245 VDD a_12727_13353# a_48398_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21246 a_45878_13476# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21247 VSS a_21479_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21248 VDD a_12895_13967# a_35346_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21249 a_19374_21540# a_16746_21538# a_19282_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2125 VSS a_16510_8760# a_16746_10494# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X21250 a_11866_27791# a_7369_24233# a_12010_28111# VSS sky130_fd_pr__nfet_01v8 ad=3.9325e+11p pd=2.51e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X21251 a_4275_36201# a_4242_35407# a_4314_40821# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21252 a_38121_48169# a_37557_32463# a_21371_50959# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X21253 a_49494_10496# a_16746_10494# a_49402_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21254 VDD a_1586_21959# a_1591_23445# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X21255 a_8533_74941# a_8489_74549# a_8367_74953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21256 a_6097_16609# a_5879_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21257 a_34434_8488# a_16746_8486# a_34342_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21258 a_2952_46805# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21259 VDD a_15439_49525# a_17274_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2126 VDD a_3983_70767# a_4060_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21260 a_49402_67214# a_16362_67214# a_49494_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21261 a_24698_56170# a_12257_56623# a_24302_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21262 vcm_commonmode a_16362_67214# a_31422_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21263 a_39854_69544# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21264 a_23669_49007# a_17682_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21265 a_36350_66210# a_10975_66407# a_36842_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21266 VDD a_12727_67753# a_43378_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21267 a_40858_64524# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21268 a_38115_32463# a_38239_32375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21269 VDD a_19594_35823# a_23451_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2127 a_25398_69222# a_16746_69224# a_25306_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21270 a_39362_59182# a_16362_59182# a_39454_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21271 a_4941_35407# a_1915_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21272 vcm_commonmode a_16362_8488# a_32426_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21273 a_43470_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21274 vcm_commonmode a_16362_59182# a_21382_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21275 a_2347_28918# a_2317_28892# a_2275_28918# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X21276 a_5913_11169# a_5695_10927# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21277 a_1644_77813# a_1823_77821# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21278 a_26402_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21279 VSS a_24893_37429# a_25312_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2128 VDD a_32319_31599# a_19807_28111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X21280 a_28714_55166# VSS a_28318_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21281 VSS a_3417_31599# a_3983_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21282 a_43774_22910# a_11067_21583# a_43378_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21283 VDD a_8531_70543# a_33697_50359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21284 a_4497_29673# a_1915_35015# a_4425_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X21285 a_41370_60186# a_12727_58255# a_41862_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21286 a_10299_11703# a_10317_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21287 VDD VSS a_30326_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21288 a_27398_50461# a_26321_50095# a_27236_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21289 a_27791_52637# a_27167_52271# a_27683_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2129 VSS config_1_in[5] a_1591_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21290 VDD a_12901_66959# a_29322_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21291 VDD a_5254_67503# a_8332_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21292 a_29718_63198# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21293 vcm_commonmode a_16362_71230# a_39454_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21294 vcm_commonmode a_16362_58178# a_25398_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21295 VSS a_4427_25071# a_6007_23145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21296 a_17739_48502# a_17488_48731# a_17280_48695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21297 a_34834_55488# a_8295_47388# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21298 VDD a_13669_38517# a_14859_38909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21299 a_47790_21906# a_12985_7663# a_47394_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_39362_59182# a_12901_58799# a_39854_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2130 VDD a_12983_63151# a_34342_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21300 VDD a_6671_51183# a_7073_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21301 a_44382_12870# a_12877_16911# a_44874_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21302 a_17766_65528# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21303 a_27688_42693# a_26815_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21304 a_27314_22910# a_10515_23975# a_27806_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21305 a_31330_71230# a_12901_66665# a_31822_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21306 a_33430_61190# a_16746_61192# a_33338_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21307 a_17274_55166# VSS a_17366_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21308 a_31822_20504# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21309 a_31422_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2131 VDD a_9507_53877# a_9465_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21310 VDD a_10964_25615# a_14482_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21311 a_37750_13874# a_12877_16911# a_37354_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21312 a_1761_43567# a_1591_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21313 VSS a_12985_16367# a_34738_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21314 a_27183_44581# a_23567_44211# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X21315 vcm_commonmode VSS a_44474_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21316 a_24497_47349# a_24279_47753# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21317 a_17274_14878# a_12877_14441# a_17766_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21318 VSS a_12985_7663# a_17670_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21319 a_15974_51843# a_15261_51433# a_15892_51843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2132 a_22690_10862# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21320 a_21782_12472# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21321 VSS a_21663_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21322 VSS a_34699_42035# a_34639_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21323 VDD a_6098_73095# a_6099_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21324 vcm_commonmode a_16362_16520# a_34434_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21325 VSS a_7676_61493# a_8201_62839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21326 a_43378_18894# a_12895_13967# a_43870_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21327 a_3203_65910# a_2952_66139# a_2744_66103# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21328 a_32334_12870# a_16362_12504# a_32426_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21329 a_9301_67503# a_9135_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2133 a_5779_18038# a_3325_18543# a_5320_18231# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X21330 VDD a_5871_47594# a_4240_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X21331 a_2886_66237# a_2840_66103# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21332 VSS a_12901_66959# a_32730_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21333 vcm_commonmode a_16362_15516# a_47486_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21334 a_21382_24552# VDD a_21290_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21335 a_7472_32937# a_6243_30662# a_7390_32693# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21336 a_5695_74031# a_5179_74031# a_5600_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X21337 a_34434_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21338 a_36746_60186# a_12981_59343# a_36350_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21339 a_12093_21583# a_11887_19087# a_11990_21583# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X2134 VDD a_5490_41365# a_5098_41641# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X21340 a_36746_19898# a_12895_13967# a_36350_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21341 vcm_commonmode a_16362_20536# a_31422_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21342 a_15775_44581# a_13984_43781# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X21343 a_19678_70226# a_12901_66665# a_19282_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21344 a_19774_9460# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21345 a_47486_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21346 a_20778_18496# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21347 a_49798_18894# a_12899_10927# a_49402_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21348 a_3112_19319# a_3325_18543# a_3254_19126# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X21349 VSS a_1586_36727# a_1591_36501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2135 a_12712_59343# a_11251_59879# a_12621_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X21350 a_13835_36649# a_15775_36965# a_16648_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X21351 a_6435_10901# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21352 a_33734_65206# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21353 VDD a_12985_19087# a_29322_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21354 a_24394_15516# a_16746_15514# a_24302_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21355 vcm_commonmode a_16362_12504# a_21382_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21356 a_31330_18894# a_16362_18528# a_31422_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21357 a_39188_38341# a_38315_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21358 VDD a_75728_40202# a_75541_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21359 a_47394_19898# a_11067_67279# a_47886_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2136 a_34434_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21360 a_3803_35523# a_2216_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21361 a_11613_59049# a_11521_58951# a_11115_59317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21362 a_7467_57863# a_3295_62083# a_7812_57711# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X21363 a_12712_62313# a_11067_13095# a_12539_62063# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21364 vcm_commonmode a_16362_62194# a_46482_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21365 a_23694_57174# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21366 VSS a_1915_51946# a_1867_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21367 a_30722_58178# a_12901_58799# a_30326_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21368 VDD a_6519_65301# a_1823_76181# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21369 a_29322_63198# a_12981_62313# a_29814_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2137 VSS a_12981_59343# a_20682_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21370 a_5637_12675# a_4812_13879# a_5546_12675# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21371 a_11587_65327# a_11141_65327# a_11491_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21372 VDD a_21267_52047# a_22094_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X21373 a_28410_14512# a_16746_14510# a_28318_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21374 vcm_commonmode a_16362_11500# a_25398_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21375 VDD a_4036_51157# a_1586_51335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21376 a_5346_33775# a_4999_33781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X21377 a_4549_52271# a_4514_52523# a_4311_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21378 a_35438_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21379 a_9913_49917# a_9869_49525# a_9747_49929# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2138 a_47790_60186# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21380 a_24794_19500# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21381 a_2121_64239# a_1643_64213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21382 a_3697_35523# a_2011_34837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21383 vcm_commonmode a_16362_64202# a_37446_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21384 a_42770_23914# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21385 a_2834_36495# a_1757_36501# a_2672_36873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21386 a_39362_22910# a_16362_22544# a_39454_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21387 a_12821_51183# a_12755_51562# a_12749_51183# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21388 a_43470_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21389 a_27067_31849# a_13357_32143# a_26985_31605# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2139 a_46482_58178# a_16746_58180# a_46390_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21390 a_28318_69222# a_12901_66959# a_28810_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21391 a_2781_51183# a_1591_51183# a_2672_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X21392 a_39758_67214# a_12727_67753# a_39362_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21393 a_9204_15113# a_8123_14741# a_8857_14709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21394 a_32826_67536# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21395 a_32334_57174# a_16362_57174# a_32426_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21396 a_5185_13967# a_4995_13103# a_4866_13967# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X21397 VSS a_12899_10927# a_48794_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21398 a_17668_49007# a_16753_49007# a_17321_49249# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21399 a_2882_64605# a_2163_64381# a_2319_64476# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X214 a_5710_12675# a_4429_14191# a_5637_12675# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X2140 vcm_commonmode VSS a_43470_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21400 VDD a_35683_50613# a_35495_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21401 VSS a_10515_23975# a_32730_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21402 a_29414_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21403 a_12584_25935# a_9670_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21404 a_41766_70226# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21405 a_28441_36389# a_28195_35327# a_29127_35561# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X21406 a_40458_68218# a_16746_68220# a_40366_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21407 a_6725_42479# a_6559_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21408 a_4255_59049# a_3016_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21409 a_10400_69513# a_9485_69141# a_10053_69109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2141 a_47790_19898# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21410 a_38358_7850# VDD a_38850_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21411 a_36833_50345# a_30928_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21412 a_7794_53903# a_7749_55535# a_7637_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21413 a_19678_24918# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21414 a_25702_17890# a_12899_11471# a_25306_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21415 a_23929_47381# a_23763_47381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21416 a_49798_13874# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21417 a_1761_52815# a_1591_52815# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X21418 a_23298_55166# VSS a_23790_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21419 a_33727_38007# a_32795_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2142 a_17366_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21420 a_24515_36965# a_23749_36929# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X21421 a_1761_31055# a_1591_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21422 a_6361_44655# a_5823_44905# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21423 vcm_commonmode a_16362_61190# a_22386_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21424 VDD a_12901_58799# a_30326_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21425 VSS a_12727_15529# a_26706_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21426 a_23694_10862# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21427 a_42709_29199# a_30565_30199# a_42721_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21428 a_33015_36161# a_30757_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21429 a_30722_11866# a_12985_16367# a_30326_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2143 a_30080_36391# a_29207_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X21430 VDD a_12947_71576# a_17274_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21431 VDD a_5447_56860# a_5378_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21432 a_35438_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21433 VSS config_1_in[8] a_1591_6031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21434 a_48794_60186# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21435 a_47486_58178# a_16746_58180# a_47394_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21436 a_42374_8854# a_16362_8488# a_42466_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21437 a_48794_19898# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21438 VSS a_10975_66407# a_38754_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21439 a_9490_56873# a_8132_53511# a_9187_56597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2144 a_29414_68218# a_16746_68220# a_29322_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21440 VSS a_4571_26677# a_7113_27253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21441 VSS a_1586_21959# a_1591_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21442 a_42770_64202# a_12355_65103# a_42374_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21443 a_36842_23516# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21444 a_36442_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21445 a_40858_72556# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21446 VDD a_12985_7663# a_40366_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21447 a_32862_27247# a_24959_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21448 a_33705_27497# a_22015_28111# a_30764_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X21449 VDD a_10975_66407# a_39362_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2145 vcm_commonmode a_16362_65206# a_26402_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21450 a_2672_30345# a_1757_29973# a_2325_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21451 a_43470_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21452 a_49894_22512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21453 a_40366_62194# a_16362_62194# a_40458_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21454 a_7692_10383# a_7255_10357# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21455 a_9943_69135# a_9319_69141# a_9835_69513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21456 a_39454_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21457 a_32730_56170# a_12257_56623# a_32334_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21458 a_9414_10383# a_9219_11471# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21459 a_28410_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2146 a_3301_27791# a_2473_34293# a_3229_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X21460 a_9263_24501# a_9955_21807# a_10767_20495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21461 a_23298_72234# VSS a_23390_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21462 a_28714_63198# a_15439_49525# a_28318_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21463 VSS a_12727_58255# a_25702_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21464 VSS a_11067_67279# a_25702_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21465 a_23790_7452# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21466 a_12369_37253# a_12677_36893# a_12343_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X21467 a_39854_14480# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21468 a_39758_20902# a_11067_67279# a_39362_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21469 VDD a_1591_36103# a_1591_35951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2147 a_31726_24918# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21470 VSS a_1923_73087# a_5497_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21471 a_37354_15882# a_16362_15516# a_37446_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21472 VDD a_10055_58791# a_43378_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21473 a_18672_38567# a_17799_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21474 a_41462_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21475 VDD a_11067_21583# a_26310_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21476 vcm_commonmode VSS a_46482_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21477 VSS a_12677_42333# a_12369_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21478 a_12621_36091# a_35647_35877# a_36520_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X21479 a_10221_74031# a_10055_74031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2148 a_28318_23914# a_16362_23548# a_28410_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21480 VDD a_7580_61751# a_7755_68591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21481 VDD a_6775_53877# a_6733_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21482 a_30418_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21483 vcm_commonmode a_16362_23548# a_36442_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21484 a_39468_37479# a_38499_37503# a_39431_37737# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X21485 VDD a_10975_66407# a_12899_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21486 a_40458_21540# a_16746_21538# a_40366_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21487 VSS a_14425_37981# a_14117_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21488 VSS config_2_in[14] a_1591_50639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21489 a_12371_53903# a_12120_54019# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2149 a_42466_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21490 VDD a_12985_16367# a_47394_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21491 a_19769_38793# a_19703_38695# a_12889_39889# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21492 VDD a_12901_66959# a_37354_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21493 a_17274_63198# a_16362_63198# a_17366_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21494 a_23535_50247# a_23631_50069# a_23933_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21495 a_38754_68218# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21496 a_31422_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21497 VSS a_2223_28617# a_3983_24233# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21498 a_27406_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21499 a_10400_69513# a_9319_69141# a_10053_69109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X215 VSS a_15548_30761# a_5363_30503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X2150 VDD a_10975_66407# a_38358_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21500 VDD a_4676_47607# a_4491_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21501 a_4065_74281# a_3978_74183# a_3275_73658# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21502 a_7565_31751# a_7295_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X21503 vcm_commonmode a_16362_67214# a_29414_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21504 a_17766_10464# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21505 a_31330_7850# VSS a_31422_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21506 a_11999_67477# a_11711_67325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21507 a_38850_64524# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21508 a_35346_61190# a_12981_59343# a_35838_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21509 a_32334_20902# a_16362_20536# a_32426_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2151 a_35838_62516# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21510 a_43378_69222# a_16362_69222# a_43470_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21511 VDD a_12981_62313# a_42374_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21512 VSS a_12257_56623# a_45782_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21513 a_36193_31375# a_32823_29397# a_36097_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21514 vcm_commonmode a_16362_59182# a_19374_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21515 a_14088_35279# a_13097_36367# a_13867_35606# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21516 VDD a_5239_65301# a_5226_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21517 VDD a_37699_27221# a_38606_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21518 VDD a_6435_47893# a_6422_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21519 a_23390_57174# a_16746_57176# a_23298_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2152 a_28152_44869# a_27183_44581# a_28056_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X21520 a_24698_18894# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21521 a_7494_46287# a_7368_46403# a_7090_46419# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X21522 a_11049_71855# a_10883_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21523 a_32641_43777# a_12357_37999# a_32555_43777# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X21524 a_47486_11500# a_16746_11498# a_47394_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21525 a_22951_52271# a_22921_52245# a_6775_53877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X21526 VSS a_7289_70767# a_7805_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21527 VDD a_12895_13967# a_46390_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21528 a_16831_51183# a_16385_51183# a_16735_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21529 a_39362_60186# a_12727_58255# a_39854_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2153 a_9215_58487# a_8592_58255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X21530 a_9970_56445# a_5682_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21531 a_31422_7484# VDD a_31330_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21532 a_20378_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21533 a_15775_34239# a_14076_35077# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X21534 a_47394_68218# a_16362_68218# a_47486_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21535 a_21519_49007# a_21003_49007# a_21424_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X21536 VDD a_14049_42869# a_14079_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21537 VDD a_15439_49525# a_28318_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21538 a_19410_43439# a_19233_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21539 a_12901_66665# a_11067_66191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2154 a_48890_22512# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21540 a_30602_50345# a_27869_50095# a_30520_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21541 VDD a_10751_59575# a_10649_58947# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X21542 a_6277_14191# a_2004_42453# a_6059_14165# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21543 a_9217_53135# a_7803_55509# a_7217_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21544 a_41462_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21545 VSS a_5877_70197# a_6791_70455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21546 a_29322_71230# a_12901_66665# a_29814_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21547 a_24394_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21548 a_2250_64605# a_2163_64381# a_1846_64491# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21549 a_40429_37479# a_40737_37692# a_40403_37683# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X2155 VSS a_28426_29941# a_12263_4391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X21550 a_41862_17492# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21551 a_41766_23914# a_10515_23975# a_41370_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21552 a_9585_68841# a_8782_65015# a_9503_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21553 a_32121_42369# a_32795_42943# a_33727_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X21554 a_21290_24918# VSS a_21782_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21555 VDD config_2_in[4] a_1591_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X21556 VSS a_35196_35425# a_36395_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21557 a_6579_42255# a_6607_42167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21558 VSS a_12202_54599# a_12120_54019# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21559 VSS a_5079_35639# a_4999_33781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2156 a_38450_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21560 a_5226_46109# a_4149_45743# a_5064_45743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21561 VDD a_19517_31751# a_18328_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X21562 VSS a_23901_42044# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21563 a_4533_55799# a_1823_58773# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21564 vcm_commonmode VSS a_37446_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21565 VDD a_3327_9308# a_9179_13737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21566 VSS a_21479_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21567 a_27406_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21568 a_8592_58255# a_7963_58255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21569 a_41462_70226# a_16746_70228# a_41370_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2157 VSS a_12907_56399# a_16362_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X21570 VSS a_24937_39306# a_12801_38517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21571 VDD a_2847_18517# a_2834_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21572 a_11400_26133# a_11251_26159# a_11696_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21573 a_44778_56170# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21574 a_38754_21906# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21575 a_42374_13874# a_12727_15529# a_42866_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21576 VSS a_2787_32679# a_7390_32693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21577 a_27710_66210# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21578 a_8753_31055# a_8215_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21579 a_4748_52637# a_4311_52245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2158 a_22294_72234# VSS a_22386_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21580 VSS a_11067_13095# a_31726_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21581 a_45878_55488# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21582 a_25306_23914# a_12947_23413# a_25798_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21583 a_25306_19898# a_16362_19532# a_25398_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21584 a_23501_42583# a_23597_42325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21585 a_35478_27791# a_19807_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21586 a_37446_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21587 VDD a_35676_49525# a_36280_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21588 vcm_commonmode a_16362_20536# a_29414_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21589 a_26321_50095# a_26155_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2159 a_27710_63198# a_15439_49525# a_27314_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21590 a_32334_65206# a_16362_65206# a_32426_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21591 a_35742_14878# a_12727_15529# a_35346_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21592 a_44474_61190# a_16746_61192# a_44382_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21593 a_28318_55166# VSS a_28410_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21594 vcm_commonmode a_16362_17524# a_41462_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21595 a_33635_47695# a_22015_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21596 VSS a_12947_56817# a_21686_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21597 a_18770_18496# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21598 a_18674_24918# a_18007_27441# a_18278_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21599 a_27406_71230# a_16746_71232# a_27314_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X216 a_8902_36469# a_8017_36495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X2160 a_18370_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21600 VDD a_12727_13353# a_22294_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21601 a_48794_13874# a_12877_16911# a_48398_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21602 VSS a_12985_16367# a_45782_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21603 vcm_commonmode a_16362_12504# a_19374_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21604 a_28318_14878# a_12877_14441# a_28810_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21605 a_12196_21583# a_12166_21501# a_12093_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21606 a_23390_10496# a_16746_10494# a_23298_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21607 a_29322_18894# a_16362_18528# a_29414_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21608 a_32826_12472# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21609 a_6956_65693# a_6519_65301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2161 VSS a_12727_58255# a_24698_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21610 a_30326_13874# a_16362_13508# a_30418_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21611 a_49402_68218# a_12727_67753# a_49894_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21612 a_2107_21807# a_1757_21807# a_2012_21807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21613 VSS a_8273_42479# a_10648_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21614 a_5957_47919# a_5913_48161# a_5791_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X21615 a_23934_48783# a_22989_48437# a_23767_48463# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X21616 a_75445_39738# a_75541_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21617 a_48490_60186# a_16746_60188# a_48398_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21618 a_4035_54965# a_4238_55123# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21619 a_48490_19532# a_16746_19530# a_48398_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2162 a_20378_55166# VDD a_20286_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21620 vcm_commonmode a_16362_16520# a_45478_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21621 a_3705_73461# a_3487_73865# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X21622 VDD a_9083_13879# a_10421_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21623 a_26319_36341# a_26495_36341# a_26447_36367# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21624 a_32426_24552# VDD a_32334_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21625 a_26447_41807# a_12641_42036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21626 VDD a_9204_15113# a_9379_15039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21627 a_2325_38645# a_2107_39049# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21628 a_2847_15039# a_2672_15113# a_3026_15101# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21629 VDD a_12139_18517# a_12126_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2163 a_21686_16886# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21630 a_45478_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21631 VDD a_5749_18297# a_5779_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21632 a_12983_63151# a_12710_63151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21633 a_26417_47919# a_25879_48169# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21634 a_26802_68540# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21635 vcm_commonmode a_16362_18528# a_18370_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21636 VDD a_12983_63151# a_30326_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21637 a_12683_51329# a_12993_50345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X21638 a_22386_16520# a_16746_16518# a_22294_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21639 VDD a_4215_51157# a_23763_47381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2164 VSS a_11067_67279# a_24698_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X21640 a_35438_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21641 a_12353_20969# a_12323_20904# a_12263_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X21642 a_11759_51959# a_11855_51959# a_12157_52047# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21643 a_3203_17620# a_3063_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21644 a_22352_37253# a_21479_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21645 a_25263_38825# a_24331_38591# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21646 a_4625_50613# a_4407_51017# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21647 a_35742_9858# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21648 a_15557_52245# a_15892_51843# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X21649 a_21686_58178# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2165 a_12869_2741# a_22026_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X21650 a_35742_71230# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21651 a_34434_69222# a_16746_69224# a_34342_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21652 VSS a_17682_50095# a_32396_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21653 VSS a_30855_41809# a_30801_41835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21654 a_29715_49667# a_29055_49525# a_29643_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21655 a_42770_72234# VDD a_42374_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21656 a_2279_33775# a_1915_35015# a_1916_33927# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X21657 a_9972_69831# a_1586_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21658 a_27314_64202# a_11067_13095# a_27806_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21659 a_31822_62516# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2166 a_9485_69141# a_9319_69141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21660 VSS a_12546_22351# a_45782_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21661 a_2497_53903# a_2327_53903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X21662 a_39454_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21663 a_16244_34973# a_15775_34239# a_16648_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X21664 a_36350_60186# a_16362_60186# a_36442_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21665 a_6435_74005# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21666 VDD a_2672_40303# a_2847_40277# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21667 a_17274_56170# a_12947_56817# a_17766_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21668 a_39758_70226# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21669 a_38450_68218# a_16746_68220# a_38358_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2167 VSS a_18703_29199# a_40219_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X21670 vcm_commonmode a_16362_65206# a_35438_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21671 a_1881_72943# a_1846_73195# a_1643_72917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21672 a_40762_24918# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21673 a_37354_23914# a_16362_23548# a_37446_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21674 VSS a_4987_52508# a_4918_52637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21675 VDD a_15259_46805# a_12355_65103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21676 vcm_commonmode a_16362_64202# a_48490_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21677 VDD a_12546_22351# a_39362_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21678 VDD a_7311_60975# a_7573_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21679 a_10755_16367# a_10239_16367# a_10660_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X2168 VDD a_11035_47893# a_7571_26151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21680 VDD a_5594_36727# a_5547_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X21681 a_2583_68047# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21682 VSS a_11619_56615# a_12565_9633# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21683 a_19629_39631# a_19203_39958# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21684 a_4701_43567# a_4535_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21685 VSS a_12727_58255# a_33734_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21686 a_22448_39429# a_21479_39141# a_22411_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X21687 VSS a_11067_67279# a_33734_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21688 a_14167_30083# a_12935_31287# a_14095_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21689 a_26155_30083# a_7939_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2169 a_38850_14480# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21690 vcm_commonmode a_16362_56170# a_38450_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21691 a_31898_30761# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21692 a_2601_72105# a_2571_72040# a_2322_72631# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X21693 a_30326_58178# a_16362_58178# a_30418_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21694 a_44382_71230# a_16362_71230# a_44474_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21695 VDD a_15069_35805# a_14675_35831# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21696 VDD a_13909_38659# a_26445_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X21697 a_43774_15882# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21698 VSS a_12895_13967# a_46786_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21699 a_22014_30761# a_20881_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X217 VSS a_10391_49855# a_6831_63303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X2170 a_38754_20902# a_11067_67279# a_38358_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21700 a_25398_64202# a_16746_64204# a_25306_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21701 VDD a_19096_36513# a_18197_36604# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X21702 a_2250_59343# a_2124_59459# a_1846_59475# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X21703 a_30326_17890# a_12899_10927# a_30818_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21704 VSS a_12947_23413# a_30722_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21705 a_29943_34789# a_29177_34753# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X21706 a_27406_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21707 a_8815_13879# a_1929_10651# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21708 VDD a_12355_15055# a_34342_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21709 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2171 a_11617_18785# a_11399_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X21710 a_18278_8854# a_12985_19087# a_18770_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21711 VSS a_12981_59343# a_19678_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21712 a_13669_35253# a_33015_36161# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X21713 VDD a_8080_47607# a_6727_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21714 a_21382_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21715 vcm_commonmode a_16362_9492# a_37446_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21716 a_22639_50639# a_22015_50645# a_22531_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21717 VSS a_12727_13353# a_20682_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21718 a_23694_18894# a_12899_10927# a_23298_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21719 a_47790_14878# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2172 VDD a_5964_35015# a_4123_37013# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21720 a_30722_9858# a_12985_19087# a_30326_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21721 VSS a_9063_71553# a_9024_71427# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21722 vcm_commonmode a_16362_70226# a_30418_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21723 a_9123_57399# a_7210_55081# a_9290_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21724 a_38850_72556# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21725 a_2121_63151# a_1643_63125# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21726 a_47486_9492# a_16746_9490# a_47394_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21727 VDD a_12901_66665# a_42374_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21728 VDD a_12981_59343# a_38358_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21729 a_41462_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2173 VDD a_10055_58791# a_42374_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21730 vcm_commonmode a_16362_62194# a_20378_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21731 VDD a_26661_34428# a_26267_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21732 a_30809_51433# a_28968_50871# a_30375_51335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21733 a_21290_58178# a_10515_22671# a_21782_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21734 a_19374_55166# VDD a_19282_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21735 a_5009_56623# a_4974_56875# a_4771_56597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21736 VSS a_12877_14441# a_24698_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21737 a_21686_11866# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21738 VSS a_29269_40741# a_30875_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21739 a_18278_10862# a_16362_10496# a_18370_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2174 VDD VDD a_23298_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21740 vcm_commonmode a_16362_61190# a_33430_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21741 VDD a_6072_56872# a_6010_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21742 a_34434_22544# a_16746_22542# a_34342_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21743 a_12723_17231# a_11251_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21744 VSS a_1929_12131# a_8167_11561# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21745 a_8636_63669# a_7155_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21746 a_6473_67825# a_6224_73095# a_5964_67655# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21747 a_6743_23555# a_4427_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21748 VDD a_10400_69513# a_10575_69439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21749 a_5791_47919# a_5345_47919# a_5695_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2175 VSS a_10055_58791# a_12901_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X21750 VDD a_12947_71576# a_28318_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21751 VSS a_12983_63151# a_36746_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21752 VDD a_27937_27247# a_28589_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X21753 a_3779_25731# a_3325_18543# a_3707_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21754 a_40762_65206# a_10975_66407# a_40366_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21755 a_2325_10081# a_2107_9839# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21756 a_3392_37949# a_2952_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21757 a_2882_63517# a_2163_63293# a_2319_63388# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21758 a_28410_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21759 VSS a_10975_66407# a_49798_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2176 a_4612_57961# a_3877_57167# a_4357_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X21760 a_14293_41807# a_13867_42134# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21761 a_38450_21540# a_16746_21538# a_38358_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21762 a_47886_23516# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21763 a_37307_51339# a_36821_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21764 a_47486_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21765 VSS a_2244_22583# a_2021_22325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21766 VDD a_22577_29111# a_23498_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21767 a_4553_64213# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X21768 a_19626_31751# a_18829_29423# a_19789_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21769 VSS a_12585_39069# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X2177 a_33261_51433# a_4482_57863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X21770 a_43774_56170# a_12257_56623# a_43378_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21771 a_37846_15484# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21772 a_29545_40193# a_28931_39679# a_29863_39913# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X21773 VDD a_12877_16911# a_41370_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21774 a_26706_66210# a_12983_63151# a_26310_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21775 a_7001_36495# a_6653_36611# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X21776 a_2369_39037# a_2325_38645# a_2203_39049# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21777 a_11455_12157# a_1586_18695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21778 VDD a_10515_23975# a_24302_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21779 a_48398_15882# a_16362_15516# a_48490_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2178 VDD a_11067_21583# a_25306_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21780 vcm_commonmode a_16362_8488# a_26402_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21781 vcm_commonmode a_16362_59182# a_40458_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21782 VDD a_3305_38671# a_3813_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21783 vcm_commonmode a_16362_69222# a_23390_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21784 a_47790_55166# VSS a_47394_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21785 a_38358_11866# a_10055_58791# a_38850_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21786 VSS VDD a_31726_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21787 a_5779_75093# a_5475_74895# a_5713_74895# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X21788 VDD a_12516_7093# a_35346_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21789 a_5179_59663# a_1952_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2179 VSS a_3491_42239# a_3425_42313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X21790 VSS a_2292_43291# a_2369_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21791 a_37699_27221# a_38436_29941# a_39409_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21792 a_9225_71855# a_9183_72007# a_8539_71829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X21793 VSS a_2339_38129# a_6743_20969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21794 a_5825_36611# a_4578_40455# a_5729_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21795 VSS a_3016_60949# a_7273_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X21796 a_25398_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21797 a_9543_65327# a_9513_65301# a_9435_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21798 VSS config_1_in[15] a_1591_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X21799 VDD a_12901_66959# a_48398_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X218 a_31009_38571# a_30943_38695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2180 a_49402_14878# a_16362_14512# a_49494_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21800 a_28318_63198# a_16362_63198# a_28410_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21801 vcm_commonmode a_16362_58178# a_44474_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21802 a_18370_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21803 vcm_commonmode a_16362_68218# a_27406_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21804 a_30561_50639# a_26397_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21805 a_25199_51183# a_24683_51183# a_25104_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X21806 a_12323_20904# a_4792_20443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21807 a_36842_65528# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21808 a_4889_55535# a_4533_55799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21809 a_7829_60431# a_7449_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2181 vcm_commonmode VSS a_36442_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21810 a_49894_64524# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21811 a_46390_61190# a_12981_59343# a_46882_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21812 a_27590_50095# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21813 a_22690_60186# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21814 a_21382_58178# a_16746_58180# a_21290_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21815 VDD a_1952_60431# a_3521_57283# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21816 a_22690_19898# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21817 VSS a_12985_25615# a_16080_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21818 VSS a_12985_7663# a_36746_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21819 VSS a_16228_28335# a_17569_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2182 a_9665_51183# a_9187_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21820 a_9707_51325# a_1586_51335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21821 a_11415_58077# a_10791_57711# a_11307_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21822 a_39854_56492# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21823 a_19282_24918# VSS a_19774_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21824 a_36520_40517# a_35647_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21825 VDD a_19591_50943# a_19578_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21826 VDD a_14049_36341# a_14079_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21827 VDD a_11812_30511# a_12786_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21828 a_34738_71230# a_12947_71576# a_34342_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21829 a_23790_22512# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2183 VSS a_29913_43457# a_30415_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21830 VDD a_12355_65103# a_26310_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21831 VSS a_25939_51157# a_25873_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21832 VSS a_7000_43541# a_15259_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21833 VDD a_6138_54599# a_6095_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21834 a_4553_64213# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21835 a_4555_55233# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21836 a_7479_17607# a_7407_18038# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21837 a_2969_41909# a_2751_42313# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21838 a_2242_24893# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21839 a_4513_32259# a_2216_28309# a_4440_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 vcm_commonmode a_16362_23548# a_35438_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21840 a_28941_48801# a_26514_47375# a_28855_48801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X21841 a_27314_72234# VDD a_27806_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21842 a_38754_70226# a_12901_66665# a_38358_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21843 VSS a_2317_28892# a_3985_22901# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21844 a_31822_70548# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21845 a_24302_14878# a_16362_14512# a_24394_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21846 a_4642_54991# a_4555_55233# a_4238_55123# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21847 a_29651_48576# a_17682_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21848 VSS a_23631_50069# a_23934_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21849 a_27806_60508# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2185 a_7289_62607# a_7199_62839# a_7071_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21850 vcm_commonmode a_16362_17524# a_39454_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21851 a_43470_15516# a_16746_15514# a_43378_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21852 vcm_commonmode a_16362_12504# a_40458_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21853 VSS a_6880_58773# a_6824_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21854 a_14365_46805# a_11067_46823# a_14611_46859# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X21855 a_11049_71855# a_10883_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21856 vcm_commonmode a_16362_22544# a_23390_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21857 a_4407_51017# a_4057_50645# a_4312_51005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21858 VSS a_35602_34191# a_36147_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21859 VDD a_29361_51727# a_30843_52521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2186 a_39362_10862# a_12985_16367# a_39854_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21860 a_12202_54599# a_12231_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21861 a_42770_57174# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21862 VSS a_28959_49783# a_29561_49667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21863 vcm_commonmode VSS a_48490_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21864 a_16746_63200# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X21865 a_25702_67214# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21866 VDD a_12202_54599# a_12202_54019# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21867 VDD a_2315_24540# a_2899_28111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21868 VDD a_2672_12937# a_2847_12863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21869 vcm_commonmode a_16362_11500# a_44474_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2187 VSS a_2787_62063# a_3484_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X21870 VSS a_51714_39886# a_52590_39936# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.55e+11p ps=1.62e+06u w=500000u l=150000u
X21871 VSS a_2775_46025# a_30716_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21872 a_43870_19500# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21873 vcm_commonmode a_16362_21540# a_27406_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21874 VSS a_3417_33231# a_3983_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21875 a_11793_67325# a_11521_66567# a_11711_67325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21876 a_42466_62194# a_16746_62196# a_42374_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21877 a_2121_59709# a_1643_59317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21878 a_41159_28585# a_29175_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X21879 a_13608_51433# a_13445_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2188 vcm_commonmode a_16362_22544# a_48490_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X21880 a_25398_72234# VDD a_25306_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21881 a_46786_14878# a_12727_15529# a_46390_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21882 VSS a_9307_30663# a_10595_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21883 a_13565_44135# a_13661_43957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21884 VSS a_12947_56817# a_32730_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21885 vcm_commonmode a_16362_13508# a_17366_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21886 a_29814_18496# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21887 a_29718_24918# VSS a_29322_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21888 a_26310_15882# a_12727_13353# a_26802_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21889 a_7075_42479# a_6725_42479# a_6980_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2189 VSS a_32397_28023# a_31263_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21890 a_28065_41601# a_27999_41495# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21891 a_21382_11500# a_16746_11498# a_21290_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21892 a_29829_49257# a_28108_48463# a_29055_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X21893 a_30818_13476# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21894 VDD a_1643_54421# a_1591_54447# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X21895 a_5438_69679# a_5091_69685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X21896 a_47394_69222# a_12901_66959# a_47886_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21897 VDD a_12895_13967# a_20286_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21898 a_3705_37557# a_3487_37961# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21899 a_19678_58178# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X219 a_19596_40743# a_18627_40767# a_19559_41001# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2190 VDD a_11771_23671# a_10286_26311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X21900 VDD a_5190_59575# a_11909_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21901 a_19678_16886# a_12727_13353# a_19282_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21902 a_33430_64202# a_16746_64204# a_33338_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21903 VSS a_2122_19087# a_2228_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X21904 VSS a_18811_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21905 a_11507_72221# a_10883_71855# a_11399_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21906 a_17668_49007# a_16587_49007# a_17321_49249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21907 VDD a_12947_8725# a_38358_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21908 VSS a_12985_19087# a_34738_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21909 a_24794_69544# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2191 a_37545_51183# a_37423_51335# a_37459_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X21910 a_48490_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21911 a_21290_66210# a_10975_66407# a_21782_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21912 a_19374_63198# a_16746_63200# a_19282_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21913 a_24497_47349# a_24279_47753# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21914 a_24302_59182# a_16362_59182# a_24394_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21915 a_44778_8854# a_12947_8725# a_44382_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21916 a_12641_43124# a_12671_42134# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X21917 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X21918 a_7009_56873# a_6835_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21919 VDD a_43227_28309# a_43175_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X2192 a_29814_72556# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21920 VDD a_29847_48734# a_29651_48576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21921 a_42374_55166# VSS a_42866_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21922 a_5393_69455# a_5208_70063# a_5295_69135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X21923 a_32730_8854# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21924 a_25306_65206# a_12355_65103# a_25798_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21925 VSS a_13743_35836# a_19743_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X21926 a_2215_14735# a_1591_14741# a_2107_15113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21927 a_46786_71230# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21928 a_45478_69222# a_16746_69224# a_45386_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21929 a_4036_54421# a_1586_51335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2193 a_37750_68218# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21930 a_12335_50639# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21931 a_7921_74581# a_7755_74581# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X21932 a_29545_28023# a_16863_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21933 VDD a_10053_69109# a_9943_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21934 a_1761_40847# a_1591_40847# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X21935 a_34145_49007# a_33681_49373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21936 VSS a_4032_53047# a_3231_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X21937 VSS a_3173_66169# a_3107_66237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21938 vcm_commonmode a_16362_71230# a_24394_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21939 a_29943_39141# a_29072_38567# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X2194 a_26402_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21940 a_42770_10862# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21941 a_7260_67753# a_6224_73095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21942 VDD a_26417_47919# a_28855_48801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21943 a_36350_8854# a_16362_8488# a_36442_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21944 a_25702_20902# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21945 VSS a_12947_23413# a_28714_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21946 a_9643_63125# a_11299_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21947 a_1645_42453# a_1778_42631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21948 VDD a_28599_28023# a_24740_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X21949 VSS a_12981_59343# a_40762_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2195 VDD a_32823_29397# a_30790_30663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X21950 a_28318_56170# a_12947_56817# a_28810_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21951 a_37446_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21952 a_22352_34215# a_21479_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21953 a_13867_41807# a_13613_42134# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21954 a_49494_68218# a_16746_68220# a_49402_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21955 vcm_commonmode a_16362_65206# a_46482_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21956 a_1643_59317# a_1846_59475# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21957 VSS a_12727_13353# a_18674_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21958 a_48398_23914# a_16362_23548# a_48490_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21959 a_22690_13874# a_12877_16911# a_22294_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2196 a_2313_12015# a_1887_12342# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21960 VSS a_33008_28853# a_32952_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21961 a_19417_39958# a_19245_39747# a_19203_39958# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21962 a_8969_42233# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X21963 VSS a_12907_27023# a_36275_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21964 a_35463_36415# a_31847_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X21965 VDD a_9314_69367# a_9319_69141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X21966 a_8195_16911# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21967 a_17766_7452# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21968 vcm_commonmode a_16362_57174# a_36442_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21969 VSS a_27411_50069# a_27345_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2197 a_23298_11866# a_16362_11500# a_23390_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X21970 a_3070_67325# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21971 a_42374_72234# VSS a_42466_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21972 a_47790_63198# a_15439_49525# a_47394_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21973 VSS a_12727_58255# a_44778_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21974 VSS a_11067_67279# a_44778_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21975 a_40458_55166# VDD a_40366_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X21976 a_41766_16886# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21977 a_3621_61519# a_2959_47113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21978 a_36442_8488# a_16746_8486# a_36350_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21979 a_11764_65845# a_11521_66567# a_11987_66191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X2198 VSS a_29943_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X21980 VSS a_12516_7093# a_27710_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21981 a_19282_58178# a_10515_22671# a_19774_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21982 a_33741_32143# a_19807_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21983 a_12785_53181# a_12755_53030# a_12713_53181# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X21984 a_12901_58799# a_11067_66191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21985 VDD a_10515_23975# a_32334_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21986 VDD a_1923_59583# a_1643_63125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21987 a_5814_13967# a_4429_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21988 a_19678_11866# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21989 a_25398_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2199 VDD a_12899_10927# a_41370_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21990 a_7640_45577# a_6559_45205# a_7293_45173# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21991 vcm_commonmode a_16362_15516# a_32426_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21992 VDD a_11067_21583# a_45386_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X21993 a_39503_43957# a_39742_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X21994 a_3392_37949# a_2952_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21995 VSS a_12355_15055# a_17670_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21996 VDD a_32672_49007# a_33515_48576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21997 a_21686_60186# a_12981_59343# a_21290_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21998 a_4853_18543# a_4809_18785# a_4687_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21999 a_21686_19898# a_12895_13967# a_21290_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_43870_23516# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X220 a_28714_15882# a_12877_14441# a_28318_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2200 VDD a_40585_42369# a_42040_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X22000 a_7833_66415# a_7567_66781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22001 a_23911_35823# a_23734_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22002 VSS a_6611_14967# a_5465_14967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22003 VDD a_12727_15529# a_35346_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22004 a_2215_49551# a_1591_49557# a_2107_49929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22005 a_32426_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22006 a_10543_16580# a_10423_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22007 a_33430_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22008 VDD a_18007_27441# a_18278_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22009 a_49894_72556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2201 VDD a_12981_59343# a_29322_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22010 a_21382_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22011 VSS a_9547_54421# a_9493_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22012 a_46482_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22013 a_43378_11866# a_16362_11500# a_43470_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22014 a_37557_32463# a_31659_31751# a_37569_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22015 a_2713_31353# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X22016 VDD a_12981_59343# a_49402_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22017 a_49402_62194# a_16362_62194# a_49494_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22018 a_32334_19898# a_11067_67279# a_32826_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22019 a_12135_69109# a_11955_69653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2202 a_19435_51727# a_19576_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X22020 a_12707_26159# a_12263_26409# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X22021 VSS a_26319_42869# a_19004_40413# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22022 vcm_commonmode a_16362_62194# a_31422_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22023 a_28607_48169# a_27393_47919# a_28524_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22024 a_15661_29967# a_8753_31055# a_15443_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22025 VSS a_11763_62581# a_11395_62037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22026 a_36842_10464# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22027 a_45478_22544# a_16746_22542# a_45386_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22028 a_19774_20504# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22029 VSS a_12727_67753# a_34738_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2203 a_29322_62194# a_16362_62194# a_29414_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22030 a_19374_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22031 a_8384_40303# a_7905_40553# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X22032 VDD VDD a_26310_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22033 a_20378_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22034 a_26402_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22035 VSS a_12983_63151# a_47790_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22036 a_3707_28995# a_1915_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22037 a_13557_37999# a_13291_37999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22038 vcm_commonmode a_16362_64202# a_22386_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22039 VSS a_2657_60949# a_2605_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2204 a_30875_39095# a_29943_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X22040 a_25398_7484# VDD a_25306_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22041 a_49494_21540# a_16746_21538# a_49402_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22042 a_24302_22910# a_16362_22544# a_24394_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22043 VDD a_3024_67191# a_9953_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22044 VSS a_12901_58799# a_37750_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22045 VDD a_1923_54591# a_5132_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22046 a_41766_57174# a_10515_22671# a_41370_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22047 VDD a_2339_38129# a_2111_38279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22048 a_35838_16488# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22049 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2205 VDD a_11430_26159# a_16865_27511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5795e+11p ps=2.99e+06u w=420000u l=150000u
X22050 a_8241_10749# a_7862_10383# a_8169_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22051 a_35346_9858# a_12546_22351# a_35838_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22052 a_24698_67214# a_12727_67753# a_24302_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22053 VDD a_15439_49525# a_47394_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22054 VSS a_33203_34191# a_33309_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22055 a_39454_13508# a_16746_13506# a_39362_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22056 vcm_commonmode a_16362_10496# a_36442_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22057 a_7324_46287# a_6655_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22058 a_76082_40202# a_76178_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22059 a_45878_9460# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2206 a_42466_12504# a_16746_12502# a_42374_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22060 a_9860_65103# a_5024_67885# a_9557_64757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22061 VDD a_2143_15271# a_11793_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22062 a_7116_30287# a_5449_25071# a_6625_29941# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=2.86e+11p ps=2.18e+06u w=650000u l=150000u
X22063 a_38378_30511# a_32970_31145# a_38209_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22064 a_38754_55166# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22065 a_39115_29423# a_34759_31029# a_38436_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22066 a_17891_36189# a_14293_37455# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22067 a_43470_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22068 a_33597_27247# a_26523_28111# a_30764_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22069 VDD a_38210_30199# a_40394_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2207 VDD a_7479_17607# a_7479_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22070 VDD a_1923_59583# a_7340_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22071 a_5190_59575# a_14985_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X22072 VDD a_23643_41569# a_23467_41237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22073 a_40366_24918# VSS a_40858_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22074 a_33903_35561# a_34297_35516# a_33963_35507# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X22075 VDD a_12516_7093# a_46390_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22076 a_18674_58178# a_12901_58799# a_18278_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22077 a_46482_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22078 a_43378_56170# a_16362_56170# a_43470_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22079 a_29414_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2208 a_42887_27247# a_20359_29199# a_42718_27497# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X22080 a_26310_66210# a_16362_66210# a_26402_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22081 VDD a_6559_22671# a_8215_25071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22082 a_7407_46529# a_1586_45431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22083 a_44382_23914# a_12947_23413# a_44874_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22084 a_44382_19898# a_16362_19532# a_44474_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22085 a_15443_29941# a_8753_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22086 a_47886_65528# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22087 VDD a_2099_59861# a_18012_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22088 a_33430_72234# VDD a_33338_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22089 a_2012_68565# a_2191_68565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2209 a_21290_7850# VSS a_21382_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22090 a_5366_63695# a_4647_63937# a_4803_63669# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X22091 a_20378_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22092 a_47394_55166# VSS a_47486_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22093 a_34342_15882# a_12727_13353# a_34834_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22094 VSS a_11067_21583# a_34738_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22095 a_37750_24918# VSS a_37354_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22096 a_33734_60186# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22097 a_32426_58178# a_16746_58180# a_32334_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22098 a_33734_19898# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22099 a_1644_76181# a_1823_76181# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X221 VSS a_12877_16911# a_25702_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2210 a_6514_37191# a_4685_37583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22100 a_46482_71230# a_16746_71232# a_46390_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22101 VDD a_5993_37039# a_6559_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22102 VSS a_10975_66407# a_23694_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22103 a_37846_57496# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22104 a_35299_32375# a_36507_31573# a_36453_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22105 VDD VSS a_41370_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22106 a_7999_48841# a_7553_48469# a_7903_48841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22107 a_47394_14878# a_12877_14441# a_47886_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22108 VSS a_12985_7663# a_47790_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22109 a_21782_23516# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2211 VDD a_2775_46025# a_33748_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.345e+12p ps=1.269e+07u w=1e+06u l=150000u M=4
X22110 a_2107_12937# a_1591_12565# a_2012_12925# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X22111 VDD a_12985_19087# a_30326_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22112 a_21382_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22113 a_21856_36513# a_21663_35327# a_22595_35561# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22114 VDD a_10975_66407# a_24302_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22115 a_2781_18543# a_1591_18543# a_2672_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X22116 a_4217_44449# a_3247_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22117 VDD a_41289_36893# a_40895_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22118 a_13795_42134# a_13613_42134# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22119 a_24394_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2212 a_8258_53359# a_7803_55509# a_8168_53359# VSS sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X22120 VDD a_39459_44527# a_39565_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22121 VSS a_8453_64757# a_5595_63125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22122 a_2369_49917# a_2325_49525# a_2203_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22123 VSS a_12877_16911# a_37750_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22124 a_6514_37191# a_5631_38127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22125 a_41766_10862# a_12546_22351# a_41370_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22126 a_8480_38127# a_4685_37583# a_7948_38377# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22127 VSS a_2595_47653# a_8165_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22128 VDD a_12899_11471# a_27314_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22129 a_24794_14480# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2213 a_25398_22544# a_16746_22542# a_25306_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22130 a_24698_20902# a_11067_67279# a_24302_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22131 a_4333_29423# a_2216_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22132 a_10973_16609# a_10755_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22133 a_11981_57487# a_11883_58575# a_11763_57399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22134 a_22294_15882# a_16362_15516# a_22386_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22135 VDD a_4811_34855# a_34098_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22136 VSS a_1591_13103# a_1768_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X22137 a_49798_70226# a_12901_66665# a_49402_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22138 vcm_commonmode a_16362_18528# a_37446_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22139 a_41462_16520# a_16746_16518# a_41370_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2214 VDD a_13390_29575# a_15661_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22140 a_11987_66191# a_11710_58487# a_11893_66191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X22141 vcm_commonmode a_16362_23548# a_21382_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22142 a_75728_39738# a_75824_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22143 a_3475_9661# a_3327_9308# a_3112_9527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22144 VSS a_1591_36103# a_1591_35951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22145 a_39758_62194# a_12981_62313# a_39362_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22146 a_28810_13476# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22147 a_25306_10862# a_12985_16367# a_25798_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22148 a_46786_7850# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22149 a_40762_58178# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2215 a_77918_39826# a_75475_40594# a_77664_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22150 a_10931_52598# a_10680_52245# a_10472_52423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22151 VDD a_12901_66959# a_22294_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22152 a_23694_68218# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22153 a_39372_42919# a_38499_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22154 VDD a_38011_42035# a_38037_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22155 VDD a_12901_58799# a_18278_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22156 a_5051_43567# a_4701_43567# a_4956_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22157 a_18674_11866# a_12985_16367# a_18278_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22158 VSS a_10472_54135# a_9547_54421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22159 a_27406_17524# a_16746_17522# a_27314_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2216 a_34342_61190# a_12981_59343# a_34834_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22160 VSS a_5320_18231# a_5271_17999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22161 a_7075_49929# a_6725_49557# a_6980_49917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22162 a_40458_63198# a_16746_63200# a_40366_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22163 a_38358_70226# a_16362_70226# a_38450_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22164 a_19282_66210# a_10975_66407# a_19774_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22165 VSS a_31280_36165# a_31243_35831# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22166 VSS a_34759_31029# a_41059_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22167 a_14951_34743# a_15345_34717# a_15011_34717# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X22168 a_23790_64524# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22169 a_26706_59182# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2217 a_8399_49159# a_8143_48246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22170 a_20286_61190# a_12981_59343# a_20778_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22171 a_2939_33535# a_2764_33609# a_3118_33597# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22172 VDD a_26397_51183# a_32318_48695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22173 a_44382_8854# a_16362_8488# a_44474_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22174 VSS a_12257_56623# a_30722_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22175 a_5274_54991# a_4516_55107# a_4711_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22176 VSS a_1761_52815# a_12191_37999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22177 vcm_commonmode a_16362_13508# a_28410_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22178 VDD a_20359_29199# a_38121_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22179 a_33734_7850# VDD a_33338_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2218 a_42374_69222# a_16362_69222# a_42466_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22180 VDD start_conversion_in a_1591_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22181 a_7100_72105# a_4119_70741# a_6927_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22182 a_32426_11500# a_16746_11498# a_32334_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22183 VSS a_18811_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X22184 a_53378_39250# a_52778_39198# a_19967_41781# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22185 a_36821_50095# a_30928_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22186 a_19743_39095# a_18811_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22187 a_4429_72943# a_2686_70223# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22188 VDD a_12895_13967# a_31330_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22189 a_5455_37039# a_5449_37191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2219 VSS a_12257_56623# a_44778_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22190 a_5504_37815# a_3949_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22191 a_24302_60186# a_12727_58255# a_24794_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22192 a_33430_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22193 a_32334_68218# a_16362_68218# a_32426_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22194 VDD a_7313_53047# a_7079_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22195 a_44474_64202# a_16746_64204# a_44382_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22196 VSS a_5767_31573# a_5547_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22197 VDD a_26319_35253# a_15968_36061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22198 a_8539_71829# a_9183_72007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22199 a_46482_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X222 VSS a_12981_62313# a_37750_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2220 a_38358_16886# a_12899_11471# a_38850_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22200 a_2215_66781# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22201 VSS VDD a_31726_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22202 a_10661_10383# a_10259_10703# a_10497_10703# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X22203 VSS a_12981_59343# a_38754_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22204 a_34434_56170# a_16746_56172# a_34342_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22205 a_35742_17890# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22206 a_24698_9858# a_12985_19087# a_24302_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22207 VDD a_4215_51157# a_22015_50645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22208 vcm_commonmode VSS a_48490_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22209 a_42770_18894# a_12899_10927# a_42374_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2221 VDD a_25939_51157# a_26397_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X22210 a_17366_66210# a_16746_66212# a_17274_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22211 a_49798_24918# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22212 a_19374_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22213 VSS a_29072_38567# a_29035_38825# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X22214 a_24305_31171# a_23626_31573# a_24223_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22215 a_2672_51183# a_1757_51183# a_2325_51425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22216 VSS a_10103_11079# a_9455_11079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22217 a_35438_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22218 a_39742_44527# a_39565_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22219 a_40366_58178# a_10515_22671# a_40858_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2222 VSS a_12983_63151# a_27710_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22220 a_38450_55166# VDD a_38358_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22221 VDD a_3667_60405# a_1823_62589# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22222 a_39758_16886# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22223 vcm_commonmode VSS a_22386_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22224 VSS a_12877_14441# a_43774_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22225 a_2191_68565# a_2847_44629# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22226 a_40762_11866# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22227 a_37354_10862# a_16362_10496# a_37446_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22228 a_8203_23145# a_5085_23047# a_8009_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X22229 a_8121_48437# a_7903_48841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2223 VDD a_2223_28617# a_3955_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22230 VSS VSS a_26706_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22231 a_10860_47919# a_9945_47919# a_10513_48161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22232 a_23694_21906# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22233 a_9305_53511# a_9240_53877# a_9468_53609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22234 a_26310_57174# a_12257_56623# a_26802_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22235 a_33338_7850# VSS a_33430_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22236 a_35438_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22237 a_11053_62607# a_10575_62911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22238 VDD a_14919_37683# a_14425_37981# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X22239 VDD a_12947_71576# a_47394_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2224 a_31726_65206# a_10975_66407# a_31330_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22240 a_30818_55488# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22241 VSS a_4681_13621# a_4629_13647# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22242 a_41820_41501# a_41443_41855# a_42375_42089# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X22243 VDD a_5595_12167# a_5399_13255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X22244 VSS a_13669_35253# a_30267_35253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22245 a_20682_14878# a_12727_15529# a_20286_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22246 a_6798_16367# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22247 a_40458_9492# a_16746_9490# a_40366_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22248 VSS a_12727_13353# a_29718_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22249 a_26706_12870# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2225 a_46482_11500# a_16746_11498# a_46390_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22250 a_38754_63198# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22251 VSS a_12985_16367# a_30722_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22252 a_4461_48981# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X22253 a_9651_67503# a_9301_67503# a_9556_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22254 a_26447_39141# a_25300_39655# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X22255 VDD a_1923_54591# a_1643_56597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22256 VDD a_4001_56377# a_4031_56118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22257 a_32730_67214# a_12727_67753# a_32334_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22258 a_17274_59182# a_12901_58799# a_17766_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22259 a_14258_34191# a_14081_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2226 VSS a_5612_58229# a_5550_58255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22260 a_30007_38695# a_30115_38695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22261 VDD a_3173_66169# a_3203_65910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22262 a_10299_47607# a_4443_46607# a_10473_47713# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X22263 a_28513_29673# a_4811_34855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22264 a_45782_66210# a_12983_63151# a_45386_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22265 vcm_commonmode a_16362_62194# a_29414_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22266 a_36350_22910# a_10515_23975# a_36842_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22267 a_6725_42479# a_6559_42479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22268 VDD a_10515_23975# a_43378_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22269 a_8485_29423# a_6752_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2227 VDD a_12895_13967# a_45386_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22270 vcm_commonmode a_16362_16520# a_30418_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22271 a_40858_20504# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22272 a_40458_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22273 VDD a_31959_34751# a_31819_35073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22274 a_7544_32937# a_6883_37019# a_7472_32937# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22275 a_43378_64202# a_16362_64202# a_43470_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22276 a_3137_37589# a_2971_37589# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22277 a_18370_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22278 a_14859_37737# a_15253_37692# a_14919_37683# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X22279 a_1761_37039# a_1591_37039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2228 a_29414_21540# a_16746_21538# a_29322_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22280 a_30418_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22281 VDD a_12877_14441# a_33338_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22282 vcm_commonmode a_16362_69222# a_42466_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22283 VDD a_19580_49159# a_19531_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22284 a_32831_35307# a_30757_37455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22285 VDD a_12727_15529# a_46390_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22286 a_44474_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22287 a_7162_59575# a_6737_60431# a_7299_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22288 a_41370_12870# a_16362_12504# a_41462_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22289 a_20378_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2229 VSS a_22243_30491# a_21879_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X22290 VDD VSS a_29322_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22291 a_47394_63198# a_16362_63198# a_47486_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22292 a_34342_66210# a_16362_66210# a_34434_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22293 a_12599_42134# a_12417_42134# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22294 a_9425_51183# a_9390_51435# a_9187_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22295 a_20682_71230# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22296 a_34834_11468# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22297 a_38315_39141# a_36708_39655# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X22298 VSS a_11067_13095# a_19678_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22299 VSS a_32167_29611# a_32397_28023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X223 VSS a_19780_39429# a_19743_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2230 a_5553_33231# a_1689_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X22300 VDD a_1586_40455# a_1775_47381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22301 a_17766_21508# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22302 a_17366_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22303 a_2885_39759# a_1689_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X22304 a_3491_42239# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22305 a_4067_15797# a_3911_16065# a_4212_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22306 a_47886_10464# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22307 VDD a_28426_29941# a_12263_4391# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22308 a_15660_49257# a_11067_13095# a_15483_49007# VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X22309 a_24394_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2231 VSS a_12901_58799# a_17670_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22310 VSS a_2419_48783# a_9913_49917# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22311 a_21290_60186# a_16362_60186# a_21382_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22312 VSS a_12727_67753# a_45782_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22313 a_39454_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22314 VSS a_25517_37455# a_41999_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22315 a_24698_70226# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22316 a_23390_68218# a_16746_68220# a_23298_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22317 vcm_commonmode a_16362_59182# a_49494_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22318 vcm_commonmode a_16362_65206# a_20378_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22319 a_13692_44527# a_13515_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2232 a_28648_50101# a_4351_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X22320 a_4935_70561# a_2952_66139# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X22321 a_22294_23914# a_16362_23548# a_22386_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22322 VDD a_10975_66407# a_32334_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22323 a_8123_28879# a_5087_29423# a_8206_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22324 a_12587_51335# a_2840_66103# a_12821_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22325 a_28056_40517# a_27183_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22326 vcm_commonmode a_16362_64202# a_33430_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22327 a_18278_13874# a_16362_13508# a_18370_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22328 VDD a_12546_22351# a_24302_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22329 a_38358_63198# a_12981_62313# a_38850_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2233 a_4985_61021# a_1823_62589# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22330 VDD a_8635_61751# a_8039_61493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X22331 a_27139_31849# a_25321_29673# a_27067_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22332 a_40675_27791# a_40402_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22333 VDD a_12355_65103# a_45386_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22334 a_42866_61512# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22335 a_2325_66657# a_2107_66415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22336 a_3357_22649# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X22337 a_37446_14512# a_16746_14510# a_37354_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22338 a_4461_48981# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22339 VSS a_30557_49783# a_30525_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2234 a_2405_20719# a_2228_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22340 a_8397_35727# a_5915_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22341 a_27710_61190# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22342 a_26402_59182# a_16746_59184# a_26310_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22343 vcm_commonmode a_16362_56170# a_23390_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22344 a_4681_13621# a_5227_13621# a_5185_13967# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22345 a_32730_20902# a_11067_67279# a_32334_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22346 VSS a_12895_13967# a_31726_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22347 VDD a_12257_56623# a_35346_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22348 VDD a_1586_40455# a_3983_48469# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22349 VDD a_12983_63151# a_18278_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2235 VSS a_38171_43983# a_38277_43983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22350 VDD a_17321_49249# a_17211_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22351 a_7090_46419# a_7407_46529# a_7365_46653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22352 a_46882_60508# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22353 VSS a_26523_28111# a_33688_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22354 a_18370_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22355 a_7373_40847# a_7107_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22356 vcm_commonmode VSS a_27406_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22357 VSS a_6072_56872# a_6010_56989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22358 a_2012_71677# a_1895_71482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22359 a_32730_14878# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2236 a_21382_7484# VDD a_21290_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22360 VSS a_11851_64391# a_11803_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22361 vcm_commonmode a_16362_22544# a_42466_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22362 a_6753_51183# a_5909_51433# a_6671_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22363 VSS a_13716_43047# a_17939_43745# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22364 a_23790_72556# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22365 a_41370_57174# a_16362_57174# a_41462_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22366 a_19774_62516# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22367 a_37750_9858# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22368 a_29718_58178# a_12901_58799# a_29322_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22369 VDD a_12355_65103# a_12899_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2237 a_2497_61519# a_2141_61635# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22370 VDD a_12981_59343# a_23298_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22371 a_44778_67214# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22372 a_8544_15101# a_8361_15529# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X22373 VDD a_23749_36929# a_24928_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X22374 a_12875_31751# a_8461_32937# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22375 a_36107_36965# a_34699_37683# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X22376 VSS a_12546_22351# a_47790_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22377 VSS a_9491_12297# a_10433_12879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22378 a_43353_27791# a_23395_32463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22379 a_34738_59182# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2238 a_21686_57174# a_10515_22671# a_21290_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22380 a_7737_74031# a_6098_73095# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22381 VDD a_4417_22671# a_9167_24011# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22382 a_34738_17890# a_12899_11471# a_34342_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22383 a_17670_69222# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22384 a_44474_72234# VDD a_44382_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22385 VSS a_12983_63151# a_21686_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22386 a_13867_38870# a_13909_38659# a_13867_38543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22387 a_48890_18496# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22388 a_45386_15882# a_12727_13353# a_45878_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22389 VSS a_11067_21583# a_45782_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2239 a_28143_52105# a_27793_51733# a_28048_52093# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X22390 VSS a_33641_29967# a_40967_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22391 VDD a_19807_28111# a_33705_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22392 vcm_commonmode a_16362_23548# a_19374_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22393 a_2461_52271# a_2417_52513# a_2295_52271# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22394 vcm_commonmode a_16362_12504# a_49494_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22395 a_23390_21540# a_16746_21538# a_23298_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22396 a_18278_58178# a_16362_58178# a_18370_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22397 a_32826_23516# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22398 a_11525_57953# a_11307_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22399 a_32426_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X224 a_4674_40277# a_7756_19087# a_6743_19881# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.99e+12p ps=2.398e+07u w=1e+06u l=150000u M=4
X2240 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22400 a_33484_39429# a_32611_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22401 a_38754_16886# a_12727_13353# a_38358_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22402 VSS a_12727_15529# a_35742_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22403 VSS a_15607_46805# a_40599_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22404 a_3801_24643# a_2315_24540# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22405 a_15074_50871# a_7050_53333# a_15211_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22406 VSS a_6619_16341# a_6553_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22407 a_18278_17890# a_12899_10927# a_18770_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22408 a_6216_28335# a_6162_28487# a_6096_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22409 a_11266_10205# a_11140_10107# a_10862_10091# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=360000u l=150000u
X2241 a_5156_18543# a_4075_18543# a_4809_18785# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X22410 a_22786_15484# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22411 VDD a_12899_10927# a_25306_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22412 a_11617_18785# a_11399_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22413 a_2215_38671# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22414 a_7815_45503# a_7640_45577# a_7994_45565# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22415 a_1644_62581# a_1823_62589# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22416 a_10571_74031# a_10221_74031# a_10476_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22417 a_43870_69544# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22418 a_40366_66210# a_10975_66407# a_40858_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22419 a_26402_12504# a_16746_12502# a_26310_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2242 a_30267_35253# a_13669_35253# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22420 a_6375_64489# a_4119_70741# a_6457_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22421 a_38450_63198# a_16746_63200# a_38358_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22422 vcm_commonmode a_16362_60186# a_35438_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22423 vcm_commonmode a_16362_19532# a_35438_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22424 a_39854_59504# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22425 VDD a_7293_45173# a_7183_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22426 a_33338_15882# a_16362_15516# a_33430_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22427 a_31543_51335# a_32091_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22428 a_36797_27497# a_32367_28309# a_36643_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22429 vcm_commonmode a_16362_70226# a_18370_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2243 VDD a_15439_49525# a_27314_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22430 a_11955_69653# a_11780_69679# a_12134_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22431 vcm_commonmode a_16362_18528# a_48490_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22432 VDD a_9011_74879# a_8998_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22433 VSS a_12257_56623# a_28714_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22434 vcm_commonmode a_16362_9492# a_39454_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22435 a_19559_41001# a_18627_40767# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22436 a_23298_11866# a_10055_58791# a_23790_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22437 a_26706_8854# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22438 a_41427_52263# a_41059_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22439 VDD a_12516_7093# a_20286_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2244 a_2250_54813# a_2163_54589# a_1846_54699# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X22440 a_44382_65206# a_12355_65103# a_44874_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22441 a_49494_9492# a_16746_9490# a_49402_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22442 a_21387_39679# a_19596_40743# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X22443 a_4177_29423# a_1915_35015# a_4095_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22444 VSS a_25987_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X22445 a_43470_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22446 VSS config_2_in[3] a_1591_34319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22447 a_25398_18528# a_16746_18526# a_25306_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22448 VDD a_2451_72373# a_4065_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22449 VDD a_12901_58799# a_29322_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2245 VSS a_2847_36799# a_2216_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X22450 VDD a_4311_52245# a_1823_63677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22451 a_34342_57174# a_12257_56623# a_34834_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22452 a_26917_47919# a_26514_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X22453 a_29718_11866# a_12985_16367# a_29322_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22454 a_44778_20902# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22455 VDD a_7640_42479# a_7815_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22456 a_17274_67214# a_12983_63151# a_17766_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22457 VSS a_26417_47919# a_30165_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22458 a_21782_65528# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22459 a_47394_56170# a_12947_56817# a_47886_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2246 a_6619_16341# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22460 a_3026_40303# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22461 a_20839_44265# a_21233_44220# a_20899_44211# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X22462 VSS a_12901_66665# a_42770_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22463 VDD a_20543_46831# a_20575_47713# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22464 VDD a_18413_47919# a_19258_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22465 a_4941_35727# a_4762_35484# a_5121_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=3.04e+06u as=0p ps=0u w=1e+06u l=150000u
X22466 a_31330_61190# a_12981_59343# a_31822_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22467 a_40458_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22468 a_34738_12870# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22469 a_16832_35303# a_15959_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2247 a_7649_17455# a_7479_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22470 VDD a_12985_7663# a_39362_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22471 vcm_commonmode a_16362_14512# a_26402_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22472 VSS a_39449_39868# a_39141_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22473 a_17670_22910# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22474 a_23467_41237# a_23643_41569# a_23595_41629# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X22475 VDD a_9731_22895# a_12935_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22476 VSS a_12985_7663# a_21686_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22477 a_24794_56492# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22478 VSS a_8015_21807# a_8583_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22479 vcm_commonmode a_16362_67214# a_38450_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 a_19374_13508# a_16746_13506# a_19282_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22480 a_2751_42313# a_2235_41941# a_2656_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22481 VSS a_12516_7093# a_46786_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22482 a_42466_65206# a_16746_65208# a_42374_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22483 a_44474_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22484 a_14912_27497# a_14287_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=150000u
X22485 a_3983_30083# a_3417_33231# a_3887_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22486 VDD a_4215_51157# a_27167_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22487 a_41370_20902# a_16362_20536# a_41462_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22488 a_5550_58255# a_4792_58371# a_4987_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22489 VDD a_6831_63303# a_30602_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2249 a_36116_50959# a_28881_52271# a_36013_50959# VSS sky130_fd_pr__nfet_01v8 ad=5.6875e+11p pd=4.35e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X22490 VSS a_12355_15055# a_36746_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22491 vcm_commonmode a_16362_8488# a_28410_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22492 a_22567_27791# a_21012_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22493 a_40762_60186# a_12981_59343# a_40366_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22494 a_40762_19898# a_12895_13967# a_40366_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22495 VSS VDD a_19678_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22496 a_28810_55488# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22497 a_23694_70226# a_12901_66665# a_23298_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22498 VSS a_12981_59343# a_49798_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22499 a_45478_56170# a_16746_56172# a_45386_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 VDD a_8177_37013# a_7244_39189# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2250 VSS a_11067_23759# a_16362_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X22500 a_46786_17890# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22501 a_34221_47695# a_33802_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22502 VDD a_3024_67191# a_9585_68841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22503 VDD VSS a_37354_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22504 vcm_commonmode a_16362_17524# a_24394_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22505 VSS a_12985_16367# a_28714_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22506 a_9624_51549# a_9187_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22507 VSS a_12907_27023# a_38115_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22508 a_26706_61190# a_12355_15055# a_26310_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22509 a_17651_30485# a_17415_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2251 a_7755_26703# a_5085_23047# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X22510 VSS a_24209_48463# a_24743_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X22511 a_1846_59475# a_2163_59585# a_2121_59709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22512 a_49494_55166# VDD a_49402_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22513 vcm_commonmode VSS a_33430_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22514 a_51330_39932# a_49750_39288# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22515 a_7901_13077# a_7999_13083# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22516 a_48398_10862# a_16362_10496# a_48490_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22517 a_38358_71230# a_12901_66665# a_38850_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22518 a_38850_20504# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22519 VDD VDD a_45386_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2252 a_49894_69544# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22520 a_38450_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22521 VSS a_32970_31145# a_32765_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22522 a_6271_72943# a_6327_72917# a_6099_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X22523 VDD a_12935_31287# a_15207_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22524 a_19703_38695# a_19919_38695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22525 a_4701_43567# a_4535_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22526 a_28410_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22527 VSS a_12899_11471# a_27710_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22528 VDD a_12546_22351# a_32334_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22529 a_31726_14878# a_12727_15529# a_31330_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2253 a_46390_66210# a_10975_66407# a_46882_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22530 a_25398_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22531 a_13543_48579# a_9989_46831# a_13461_48579# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22532 VSS a_27183_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X22533 a_13692_34191# a_13515_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22534 a_2199_31599# a_1683_31599# a_2104_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22535 a_39362_12870# a_16362_12504# a_39454_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22536 VSS a_7210_55081# a_8853_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22537 a_18370_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22538 VSS a_12901_66959# a_39758_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22539 a_36746_66210# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2254 VDD rst_n a_1591_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22540 VDD a_4503_10687# a_4490_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22541 a_32334_69222# a_12901_66959# a_32826_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22542 a_43774_67214# a_12727_67753# a_43378_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22543 vcm_commonmode a_16362_63198# a_27406_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22544 VSS a_11067_13095# a_40762_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22545 a_28318_59182# a_12901_58799# a_28810_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22546 a_16385_51183# a_16219_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22547 vcm_commonmode a_16362_20536# a_38450_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22548 a_41370_65206# a_16362_65206# a_41462_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22549 a_40967_30511# a_34759_31029# a_40861_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2255 VDD a_32970_31145# a_40691_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22550 a_19774_70548# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22551 a_33734_59182# a_12727_58255# a_33338_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22552 a_12073_71855# a_10883_71855# a_11964_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22553 a_19282_60186# a_16362_60186# a_19374_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22554 a_11613_59049# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22555 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22556 VSS a_12663_40871# a_14088_41807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22557 a_7074_15279# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22558 a_35683_50613# a_28881_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22559 a_17449_46831# a_17171_46859# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2256 a_32971_35281# a_1761_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X22560 a_29414_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22561 a_19684_37253# a_18811_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22562 VDD a_12877_14441# a_44382_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22563 a_38358_18894# a_16362_18528# a_38450_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22564 VSS a_6473_40277# a_7197_41213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X22565 VSS a_2939_31573# a_2873_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22566 a_29804_39655# a_28931_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22567 VSS a_1586_66567# a_9135_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22568 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22569 a_8105_21263# a_7757_21379# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2257 a_7090_46419# a_7368_46403# a_7324_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22570 a_2163_56765# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22571 a_9911_18870# a_9729_18870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22572 a_10097_69501# a_10053_69109# a_9931_69513# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22573 a_37750_58178# a_12901_58799# a_37354_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22574 VDD a_1915_21482# a_1867_21263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22575 a_12713_43011# a_18811_42405# a_19684_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22576 a_9215_61127# a_8500_58799# a_9560_60975# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X22577 a_2464_58077# a_2250_58077# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22578 a_2107_40303# a_1591_40303# a_2012_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22579 VSS a_12355_65103# a_17670_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2258 a_18674_55166# a_18602_55312# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X22580 a_2509_47349# a_2291_47753# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22581 VSS a_2775_46025# a_31953_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22582 a_48490_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22583 a_21479_38053# a_19780_38341# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X22584 a_45386_66210# a_16362_66210# a_45478_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22585 VSS a_7841_22895# a_10411_23759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22586 a_31726_71230# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22587 VSS a_1823_67668# a_1775_67503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22588 a_30418_69222# a_16746_69224# a_30326_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22589 a_9705_11989# a_3327_9308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2259 a_41862_9460# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22590 a_45878_11468# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22591 a_35838_68540# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22592 a_6835_31055# a_6243_30662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22593 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X22594 a_35601_27497# a_26523_28111# a_35447_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22595 a_28883_52031# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22596 a_11491_60975# a_11141_60975# a_11396_60975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22597 VDD a_12355_15055# a_17274_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22598 a_14471_28585# a_9731_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22599 a_33856_40743# a_32887_40767# a_33819_41001# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X226 a_5023_13255# a_4812_13879# a_5169_13103# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X2260 VSS a_10506_29967# a_15207_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.3585e+12p ps=1.328e+07u w=650000u l=150000u M=4
X22600 a_22386_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22601 VDD a_12985_19087# a_24302_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22602 vcm_commonmode a_16362_65206# a_31422_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22603 a_39854_67536# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22604 a_36350_64202# a_11067_13095# a_36842_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22605 a_33338_23914# a_16362_23548# a_33430_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22606 VDD a_10975_66407# a_43378_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22607 VSS a_2847_40277# a_2781_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22608 a_40858_62516# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22609 a_49402_24918# VSS a_49894_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2261 a_23390_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22610 a_12507_44310# a_12325_44310# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22611 a_1881_56623# a_1846_56875# a_1643_56597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22612 a_2463_24893# a_2315_24540# a_2100_24759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22613 a_39362_57174# a_16362_57174# a_39454_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22614 VSS a_1923_73087# a_3749_73853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22615 a_25702_62194# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22616 a_43470_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22617 a_38295_29967# a_38436_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22618 vcm_commonmode a_16362_57174# a_21382_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22619 VSS a_4571_26677# a_4351_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2262 a_49402_59182# a_16362_59182# a_49494_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22620 a_23595_41629# a_19629_39631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22621 VDD a_10515_22671# a_33338_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22622 a_2369_30333# a_2325_29941# a_2203_30345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22623 VSS a_10515_23975# a_39758_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22624 a_2012_36861# a_1761_35951# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22625 a_43870_14480# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22626 a_43774_20902# a_11067_67279# a_43378_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22627 VDD a_4719_33239# a_4191_33449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X22628 a_29147_50069# a_29561_49667# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X22629 VDD a_12257_56623# a_46390_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2263 a_4404_48829# a_4287_48634# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X22630 a_26802_24520# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22631 VSS a_12985_19087# a_36746_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22632 VDD a_3705_37557# a_3595_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22633 VDD a_11067_21583# a_30326_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22634 a_8980_71311# a_8459_71285# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X22635 VDD a_12983_63151# a_29322_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22636 a_4600_62069# a_1591_64239# a_4528_62069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22637 a_7794_53903# a_7803_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22638 a_6377_67503# a_6515_67477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22639 VSS a_23172_31573# a_23119_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X2264 VDD a_6651_31599# a_2235_30503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X22640 a_33734_12870# a_10055_58791# a_33338_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22641 a_2007_10901# a_1887_10422# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22642 a_29414_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22643 a_11143_31599# a_10870_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22644 a_46786_8854# a_12947_8725# a_46390_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22645 vcm_commonmode a_16362_23548# a_40458_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22646 VDD a_13837_38772# a_15039_38909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22647 a_16891_44265# a_15959_44031# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22648 a_21719_48285# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22649 VDD a_12727_15529# a_20286_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2265 vcm_commonmode a_16362_59182# a_31422_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22650 a_4437_10761# a_3247_10389# a_4328_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22651 a_44382_10862# a_12985_16367# a_44874_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22652 a_2834_40669# a_1757_40303# a_2672_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22653 VDD a_9215_61127# a_2794_62697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X22654 a_27314_20902# a_12985_7663# a_27806_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22655 a_10430_53181# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22656 a_42770_68218# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22657 a_27314_16886# a_16362_16520# a_27406_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22658 a_38171_34191# a_37994_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22659 a_14031_38007# a_14425_37981# a_13909_37571# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2266 a_8625_20175# a_8015_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X22660 a_33430_18528# a_16746_18526# a_33338_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X22661 VDD a_12901_58799# a_37354_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22662 a_24413_39087# a_23987_39126# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22663 a_31422_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22664 VDD a_3987_19623# a_5797_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22665 a_37750_11866# a_12985_16367# a_37354_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22666 a_7825_64239# a_2840_53511# a_7741_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22667 a_46482_17524# a_16746_17522# a_46390_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22668 VDD a_12404_34191# a_12510_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22669 a_7815_19319# a_5825_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2267 a_26889_50337# a_26671_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X22670 a_17274_12870# a_12877_16911# a_17766_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22671 VDD a_6515_67477# a_6473_67825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22672 a_21782_10464# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22673 VDD a_2847_69439# a_2834_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22674 a_30418_22544# a_16746_22542# a_30326_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22675 a_9705_11989# a_3327_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22676 a_38358_8854# a_16362_8488# a_38450_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22677 a_45782_59182# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22678 a_2215_26525# a_1591_26159# a_2107_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22679 vcm_commonmode a_16362_14512# a_34434_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2268 a_7657_64489# a_7987_64213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=7.72e+06u as=0p ps=0u w=1e+06u l=150000u
X22680 a_43378_16886# a_12899_11471# a_43870_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22681 a_28714_69222# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22682 a_7187_37583# a_6559_37583# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22683 a_31669_51433# a_2959_47113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22684 VSS a_12983_63151# a_32730_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22685 vcm_commonmode VSS a_17366_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22686 vcm_commonmode a_16362_13508# a_47486_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22687 a_5147_19605# a_4839_21495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X22688 a_7493_10749# a_7458_10515# a_7255_10357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22689 a_34434_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2269 a_40762_23914# a_10515_23975# a_40366_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X22690 a_24331_39679# a_22448_39429# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X22691 VDD a_29791_52436# a_19720_55394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22692 a_2375_49172# a_2467_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22693 VDD a_2899_27023# a_3301_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22694 a_19774_7452# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22695 VSS a_12901_58799# a_22690_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22696 a_49798_58178# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22697 a_21479_44581# a_17863_44211# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X22698 a_49798_16886# a_12727_13353# a_49402_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22699 a_20778_16488# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X227 VSS a_23993_37981# a_23685_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X2270 a_7089_29423# a_6649_25615# a_6743_29673# VSS sky130_fd_pr__nfet_01v8 ad=2.275e+11p pd=2e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X22700 a_38450_8488# a_16746_8486# a_38358_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22701 VDD VDD a_29322_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22702 VSS VDD a_25702_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22703 a_24394_13508# a_16746_13506# a_24302_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22704 vcm_commonmode a_16362_10496# a_21382_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22705 a_7113_27253# a_4427_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22706 a_37446_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22707 a_15941_31055# a_16101_31029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22708 a_23540_48981# a_23019_48463# a_23763_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22709 a_19559_34473# a_18627_34239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2271 a_40858_56492# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22710 a_49494_63198# a_16746_63200# a_49402_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22711 vcm_commonmode a_16362_60186# a_46482_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22712 vcm_commonmode a_16362_19532# a_46482_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22713 a_39176_44527# a_38999_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22714 VSS a_10515_22671# a_26706_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22715 a_23694_55166# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22716 a_36442_66210# a_16746_66212# a_36350_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22717 VSS a_11335_10076# a_11266_10205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22718 a_29322_61190# a_12981_59343# a_29814_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22719 a_35346_21906# a_16362_21540# a_35438_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2272 VDD a_18197_44220# a_17803_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X22720 a_38450_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22721 a_12787_31421# a_8461_32937# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22722 VDD a_5616_43567# a_5791_43541# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22723 VDD a_3391_15797# a_3023_16341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22724 a_12985_16367# a_12815_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X22725 a_38557_32143# a_38288_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X22726 a_5897_36611# a_3305_38671# a_5825_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22727 a_36001_31055# a_27535_30503# a_35907_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X22728 VDD a_7640_49929# a_7815_49855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22729 a_23390_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2273 a_30967_44535# a_31004_44869# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X22730 VDD a_12516_7093# a_31330_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22731 a_7197_41213# a_6927_40847# a_7107_40847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22732 a_16648_44869# a_15775_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22733 a_16843_51549# a_16219_51183# a_16735_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22734 a_77086_40693# a_76346_38962# a_76971_38925# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X22735 a_17670_71230# a_12947_71576# a_17274_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22736 a_31422_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22737 a_42770_21906# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22738 a_39362_20902# a_16362_20536# a_39454_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22739 a_45386_57174# a_12257_56623# a_45878_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2274 a_20286_24918# VSS a_20778_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22740 a_2012_26159# a_1853_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22741 VSS VDD a_40762_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22742 vcm_commonmode VSS a_41462_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22743 a_28318_67214# a_12983_63151# a_28810_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22744 a_39758_65206# a_10975_66407# a_39362_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22745 a_8395_37289# a_5915_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22746 a_32826_65528# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22747 a_3291_67325# a_3143_66972# a_2928_67191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22748 a_11136_74031# a_10055_74031# a_10789_74273# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22749 a_33430_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2275 a_2830_15431# a_2873_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22750 vcm_commonmode VSS a_17366_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22751 a_32334_55166# VSS a_32426_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22752 VSS a_12727_13353# a_48794_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22753 a_45782_12870# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22754 a_22690_24918# VSS a_22294_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22755 a_31422_71230# a_16746_71232# a_31330_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22756 a_5411_59317# a_5091_60981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X22757 a_22786_57496# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22758 a_28714_22910# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22759 vcm_commonmode a_16362_68218# a_36442_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2276 a_19789_29673# a_19442_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X22760 a_27406_7484# VDD a_27314_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22761 a_32334_14878# a_12877_14441# a_32826_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22762 VSS a_12985_7663# a_32730_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22763 a_27981_37477# a_27183_36965# a_28056_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22764 VSS a_1803_19087# a_30855_41809# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X22765 a_10391_67477# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22766 VDD a_1775_60663# a_2785_60151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22767 a_35647_41317# a_33764_41831# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X22768 a_49402_58178# a_10515_22671# a_49894_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22769 a_37354_9858# a_12546_22351# a_37846_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2277 VSS a_30155_32375# a_30105_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22770 a_28143_52105# a_27627_51733# a_28048_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22771 VDD a_5599_74549# a_6619_73719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22772 a_25702_15882# a_12877_14441# a_25306_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22773 VSS a_12877_16911# a_22690_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22774 a_5226_65693# a_4149_65327# a_5064_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22775 VSS a_12981_62313# a_34738_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22776 a_49798_11866# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22777 VDD a_3143_66972# a_7142_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22778 a_16865_27511# a_12349_25847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22779 a_47886_9460# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2278 VDD a_12516_7093# a_26310_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22780 a_25221_41281# a_24423_40229# a_25296_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22781 VSS a_12355_15055# a_47790_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22782 a_27983_40871# a_12725_44527# a_28157_40747# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22783 a_39210_48783# a_37427_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22784 a_13670_35862# a_12663_35431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X22785 vcm_commonmode a_16362_18528# a_22386_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22786 a_26802_58500# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22787 a_15017_47375# a_11067_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22788 VDD a_5975_71829# a_5962_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22789 a_7159_50260# a_7251_50069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2279 VDD a_32227_48169# a_33515_48576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X22790 VSS a_10055_58791# a_26706_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22791 a_4761_65327# a_4717_65569# a_4595_65327# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X22792 a_8263_45908# a_8308_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22793 a_24698_62194# a_12981_62313# a_24302_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22794 a_12714_30761# a_2787_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X22795 a_2713_31353# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22796 VSS a_11067_13095# a_38754_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22797 VDD a_12707_26159# a_13919_27904# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22798 a_36350_72234# VDD a_36842_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22799 a_36842_21508# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X228 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u M=254
X2280 VDD a_12985_19087# a_27314_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X22800 a_40858_70548# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22801 a_36442_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22802 a_2163_73085# a_1586_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22803 a_39362_65206# a_16362_65206# a_39454_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22804 a_2475_68425# a_2125_68053# a_2380_68413# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22805 a_43470_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22806 a_40366_60186# a_16362_60186# a_40458_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22807 a_49894_20504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22808 VDD a_1950_59887# a_3983_68591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22809 a_49494_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2281 VDD a_5331_18517# a_4792_20443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X22810 a_23298_70226# a_16362_70226# a_23390_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22811 a_7622_57711# a_7580_61751# a_7812_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22812 a_5261_59343# a_5190_59575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X22813 a_4607_48463# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22814 VSS a_1586_9991# a_1591_12565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22815 VSS a_7580_61751# a_8152_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22816 a_39854_12472# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22817 a_25419_50959# a_28671_30539# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X22818 a_11696_26409# a_10286_26311# a_11612_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22819 a_37354_13874# a_16362_13508# a_37446_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2282 VDD a_19096_44129# a_18197_44220# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X22820 VDD a_12546_22351# a_43378_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22821 a_6516_53511# a_6666_53359# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22822 a_7390_32693# a_6883_37019# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22823 VDD a_11067_67279# a_26310_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22824 a_41766_68218# a_12901_66959# a_41370_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22825 a_4127_63669# a_4330_63827# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22826 VDD a_12263_4391# a_12815_4399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22827 a_12985_25615# a_12394_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22828 a_29414_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22829 a_26310_61190# a_16362_61190# a_26402_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2283 a_7519_59575# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22830 VSS a_12935_31287# a_15207_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22831 VDD a_1761_25615# a_1959_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X22832 vcm_commonmode a_16362_56170# a_42466_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22833 a_39454_24552# VDD a_39362_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22834 a_35337_52093# a_29361_51727# a_35237_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22835 vcm_commonmode a_16362_21540# a_36442_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22836 a_29718_71230# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22837 VDD a_1586_69367# a_1591_69141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22838 a_28410_69222# a_16746_69224# a_28318_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22839 vcm_commonmode a_16362_66210# a_25398_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2284 a_22438_49007# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X22840 VSS a_19807_28111# a_33635_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22841 VDD a_1923_59583# a_3667_60405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22842 a_27314_24918# VSS a_27406_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22843 VDD a_12983_63151# a_37354_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22844 VDD a_17763_35797# a_17585_37477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X22845 a_34834_63520# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22846 a_31422_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22847 a_44778_59182# a_12727_58255# a_44382_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22848 a_27406_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22849 VSS a_8123_56399# a_8219_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2285 a_26402_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22850 VDD a_9314_69367# a_10055_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22851 VSS a_12981_59343# a_23694_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22852 a_20682_17890# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22853 a_32135_49007# a_28108_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22854 a_10648_28995# a_7841_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22855 vcm_commonmode a_16362_65206# a_29414_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22856 a_2834_12559# a_1757_12565# a_2672_12937# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22857 a_30326_9858# a_16362_9492# a_30418_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22858 a_38850_62516# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22859 a_48794_7850# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 a_23298_56170# a_16362_56170# a_23390_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X22860 a_48794_58178# a_12901_58799# a_48398_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22861 VSS a_14646_29423# a_23172_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22862 a_43378_67214# a_16362_67214# a_43470_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22863 VDD a_12981_59343# a_42374_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22864 VSS VSS a_45782_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22865 a_9379_15039# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22866 VSS a_5428_63669# a_5366_63695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22867 a_12126_18909# a_11049_18543# a_11964_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22868 a_27234_29789# a_5363_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22869 vcm_commonmode a_16362_57174# a_19374_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2287 a_3316_42313# a_2235_41941# a_2969_41909# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X22870 a_23390_55166# VDD a_23298_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22871 a_24698_16886# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22872 VDD config_1_in[11] a_1626_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22873 a_7097_67655# a_5254_67503# a_7260_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22874 a_22294_10862# a_16362_10496# a_22386_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22875 a_16928_35303# a_15959_35327# a_16832_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22876 a_1761_46287# a_1591_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22877 a_20378_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22878 a_1757_71317# a_1591_71317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22879 VDD a_7203_10383# a_9219_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2288 a_37750_21906# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X22880 VDD a_12355_15055# a_28318_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22881 VSS a_2292_17179# a_2369_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22882 a_1895_38842# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22883 a_5064_20719# a_3983_20719# a_4717_20961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22884 a_15305_38543# a_15039_38909# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X22885 VDD a_12895_13967# a_19282_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22886 a_37354_58178# a_16362_58178# a_37446_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22887 a_5553_63401# a_5497_63303# a_2944_64488# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22888 a_41211_28023# a_11067_46823# a_41385_28129# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X22889 a_31004_44869# a_30035_44581# a_30908_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2289 vcm_commonmode a_16362_71230# a_49494_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22890 a_23694_63198# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22891 a_3980_35523# a_1915_35015# a_3885_35523# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22892 a_35742_7850# VDD a_35346_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22893 VDD a_16101_31029# a_18053_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22894 VSS a_33656_43439# a_33762_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22895 a_19541_29423# a_18829_29423# a_19459_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22896 a_37354_17890# a_12899_10927# a_37846_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22897 VSS a_12947_23413# a_37750_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22898 VDD a_2235_30503# a_23731_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22899 a_4075_14191# a_3023_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X229 a_1761_22895# a_1591_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2290 a_4495_35925# a_5405_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X22900 VSS a_12546_22351# a_40762_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22901 a_17711_40183# a_18105_40157# a_13576_40413# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X22902 VSS a_12659_54965# a_12785_53181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22903 a_41862_15484# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22904 a_41766_21906# a_12985_7663# a_41370_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22905 a_18811_41317# a_18045_41281# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X22906 a_7571_72512# a_6453_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22907 a_30722_66210# a_12983_63151# a_30326_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22908 VDD a_10515_22671# a_44382_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22909 a_10045_14013# a_7841_12167# a_9963_13760# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2291 a_22062_31287# a_20881_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22910 a_21290_22910# a_10515_23975# a_21782_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22911 VSS a_35615_30199# a_33839_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X22912 a_28410_22544# a_16746_22542# a_28318_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22913 vcm_commonmode a_16362_70226# a_37446_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22914 a_18022_49007# a_17039_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22915 VDD a_1586_40455# a_4535_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22916 a_27406_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22917 a_26706_9858# a_12985_19087# a_26310_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22918 a_44778_12870# a_10055_58791# a_44382_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22919 VDD a_3417_33231# a_3983_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2292 a_35739_39679# a_34699_38771# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X22920 a_42374_11866# a_10055_58791# a_42866_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22921 a_27710_64202# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22922 a_2672_18543# a_1757_18543# a_2325_18785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22923 a_25306_21906# a_11067_21583# a_25798_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22924 VDD a_3421_57167# a_3521_57283# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22925 a_25306_17890# a_16362_17524# a_25398_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22926 VDD a_12727_15529# a_31330_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22927 a_37446_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22928 VDD a_12727_58255# a_35346_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22929 a_9123_55223# a_9695_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2293 a_10835_52271# a_10687_52553# a_10472_52423# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X22930 a_32334_63198# a_16362_63198# a_32426_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22931 a_17670_56170# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22932 VDD a_12901_58799# a_48398_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22933 vcm_commonmode a_16362_15516# a_41462_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22934 a_44474_18528# a_16746_18526# a_44382_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22935 a_18770_16488# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22936 a_5483_11140# a_5601_11471# a_5645_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22937 a_48794_11866# a_12985_16367# a_48398_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22938 a_2215_19997# a_1591_19631# a_2107_19631# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22939 vcm_commonmode a_16362_10496# a_19374_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2294 VDD a_12815_16519# a_12815_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X22940 a_12549_44212# a_12671_43222# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22941 a_28318_12870# a_12877_16911# a_28810_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22942 a_32826_10464# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22943 a_49402_66210# a_10975_66407# a_49894_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22944 a_17366_61190# a_16746_61192# a_17274_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22945 a_7987_15431# a_2004_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22946 a_22062_31287# a_20905_32143# a_22365_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22947 a_18501_50645# a_18335_50645# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X22948 VSS a_12727_67753# a_30722_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22949 a_4220_57685# a_4674_57685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2295 a_27337_38565# a_26447_39141# a_27379_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X22950 a_11763_57399# a_11883_58575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22951 a_2375_13268# a_2313_12015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X22952 VSS a_2835_62215# a_2787_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22953 vcm_commonmode a_16362_14512# a_45478_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22954 a_10317_13647# a_9963_13760# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22955 a_7436_46983# a_6835_46823# a_7578_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22956 a_41370_19898# a_11067_67279# a_41862_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22957 vcm_commonmode VSS a_28410_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22958 a_42466_9492# a_16746_9490# a_42374_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22959 a_12010_28111# a_8935_27791# a_11711_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2296 a_16928_42919# a_15959_42943# a_16832_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X22960 VDD a_17939_43745# a_17763_43413# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22961 a_12800_43983# a_12549_44212# a_12579_44310# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22962 a_43870_56492# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22963 a_2250_73309# a_2124_73211# a_1846_73195# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X22964 a_7439_64213# a_7567_64391# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22965 a_45478_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22966 VDD a_11136_74031# a_11311_74005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22967 VDD a_2764_31599# a_2939_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22968 a_26802_66532# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22969 a_18370_9492# a_16746_9490# a_18278_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2297 VDD a_4711_54965# a_4642_54991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X22970 a_23298_63198# a_12981_62313# a_23790_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22971 a_13353_30511# a_12786_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X22972 vcm_commonmode a_16362_16520# a_18370_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22973 VDD a_12355_65103# a_30326_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22974 a_22386_14512# a_16746_14510# a_22294_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22975 a_4529_40553# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22976 a_35438_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22977 VSS a_1761_4399# a_1683_5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22978 VDD a_26495_35253# a_26319_35253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22979 VSS a_38044_44759# a_37857_44501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2298 a_44874_55488# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22980 a_22319_38825# a_21387_38591# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22981 VSS config_2_in[5] a_1591_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X22982 VSS a_7019_30511# a_7116_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22983 VDD a_12257_56623# a_20286_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22984 VSS VDD a_38754_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22985 VDD a_6098_73095# a_7571_72512# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22986 a_34434_67214# a_16746_67216# a_34342_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22987 a_42770_70226# a_12901_66665# a_42374_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22988 VDD a_7005_55223# a_6138_54599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X22989 VSS a_24331_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X2299 VSS VDD a_35742_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22990 a_10949_72719# a_10509_73193# a_10865_72719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22991 a_27314_62194# a_12355_15055# a_27806_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22992 a_31822_60508# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22993 a_47486_66210# a_16746_66212# a_47394_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22994 VSS a_19127_43439# a_19233_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X22995 a_49494_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22996 a_2957_72105# a_2843_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22997 a_46390_21906# a_16362_21540# a_46482_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X22998 a_32730_62194# a_12981_62313# a_32334_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22999 a_2345_33749# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23 a_12161_31599# a_11143_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X230 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2300 a_24302_23914# a_12947_23413# a_24794_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23000 a_45782_61190# a_12355_15055# a_45386_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23001 a_2121_57711# a_1643_57685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23002 VSS a_12899_10927# a_42770_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23003 a_24331_38591# a_23565_38565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X23004 a_2250_58077# a_2163_57853# a_1846_57963# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23005 a_28714_71230# a_12947_71576# a_28318_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23006 vcm_commonmode a_16362_8488# a_21382_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23007 VDD a_5993_32687# a_7545_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23008 VDD a_30125_47919# a_30479_48576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23009 a_19877_41972# a_19967_41781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2301 VDD a_2325_66657# a_2215_66781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X23010 VSS a_12899_11471# a_46786_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23011 a_43774_13874# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23012 a_44474_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23013 a_20195_49793# a_4191_33449# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23014 a_8639_15113# a_8123_14741# a_8544_15101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23015 a_34834_71552# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23016 a_26706_23914# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23017 VDD a_4248_29967# a_8493_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23018 a_30326_15882# a_12727_13353# a_30818_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23019 VSS a_11067_21583# a_30722_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2302 VDD a_30835_39783# a_14963_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X23020 VSS a_1803_19087# a_1945_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23021 a_27406_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23022 a_2882_58077# a_2163_57853# a_2319_57948# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23023 a_34342_61190# a_16362_61190# a_34434_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23024 VDD a_4075_64239# a_4167_64783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23025 VSS a_4495_35925# a_4443_36611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23026 a_38292_30511# a_34759_31029# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23027 a_17274_71230# a_16362_71230# a_17366_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23028 VDD a_37888_34191# a_37994_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23029 a_47394_59182# a_12901_58799# a_47886_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2303 a_24302_19898# a_16362_19532# a_24394_19532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23030 VSS a_12895_13967# a_19678_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23031 a_13867_42134# a_12889_40977# a_13795_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X23032 a_17103_49007# a_16587_49007# a_17008_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23033 a_31611_43447# a_30679_43493# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23034 a_23694_16886# a_12727_13353# a_23298_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23035 VSS a_12727_15529# a_20682_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23036 a_13528_36055# a_13743_35836# a_13670_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23037 a_18627_42943# a_17711_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X23038 a_38850_70548# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23039 a_4734_63695# a_4647_63937# a_4330_63827# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2304 a_27806_65528# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23040 VSS a_12981_62313# a_45782_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23041 a_3005_56079# a_2727_56417# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X23042 a_35742_69222# a_12516_7093# a_35346_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23043 a_16257_38517# a_12663_39783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23044 VDD a_2503_34319# a_3217_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23045 a_19578_50639# a_18501_50645# a_19416_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23046 a_23390_63198# a_16746_63200# a_23298_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23047 vcm_commonmode a_16362_60186# a_20378_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23048 VDD a_11521_66567# a_12066_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23049 a_10995_14333# a_1586_18695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2305 VDD a_33515_30511# a_33694_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X23050 a_13669_37429# a_31083_36395# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X23051 a_2040_43401# a_1757_43029# a_1945_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23052 a_48490_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23053 vcm_commonmode a_16362_19532# a_20378_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23054 VDD a_29915_41959# a_18127_35797# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X23055 a_24794_59504# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23056 a_30609_49159# a_30479_48576# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23057 a_12227_51017# a_11877_50645# a_12132_51005# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23058 a_2325_26401# a_2107_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23059 a_10288_53047# a_6559_59663# a_10430_53181# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X2306 a_1761_32143# a_1591_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23060 a_34434_20536# a_16746_20534# a_34342_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23061 vcm_commonmode a_16362_18528# a_33430_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23062 VSS a_7255_10357# a_7203_10383# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23063 a_32795_38591# a_32029_38565# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23064 VSS a_18627_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23065 VSS a_6559_22671# a_7431_22441# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23066 VSS a_17843_48981# a_17777_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23067 a_26447_35279# a_12549_35836# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23068 a_11709_65569# a_11491_65327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23069 VSS a_12355_65103# a_36746_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2307 VSS a_19675_49525# a_14985_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23070 a_35739_39679# a_34699_38771# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23071 VDD a_12899_11471# a_36350_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23072 a_39758_9858# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23073 a_32672_49007# a_32135_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X23074 VSS a_41443_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23075 a_34434_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23076 VDD a_13620_40871# a_12641_42036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23077 a_9370_69831# a_9466_69653# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23078 VSS a_11067_13095# a_49798_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23079 VSS a_1586_18695# a_1591_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2308 a_18672_38567# a_18045_39105# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X23080 a_47886_21508# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23081 a_47486_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23082 VSS a_12546_22351# a_49798_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23083 VDD a_22351_47893# a_22338_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23084 a_2325_14709# a_2107_15113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23085 a_8168_53359# a_8132_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23086 VDD a_11155_30663# a_11183_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23087 VSS a_12947_56817# a_39758_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23088 VSS a_4719_51183# a_4215_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X23089 a_32334_56170# a_12947_56817# a_32826_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2309 a_43470_61190# a_16746_61192# a_43378_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23090 a_41462_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23091 a_37846_13476# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23092 VDD a_12985_16367# a_41370_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23093 a_26706_64202# a_12355_65103# a_26310_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23094 a_23784_42583# a_23880_42325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23095 a_11372_30511# a_10899_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23096 VDD a_12985_7663# a_24302_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23097 a_48398_13874# a_16362_13508# a_48490_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23098 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23099 a_27406_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X231 a_32334_7850# VSS a_32426_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2310 a_27314_55166# VSS a_27406_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23100 a_12191_39095# a_12585_39069# a_12251_39069# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X23101 a_44778_62194# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23102 vcm_commonmode a_16362_57174# a_40458_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23103 a_8541_44449# a_8475_44343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23104 a_2325_69109# a_2107_69513# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23105 a_24423_40229# a_23415_41263# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X23106 a_27710_72234# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23107 VDD a_7387_46831# a_7387_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23108 vcm_commonmode a_16362_67214# a_23390_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23109 a_31898_30761# a_19807_28111# a_31741_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2311 vcm_commonmode a_16362_17524# a_40458_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23110 a_15812_31029# a_14625_30761# a_15941_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X23111 VSS a_12516_7093# a_31726_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23112 VSS a_7155_55509# a_7101_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23113 VDD a_12727_67753# a_35346_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23114 a_2203_36873# a_1757_36501# a_2107_36873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23115 a_6451_22895# a_6007_23145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X23116 a_13835_43177# a_27183_43493# a_28115_43447# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X23117 a_46390_8854# a_12985_19087# a_46882_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23118 a_25398_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23119 a_5393_69455# a_5213_70223# a_5484_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2312 a_2369_44655# a_2325_44897# a_2203_44655# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X23120 VDD a_12983_63151# a_48398_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23121 a_45878_63520# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23122 VSS a_12355_15055# a_21686_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23123 a_28305_28879# a_28027_29217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X23124 a_7553_62927# a_7523_62581# a_7457_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23125 a_18370_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23126 a_1757_21807# a_1591_21807# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23127 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23128 a_3040_68425# a_1959_68053# a_2693_68021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23129 a_48490_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2313 a_17670_24918# VSS a_17274_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23130 a_35742_22910# a_11067_21583# a_35346_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23131 a_30418_56170# a_16746_56172# a_30326_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23132 a_31726_17890# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23133 a_16257_38517# a_12663_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23134 VSS a_13669_39605# a_13613_39958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23135 a_28714_8854# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23136 a_41370_68218# a_16362_68218# a_41462_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23137 VDD VSS a_22294_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23138 a_5437_11791# a_4812_13879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23139 a_3118_52271# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2314 a_39409_28585# a_38210_30199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X23140 a_7203_71017# a_6224_73095# a_7457_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X23141 vcm_commonmode a_16362_58178# a_17366_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23142 a_49894_62516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23143 a_28172_31415# a_27797_29423# a_28089_31157# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23144 a_2325_49525# a_2107_49929# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23145 a_2873_33609# a_1683_33237# a_2764_33609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23146 a_28909_49871# a_27869_50095# a_28691_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23147 VDD a_9914_68279# a_9865_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23148 VDD a_12056_60975# a_12231_60949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23149 VSS a_15345_34717# a_15037_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2315 a_4515_50639# a_3891_50645# a_4407_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X23150 VDD a_21712_43781# a_21049_41245# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X23151 VDD a_28757_27247# a_41795_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23152 a_2813_56417# a_1591_56623# a_2727_56417# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X23153 a_12605_54991# a_12755_53030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23154 VDD a_30991_29397# a_27752_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23155 VDD a_12947_8725# a_33338_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23156 a_33338_10862# a_16362_10496# a_33430_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23157 a_19282_22910# a_10515_23975# a_19774_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23158 a_23298_71230# a_12901_66665# a_23790_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23159 a_23790_20504# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2316 a_26402_71230# a_16746_71232# a_26310_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23160 VDD VDD a_30326_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23161 a_23390_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23162 a_6821_26311# a_5211_24759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23163 VDD a_12981_62313# a_26310_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23164 VDD a_7072_56053# a_6072_56872# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23165 a_47790_69222# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23166 a_36904_28879# a_36425_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X23167 VDD a_2805_22869# a_2835_23222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23168 VSS a_5959_13621# a_5903_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23169 a_5755_14709# a_6895_15253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2317 a_47790_13874# a_12877_16911# a_47394_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23170 vcm_commonmode a_16362_23548# a_49494_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23171 a_21873_47919# a_21829_48161# a_21707_47919# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23172 a_31822_8456# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23173 a_27314_70226# a_12516_7093# a_27806_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23174 a_48398_58178# a_16362_58178# a_48490_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23175 a_18811_34789# a_16928_36391# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23176 VSS a_32327_35839# a_32273_36161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23177 VSS a_12901_58799# a_41766_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23178 a_35346_18894# a_12895_13967# a_35838_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23179 VSS VSS a_35742_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2318 VSS a_12985_16367# a_44778_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23180 a_2788_43389# a_1591_43029# a_2592_43023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23181 a_24302_12870# a_16362_12504# a_24394_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23182 a_34895_30511# a_34759_31029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23183 a_11893_66191# a_11619_63151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23184 a_33764_38567# a_32795_38591# a_33668_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23185 VDD a_2672_51183# a_2847_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23186 VSS a_12901_66959# a_24698_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23187 a_21686_66210# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23188 vcm_commonmode a_16362_15516# a_39454_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23189 a_48398_17890# a_12899_10927# a_48890_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2319 a_17766_57496# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23190 a_43470_13508# a_16746_13506# a_43378_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23191 vcm_commonmode a_16362_10496# a_40458_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23192 a_12549_35836# a_13867_35606# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23193 VSS a_1770_14441# a_1824_61127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23194 vcm_commonmode a_16362_20536# a_23390_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23195 a_26402_23548# a_16746_23546# a_26310_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23196 a_39454_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23197 a_25398_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23198 VSS a_2606_41079# a_7889_48246# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23199 a_42770_55166# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X232 VSS a_13445_50639# a_15211_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X2320 VDD a_13576_40413# a_12677_40157# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X23200 a_10701_31849# a_8273_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23201 vcm_commonmode a_16362_70226# a_48490_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23202 VSS a_12727_67753# a_28714_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23203 a_25702_65206# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23204 a_25798_17492# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23205 a_23298_18894# a_16362_18528# a_23390_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23206 a_17366_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23207 a_39362_19898# a_11067_67279# a_39854_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23208 a_1643_63125# a_1846_63403# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23209 a_43378_68218# a_12727_67753# a_43870_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2321 a_24194_35823# a_24017_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23210 vcm_commonmode a_16362_62194# a_38450_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23211 VSS a_5871_47594# a_4240_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X23212 a_42466_60186# a_16746_60188# a_42374_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23213 a_42466_19532# a_16746_19530# a_42374_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23214 VDD a_12727_58255# a_46390_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23215 VSS a_2695_58951# a_2695_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X23216 a_9405_10927# a_9414_10383# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23217 a_22690_58178# a_12901_58799# a_22294_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23218 a_25263_29981# a_25368_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23219 a_33760_42693# a_32887_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2322 VDD VSS a_21290_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X23220 a_25398_70226# a_16746_70228# a_25306_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23221 a_28714_56170# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23222 a_30326_66210# a_16362_66210# a_30418_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23223 vcm_commonmode a_16362_11500# a_17366_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23224 a_29814_16488# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23225 a_26310_13874# a_12727_15529# a_26802_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23226 a_1895_38842# a_2927_39733# a_2885_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23227 a_18844_43439# a_18667_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23228 a_30818_11468# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23229 a_20778_68540# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2323 a_27314_14878# a_12877_14441# a_27806_14480# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23230 VDD a_6625_29941# a_6039_30663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X23231 a_47394_67214# a_12983_63151# a_47886_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23232 VDD a_2375_48084# a_2079_47546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23233 a_11699_58799# a_11521_66567# a_11115_59317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23234 a_1761_35407# a_1591_35407# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23235 a_4241_18543# a_4075_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23236 a_39305_48169# a_37557_32463# a_39222_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23237 a_7079_52815# a_7217_53047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23238 a_19678_14878# a_12727_15529# a_19282_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23239 a_1644_54965# a_1823_54973# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2324 VSS a_12985_7663# a_27710_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23240 a_1925_18231# a_2021_17973# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23241 VDD config_1_in[6] a_1591_2767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23242 a_34738_23914# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23243 VDD a_2473_34293# a_4055_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23244 a_33826_50075# a_33515_48576# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23245 a_26576_50095# a_6559_59663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23246 a_41862_57496# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23247 a_47790_22910# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23248 a_10382_58487# a_10478_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23249 a_24794_67536# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2325 VSS a_14354_32117# a_15162_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X23250 a_21290_64202# a_11067_13095# a_21782_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23251 a_18835_48502# a_18653_48502# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23252 a_13565_44135# a_13661_43957# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23253 a_32402_48463# a_32318_48695# a_32319_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23254 a_24302_57174# a_16362_57174# a_24394_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23255 a_19611_28335# a_11902_27497# a_19442_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23256 VSS a_12877_16911# a_41766_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23257 VDD a_5239_48767# a_5226_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23258 a_2375_76372# a_2361_74575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23259 VSS a_10515_23975# a_24698_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 a_31822_12472# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23260 a_37423_51335# a_37512_50755# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X23261 VDD a_12257_56623# a_31330_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23262 a_45478_67214# a_16746_67216# a_45386_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23263 VDD a_25971_29967# a_25971_29789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X23264 a_17670_17890# a_12899_11471# a_17274_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23265 a_20378_7484# VDD a_20286_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23266 a_35647_39141# a_33764_38567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X23267 a_36746_61190# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23268 VSS a_11067_21583# a_28714_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23269 a_35438_59182# a_16746_59184# a_35346_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2327 a_25306_9858# a_16362_9492# a_25398_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23270 a_43774_62194# a_12981_62313# a_43378_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23271 VSS a_12895_13967# a_40762_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23272 a_26706_72234# VDD a_26310_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23273 a_1915_11092# a_2007_10901# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23274 VDD a_12901_58799# a_22294_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23275 VSS a_8958_65961# a_8753_66103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23276 VSS a_12727_15529# a_18674_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23277 a_22690_11866# a_12985_16367# a_22294_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23278 a_40858_9460# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23279 a_31422_17524# a_16746_17522# a_31330_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2328 VSS a_22015_28111# a_35132_47695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23280 VSS a_28757_27247# a_35687_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23281 a_39454_58178# a_16746_58180# a_39362_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23282 vcm_commonmode VSS a_36442_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23283 a_42374_70226# a_16362_70226# a_42466_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23284 a_41766_14878# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23285 a_30722_59182# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23286 VDD a_12985_7663# a_32334_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23287 a_9832_60797# a_9424_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23288 a_5381_68345# a_2843_71829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23289 VDD a_12985_19087# a_26310_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2329 a_36613_48169# a_21187_29415# a_36541_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X23290 VSS a_2419_48783# a_12489_51005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23291 VSS a_18351_37503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23292 a_38013_47919# a_13643_28327# a_21371_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23293 a_45878_71552# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23294 VDD a_11067_67279# a_45386_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23295 VSS a_1923_54591# a_2461_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23296 vcm_commonmode a_16362_13508# a_32426_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23297 VSS a_12727_58255# a_17670_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23298 VSS a_4036_54421# a_3295_54421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X23299 VDD a_10317_55223# a_9695_54965# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X233 VSS a_12447_29199# a_38210_30199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X2330 VSS a_4351_67279# a_37459_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X23300 VSS a_11067_67279# a_17670_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23301 a_48490_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23302 a_45386_61190# a_16362_61190# a_45478_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23303 VDD a_2292_17179# a_3391_15797# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23304 VSS a_43678_31029# a_43319_31029# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23305 a_28318_71230# a_16362_71230# a_28410_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23306 vcm_commonmode a_16362_66210# a_44474_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23307 VDD a_10055_58791# a_35346_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23308 a_33430_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23309 VSS config_2_in[12] a_1591_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2331 VDD a_5105_47673# a_5135_47414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X23310 a_35463_44031# a_33856_44869# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23311 VDD a_11067_21583# a_18278_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23312 a_49894_70548# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23313 a_5502_33053# a_4425_32687# a_5340_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23314 a_46482_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23315 a_12166_21501# a_5535_18012# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X23316 a_30415_43177# a_29483_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23317 VDD a_12381_35836# a_12325_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X23318 a_22386_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23319 a_46786_69222# a_12516_7093# a_46390_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2332 vcm_commonmode a_16362_16520# a_44474_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23320 a_49402_60186# a_16362_60186# a_49494_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23321 VSS a_12985_19087# a_38754_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23322 a_11495_16341# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23323 a_11771_68021# a_11947_68279# a_12157_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X23324 vcm_commonmode a_16362_60186# a_31422_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23325 vcm_commonmode a_16362_19532# a_31422_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23326 a_21382_66210# a_16746_66212# a_21290_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23327 a_1915_45908# a_2007_45717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23328 a_48794_8854# a_12947_8725# a_48398_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23329 a_24184_47741# a_7479_54439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X2333 VSS a_12877_16911# a_17670_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23330 a_45478_20536# a_16746_20534# a_45386_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23331 a_23390_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23332 VDD a_13445_50639# a_16902_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23333 a_20286_21906# a_16362_21540# a_20378_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23334 a_7037_19385# a_3247_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23335 VDD a_12901_66665# a_26310_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23336 a_19374_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23337 a_15661_29967# a_15799_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23338 VDD a_12899_10927# a_34342_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23339 VSS a_2216_28309# a_4177_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2334 VDD a_7623_13621# a_6738_19783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23340 a_1916_33927# a_2011_34837# a_2058_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23341 VDD a_3040_68425# a_3215_68351# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23342 a_33597_50141# a_30928_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23343 a_26402_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23344 VDD a_9529_28335# a_15146_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23345 VSS a_12355_65103# a_47790_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23346 a_5173_48841# a_3983_48469# a_5064_48841# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23347 a_6154_71855# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23348 a_2497_53903# a_2327_53903# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23349 a_35438_12504# a_16746_12502# a_35346_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2335 a_21686_10862# a_12546_22351# a_21290_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23350 a_45478_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23351 a_13097_35279# a_12831_35645# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23352 VSS a_36324_34191# a_36430_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23353 a_25493_29967# a_25145_30083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X23354 a_2746_16885# a_2596_16911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X23355 a_24302_20902# a_16362_20536# a_24394_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23356 a_35346_69222# a_16362_69222# a_35438_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23357 VSS a_12257_56623# a_37750_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23358 a_30326_57174# a_12257_56623# a_30818_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23359 a_41766_55166# VSS a_41370_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2336 VDD a_51330_39932# a_51936_39932# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u M=2
X23360 a_5366_63695# a_4608_63811# a_4803_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23361 a_35346_7850# VDD a_35838_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23362 a_24698_65206# a_10975_66407# a_24302_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23363 VDD a_12355_15055# a_47394_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23364 a_14081_42134# a_13909_41923# a_13867_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X23365 a_14577_27247# a_11430_26159# a_14287_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23366 a_39454_11500# a_16746_11498# a_39362_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23367 VDD a_77568_39738# a_77381_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23368 a_13670_36189# a_12663_35431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23369 a_28410_56170# a_16746_56172# a_28318_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2337 a_21479_44581# a_17863_44211# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23370 a_29718_17890# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23371 VDD a_12895_13967# a_38358_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23372 a_45878_7452# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23373 a_41766_7850# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23374 a_30722_12870# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23375 a_42770_63198# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23376 VSS a_17358_31069# a_17187_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23377 a_39362_68218# a_16362_68218# a_39454_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23378 a_32406_47919# a_6831_63303# a_32227_48169# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u w=650000u l=150000u
X23379 VDD a_2672_23817# a_2847_23743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2338 a_6194_30511# a_2787_32679# a_5915_30511# VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=3.9975e+11p ps=3.83e+06u w=650000u l=150000u
X23380 vcm_commonmode a_16362_68218# a_21382_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23381 a_16744_40517# a_15775_40229# a_16648_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23382 a_17670_7850# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23383 a_13867_35279# a_13613_35606# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23384 a_4549_58621# a_4514_58387# a_4311_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23385 VDD a_10531_31055# a_14625_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X23386 VSS a_14963_39783# a_19424_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23387 VDD a_4215_51157# a_24683_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23388 a_40366_22910# a_10515_23975# a_40858_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23389 VSS a_6743_23555# a_7187_23439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X2339 a_31422_24552# VDD a_31330_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23390 VSS VDD a_27710_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23391 a_12953_53339# a_12631_52928# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23392 a_33430_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23393 VDD a_12727_67753# a_46390_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23394 a_7340_65693# a_7126_65693# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23395 a_30311_35877# a_29545_35841# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23396 a_23172_31573# a_23626_31573# a_23564_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X23397 a_29498_31171# a_8491_41383# a_29416_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23398 a_46482_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23399 a_4067_15797# a_3872_15939# a_4377_16189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X234 a_28410_52637# a_27333_52271# a_28248_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2340 VDD a_20957_36604# a_20563_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X23400 a_10651_53181# a_10503_52828# a_10288_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23401 a_5249_56623# a_4771_56597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23402 a_33830_17492# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23403 a_33734_23914# a_10515_23975# a_33338_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23404 VSS a_12355_15055# a_32730_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23405 a_29414_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23406 VSS a_36904_28879# a_37919_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23407 VSS a_2451_72373# a_1895_71482# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X23408 a_46786_22910# a_11067_21583# a_46390_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23409 a_12901_52521# a_12659_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2341 VSS a_39272_31573# a_32970_31145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X23410 VDD a_12516_7093# a_19282_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23411 a_44382_21906# a_11067_21583# a_44874_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23412 a_44382_17890# a_16362_17524# a_44474_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23413 a_18811_39141# a_18045_39105# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X23414 VDD a_28757_27247# a_35458_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23415 VDD a_32227_48169# a_33681_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23416 a_19374_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23417 VDD a_21948_34973# a_21049_34717# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X23418 a_33430_70226# a_16746_70228# a_33338_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X23419 a_26495_42869# a_12381_43957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2342 a_15095_41781# a_15193_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23420 vcm_commonmode a_16362_58178# a_28410_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23421 VDD a_4127_50069# a_4031_50247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X23422 a_34342_13874# a_12727_15529# a_34834_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23423 a_19678_66210# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23424 VSS a_11067_13095# a_23694_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23425 a_37846_55488# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23426 a_17274_23914# a_12947_23413# a_17766_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23427 a_21290_72234# VDD a_21782_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23428 a_17274_19898# a_16362_19532# a_17366_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23429 a_47394_12870# a_12877_16911# a_47886_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2343 a_44474_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23430 a_21782_21508# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23431 VDD VDD a_30326_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23432 a_21382_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23433 VDD a_6895_15253# a_6882_15645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23434 VSS a_52778_39198# a_7841_12167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23435 a_24302_65206# a_16362_65206# a_24394_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23436 a_36442_61190# a_16746_61192# a_36350_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23437 VDD a_76346_38962# a_77451_38925# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X23438 vcm_commonmode VSS a_43470_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23439 a_3112_9527# a_3327_9308# a_3254_9334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X2344 a_46786_60186# a_12981_59343# a_46390_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23440 a_19374_71230# a_16746_71232# a_19282_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23441 a_8263_45908# a_8308_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23442 VSS a_12985_16367# a_37750_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23443 a_1757_21807# a_1591_21807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23444 a_3026_45565# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23445 vcm_commonmode VSS a_19374_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23446 vcm_commonmode VSS a_47486_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23447 VDD a_12877_14441# a_27314_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23448 a_24794_12472# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23449 a_22294_13874# a_16362_13508# a_22386_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2345 a_46786_19898# a_12895_13967# a_46390_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23450 VSS a_20743_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23451 a_42374_63198# a_12981_62313# a_42866_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23452 a_29414_7484# VDD a_29322_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23453 vcm_commonmode a_16362_16520# a_37446_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23454 a_46390_18894# a_12895_13967# a_46882_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23455 a_41462_14512# a_16746_14510# a_41370_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23456 a_39362_9858# a_12546_22351# a_39854_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23457 a_24394_24552# VDD a_24302_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23458 a_34267_31599# a_34016_31849# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X23459 vcm_commonmode a_16362_21540# a_21382_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2346 VSS a_4842_45467# a_6169_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X23460 a_9275_15253# a_9379_15039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23461 a_29391_44031# a_28152_44869# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23462 a_37446_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23463 a_39758_60186# a_12981_59343# a_39362_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23464 a_28810_11468# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23465 a_39758_19898# a_12895_13967# a_39362_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23466 VDD a_5136_34551# a_5079_35639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X23467 a_18770_68540# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23468 VSS a_15069_35805# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23469 a_9204_30663# a_8733_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X2347 a_40895_36919# a_25133_37571# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X23470 a_49894_9460# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23471 VDD a_12983_63151# a_22294_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23472 a_16043_38825# a_15683_39141# a_16615_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X23473 VSS a_3355_25071# a_4351_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23474 a_1643_56597# a_1846_56875# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23475 a_24029_39355# a_35647_40229# a_36579_40183# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X23476 VSS a_23993_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23477 a_30415_50871# a_30573_52271# a_30561_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23478 a_41370_69222# a_12901_66959# a_41862_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23479 a_27406_15516# a_16746_15514# a_27314_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2348 a_7183_42845# a_6559_42479# a_7075_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X23480 vcm_commonmode a_16362_63198# a_36442_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23481 VSS a_4343_60405# a_4274_60431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23482 a_9983_18870# a_5671_21495# a_9911_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23483 VSS a_1923_73087# a_10097_69501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23484 a_13984_43781# a_13015_43493# a_13888_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23485 a_6713_37903# a_6683_37815# a_6641_37903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23486 a_19282_64202# a_11067_13095# a_19774_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23487 a_26706_57174# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23488 a_23790_62516# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23489 a_38101_38565# a_38315_39141# a_39188_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2349 a_32795_44031# a_31004_44869# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X23490 a_47790_71230# a_12947_71576# a_47394_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23491 VSS VSS a_30722_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23492 a_2847_51157# a_2672_51183# a_3026_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23493 a_42466_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23494 vcm_commonmode a_16362_11500# a_28410_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23495 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23496 a_11179_9981# a_1586_18695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23497 VDD a_2235_30503# a_25450_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23498 a_11978_29967# a_12120_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23499 a_27806_19500# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X235 a_28410_62194# a_16746_62196# a_28318_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2350 a_29718_70226# a_12901_66665# a_29322_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23500 VDD a_13576_37149# a_12677_36893# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X23501 a_12369_40517# a_12677_40157# a_12249_43457# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X23502 a_15959_36415# a_13097_35279# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23503 VSS a_4187_60673# a_4148_60547# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23504 a_11035_47893# a_10860_47919# a_11214_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23505 a_3229_16617# a_3023_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23506 a_3487_73865# a_3137_73493# a_3392_73853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23507 a_45782_23914# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23508 a_4404_45743# a_4259_45199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23509 a_2518_22895# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2351 vcm_commonmode a_16362_18528# a_17366_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23510 a_46482_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23511 VDD a_3063_9295# a_3247_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23512 a_27183_34789# a_23567_35507# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23513 a_31004_40743# a_30035_40767# a_30908_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23514 a_5418_65327# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23515 a_12579_44310# a_12549_44212# a_12507_44310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23516 a_22294_58178# a_16362_58178# a_22386_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23517 a_35742_15882# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23518 VSS a_12895_13967# a_38754_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23519 a_42770_16886# a_12727_13353# a_42374_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2352 VDD a_11619_56615# a_12754_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X23520 VSS a_18844_43439# a_18950_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23521 a_17366_64202# a_16746_64204# a_17274_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23522 a_22294_17890# a_12899_10927# a_22786_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23523 VSS a_12947_23413# a_22690_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23524 a_19374_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23525 a_4255_59049# a_3141_59887# a_4037_58773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23526 a_7567_66781# a_7387_66781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23527 VSS a_30007_38695# a_13669_39605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X23528 a_34434_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23529 a_43870_59504# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2353 a_17569_29423# a_14926_31849# a_17497_29423# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23530 a_11667_63303# a_11145_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23531 a_39758_14878# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23532 a_76365_40202# a_76461_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23533 vcm_commonmode a_16362_70226# a_22386_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23534 VSS a_1643_64213# a_1591_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23535 a_28714_17890# a_12899_11471# a_28318_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23536 VDD a_12985_25615# a_16961_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23537 VSS a_10899_28879# a_13047_29575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23538 VDD a_6607_13879# a_6327_14343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23539 a_41766_63198# a_15439_49525# a_41370_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2354 a_9529_71677# a_9150_71311# a_9457_71677# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X23540 a_26310_55166# VSS a_26802_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23541 a_32334_9858# a_16362_9492# a_32426_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23542 VSS a_4842_45467# a_5173_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23543 VDD a_12727_58255# a_20286_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23544 a_9983_18543# a_9729_18870# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23545 vcm_commonmode a_16362_61190# a_25398_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23546 a_35838_24520# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23547 a_33049_28585# a_30788_28487# a_32772_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23548 VSS a_7050_53333# a_6996_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23549 VSS a_12727_15529# a_29718_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2355 a_21382_16520# a_16746_16518# a_21290_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23550 a_26706_10862# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23551 a_7637_69679# a_2686_70223# a_7553_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23552 a_9654_65577# a_9624_65301# a_9280_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23553 a_32730_65206# a_10975_66407# a_32334_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23554 a_11141_65327# a_10975_65327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23555 VSS a_3759_39991# a_3705_40079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23556 a_45782_64202# a_12355_65103# a_45386_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23557 vcm_commonmode a_16362_60186# a_29414_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23558 vcm_commonmode a_16362_19532# a_29414_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23559 a_36350_20902# a_12985_7663# a_36842_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2356 VSS a_6791_70455# a_6598_69653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X23560 a_39854_23516# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23561 a_39454_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23562 a_36350_16886# a_16362_16520# a_36442_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23563 vcm_commonmode a_16362_14512# a_30418_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23564 VDD a_12985_7663# a_43378_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23565 a_40458_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23566 VSS a_7624_68021# a_7571_68047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X23567 a_46482_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23568 a_43378_62194# a_16362_62194# a_43470_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23569 VDD a_2847_9813# a_2834_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2357 a_30818_18496# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23570 a_35742_56170# a_12257_56623# a_35346_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23571 a_26310_72234# VSS a_26402_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23572 a_37750_7850# VDD a_37354_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23573 VDD a_12877_16911# a_33338_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23574 a_18579_27399# a_7571_29199# a_18753_27275# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23575 VDD a_30091_35253# a_29177_34753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23576 a_30418_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23577 vcm_commonmode a_16362_67214# a_42466_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23578 VSS a_2847_45503# a_2781_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X23579 a_18674_66210# a_12983_63151# a_18278_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2358 a_36579_35831# a_12621_36091# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X23580 a_25145_30083# a_25263_29981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23581 VSS a_8569_25071# a_9043_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23582 a_28430_32143# a_14646_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23583 VSS a_12546_22351# a_42770_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23584 VDD a_10055_58791# a_46390_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23585 a_44474_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23586 VDD a_11067_21583# a_29322_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23587 a_20378_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23588 VSS a_12546_22351# a_18674_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23589 a_2107_23817# a_1591_23445# a_2012_23805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2359 VSS a_11803_55311# a_16746_69224# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X23590 VSS a_7637_53877# a_3228_54171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X23591 VSS VDD a_23694_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23592 a_9740_62973# a_7676_61493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X23593 VSS a_3016_60949# a_5443_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23594 a_28714_9858# a_12985_19087# a_28318_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23595 VDD a_12727_15529# a_19282_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23596 a_28618_32143# a_14646_29423# a_27417_32509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23597 a_27251_30083# a_14926_31849# a_27169_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23598 VDD a_13445_50639# a_12683_51329# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23599 a_17366_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X236 a_6649_25615# a_4571_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=0p ps=0u w=650000u l=150000u M=4
X2360 a_9931_62985# a_9485_62613# a_9835_62985# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X23600 a_32426_66210# a_16746_66212# a_32334_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23601 a_11304_18543# a_10961_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23602 a_31330_21906# a_16362_21540# a_31422_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23603 VSS a_4889_55535# a_5258_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23604 VDD a_15439_49525# a_41370_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23605 VSS a_35217_44509# a_34909_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23606 a_9544_61635# a_9526_61751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23607 a_39454_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23608 a_4174_53181# a_3668_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23609 vcm_commonmode a_16362_68218# a_19374_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2361 VSS a_32649_28853# a_31768_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23610 a_7505_65327# a_7126_65693# a_7433_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23611 VDD a_12663_40871# a_14081_42134# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23612 vcm_commonmode a_16362_57174# a_49494_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23613 a_30722_61190# a_12355_15055# a_30326_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23614 VSS a_29927_29199# a_33689_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23615 a_27425_47375# a_4891_47388# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23616 VSS a_10515_22671# a_35742_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23617 a_42374_71230# a_12901_66665# a_42866_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23618 a_8638_65103# a_8782_65015# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23619 a_38358_61190# a_12981_59343# a_38850_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2362 a_14079_36694# a_13349_37973# a_13620_36519# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X23620 a_46390_69222# a_16362_69222# a_46482_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23621 a_32509_47919# a_27869_50095# a_32406_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23622 VDD a_12981_62313# a_45386_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23623 a_10863_16733# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23624 a_14109_31055# a_9765_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23625 VSS a_4811_34855# a_32319_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X23626 VDD a_26514_47375# a_30079_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23627 a_32611_39141# a_30912_39429# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23628 VDD a_2847_44629# a_2834_45021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23629 a_36097_51727# a_29361_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2363 VSS a_16928_36391# a_16891_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X23630 VDD a_7841_22895# a_11771_23671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23631 VDD a_2713_35925# a_2743_36278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23632 a_35463_42943# a_33856_42693# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23633 vcm_commonmode a_16362_9492# a_34434_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23634 a_29915_29423# a_28841_29575# a_28963_28853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23635 a_26402_57174# a_16746_57176# a_26310_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23636 a_27710_18894# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23637 a_4333_22895# a_3985_22901# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X23638 a_25798_8456# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23639 VSS a_12899_11471# a_31726_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2364 VSS a_6792_43719# a_5715_44343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23640 a_21686_8854# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23641 a_30875_34743# a_29943_34789# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23642 a_15211_50959# a_14985_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23643 a_40458_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23644 a_44474_9492# a_16746_9490# a_44382_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23645 VDD a_12895_13967# a_49402_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23646 a_38524_28585# a_36904_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23647 VDD a_12355_65103# a_18278_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23648 VSS a_3339_43023# a_12227_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23649 a_2865_58799# a_2695_58799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2365 a_34434_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23650 VSS a_12901_66959# a_43774_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23651 a_40762_66210# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23652 a_4974_56875# a_5252_56891# a_5208_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23653 VDD a_10791_15529# a_11714_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23654 a_32334_59182# a_12901_58799# a_32826_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23655 a_6829_15055# a_5755_14709# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23656 a_22352_40517# a_21479_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23657 a_20853_47375# a_20575_47713# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X23658 VSS a_23784_42583# a_23597_42325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23659 a_19282_72234# VDD a_19774_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2366 VDD a_9187_10901# a_8556_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X23660 vcm_commonmode a_16362_20536# a_42466_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23661 a_17211_49373# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23662 VSS a_5239_65301# a_5173_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23663 VDD a_3449_54201# a_3479_53942# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23664 a_23790_70548# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23665 a_44474_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23666 a_41370_55166# VSS a_41462_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23667 VSS a_12981_62313# a_30722_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23668 VSS a_1929_12131# a_8815_13879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23669 a_3254_9334# a_1689_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2367 vcm_commonmode a_16362_12504# a_31422_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23670 a_5957_74031# a_5913_74273# a_5791_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X23671 a_19774_60508# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23672 a_40458_71230# a_16746_71232# a_40366_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23673 a_7938_11587# a_1929_10651# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23674 a_27406_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23675 a_7445_63695# a_6913_64239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23676 a_20682_69222# a_12516_7093# a_20286_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23677 a_44778_65206# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23678 a_44874_17492# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23679 a_44778_23914# a_10515_23975# a_44382_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2368 vcm_commonmode a_16362_63198# a_43470_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23680 a_7267_62063# a_7213_62215# a_7077_62313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23681 a_41370_14878# a_12877_14441# a_41862_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23682 a_77568_40202# a_77664_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23683 a_42374_18894# a_16362_18528# a_42466_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23684 a_8011_48463# a_7387_48469# a_7903_48841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23685 VSS a_1923_59583# a_4761_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23686 a_34738_57174# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23687 a_11990_21583# a_9955_21807# a_11763_21237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9825e+11p ps=1.91e+06u w=650000u l=150000u
X23688 VSS a_4339_64521# a_9177_60214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23689 a_34738_15882# a_12877_14441# a_34342_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2369 a_19678_62194# a_12981_62313# a_19282_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23690 a_17670_67214# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23691 a_44474_70226# a_16746_70228# a_44382_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23692 a_12786_30761# a_12161_31849# a_12714_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23693 a_8177_37013# a_6372_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23694 VSS a_12355_65103# a_21686_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23695 a_47790_56170# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23696 VDD a_12899_11471# a_21290_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23697 a_48890_16488# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23698 a_45386_13874# a_12727_15529# a_45878_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23699 a_10521_25731# a_9751_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X237 vcm_commonmode a_16362_18528# a_25398_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2370 a_20682_58178# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23700 a_20897_42917# a_21479_42405# a_22411_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X23701 vcm_commonmode a_16362_21540# a_19374_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23702 a_28318_23914# a_12947_23413# a_28810_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23703 a_28318_19898# a_16362_19532# a_28410_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23704 a_34434_62194# a_16746_62196# a_34342_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23705 vcm_commonmode a_16362_10496# a_49494_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23706 vcm_commonmode a_16362_8488# a_23390_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23707 a_13067_38517# a_27219_44011# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X23708 a_35838_58500# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23709 VSS a_11763_20407# a_10275_21495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2371 a_10901_54201# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23710 a_32826_21508# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23711 a_32426_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23712 a_12921_40719# a_12651_41085# a_12831_41085# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23713 a_17366_72234# VDD a_17274_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23714 a_38754_14878# a_12727_15529# a_38358_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23715 VSS a_10055_58791# a_35742_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23716 a_47486_61190# a_16746_61192# a_47394_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23717 VDD a_10409_18543# a_10791_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23718 a_27710_59182# a_12727_58255# a_27314_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23719 VSS a_12947_56817# a_24698_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2372 a_34738_71230# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23720 a_18278_15882# a_12727_13353# a_18770_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23721 a_5333_59343# a_1952_60431# a_5261_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23722 VSS a_19492_52245# a_12659_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X23723 VDD a_12727_13353# a_25306_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23724 a_22786_13476# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23725 a_24743_48437# a_25015_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23726 a_5291_56765# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X23727 a_39362_69222# a_12901_66959# a_39854_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23728 a_53218_40254# a_52778_39198# a_7841_12167# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23729 a_43870_67536# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2373 a_33430_69222# a_16746_69224# a_33338_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23730 a_10403_48285# a_9779_47919# a_10295_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23731 a_40366_64202# a_11067_13095# a_40858_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23732 a_26402_10496# a_16746_10494# a_26310_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23733 a_7381_35727# a_5963_36585# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23734 a_33338_13874# a_16362_13508# a_33430_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23735 a_11415_58077# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23736 a_9835_62985# a_9485_62613# a_9740_62973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23737 vcm_commonmode a_16362_16520# a_48490_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23738 VSS VSS a_28714_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23739 a_32765_31287# a_4811_34855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2374 a_46882_7452# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23740 a_1823_53885# a_2939_52245# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23741 a_8268_35381# a_6372_38279# a_8491_35727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23742 a_28638_30083# a_20267_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23743 VSS a_1586_40455# a_4535_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23744 VSS a_10515_23975# a_43774_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23745 VDD a_12727_67753# a_20286_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23746 a_10969_59663# a_11115_59317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23747 VDD a_4095_29423# a_4497_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23748 VDD a_19576_51701# a_21095_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23749 VSS a_6786_37557# a_6713_37903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2375 a_42770_7850# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X23750 a_29814_68540# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23751 a_2872_59893# a_2685_59933# a_2785_60151# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X23752 VSS a_2216_42997# a_2150_43401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23753 a_8500_58799# a_7871_59049# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X23754 a_30818_63520# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23755 a_25398_16520# a_16746_16518# a_25306_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23756 VSS a_76648_39738# a_76461_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23757 a_37888_34191# a_37711_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23758 a_1846_73195# a_2163_73085# a_2121_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23759 a_34342_55166# a_8295_47388# a_34834_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2376 VDD a_17843_48981# a_17830_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X23760 a_20682_22910# a_11067_21583# a_20286_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23761 VDD a_24844_47753# a_25019_47679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23762 a_27105_48169# a_26465_48463# a_26917_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23763 a_27245_41829# a_26815_42405# a_27688_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23764 a_17274_65206# a_12355_65103# a_17766_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23765 a_10253_23759# a_7841_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23766 a_38754_71230# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23767 a_37446_69222# a_16746_69224# a_37354_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23768 a_45782_72234# VDD a_45386_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23769 a_38115_52263# a_38524_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2377 VDD a_12381_43957# a_12793_44310# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23770 a_36350_24918# VSS a_36442_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23771 a_2244_18231# config_1_in[10] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23772 a_34738_10862# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23773 a_40458_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23774 a_10973_16609# a_10755_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23775 VDD a_12801_38517# a_24382_41629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23776 a_10053_62581# a_9835_62985# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23777 a_1761_47919# a_1591_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X23778 a_17670_20902# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23779 VDD a_11067_63143# a_12541_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2378 VSS a_2292_43291# a_7125_46653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X23780 a_35581_31849# a_11067_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23781 VDD a_10515_22671# a_27314_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23782 a_36465_49551# a_36551_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23783 vcm_commonmode a_16362_65206# a_38450_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23784 VSS a_8453_51727# a_9278_55311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23785 a_43774_24918# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23786 a_2744_66103# a_2952_66139# a_2886_66237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23787 a_32730_69222# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23788 a_11801_68047# a_11947_68279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23789 a_14039_34743# a_13107_34789# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2379 a_33734_57174# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23790 a_27710_12870# a_10055_58791# a_27314_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23791 a_5791_74031# a_5345_74031# a_5695_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23792 a_34342_72234# VSS a_34434_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23793 VSS a_12727_58255# a_36746_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23794 VDD a_3911_16065# a_3872_15939# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23795 VSS a_11067_67279# a_36746_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23796 a_12263_20969# a_12323_20904# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23797 VSS a_12516_7093# a_19678_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23798 a_33338_58178# a_16362_58178# a_33430_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23799 a_47394_71230# a_16362_71230# a_47486_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X238 a_35838_22512# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2380 a_35099_43447# a_35493_43421# a_30412_42589# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X23800 a_46786_15882# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23801 VSS a_12895_13967# a_49798_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23802 a_20286_18894# a_12895_13967# a_20778_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23803 VSS VSS a_20682_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23804 a_17366_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23805 a_10543_16580# a_10423_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23806 VDD a_10103_48682# a_9392_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23807 VDD a_11067_21583# a_37354_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23808 vcm_commonmode a_16362_15516# a_24394_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23809 VDD a_12947_71576# a_41370_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2381 a_35838_70548# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23810 a_33338_17890# a_12899_10927# a_33830_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23811 a_14859_38909# a_13669_38517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23812 a_37733_37477# a_38315_38053# a_39188_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X23813 a_48398_8854# a_12985_19087# a_48890_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23814 a_41462_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23815 a_10984_58487# a_11080_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23816 VDD a_7571_29199# a_18487_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23817 a_17799_38591# a_17033_38565# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X23818 a_11507_72221# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23819 a_7126_65693# a_7039_65469# a_6722_65579# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X2382 VSS a_12546_22351# a_35742_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23820 a_24394_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23821 a_11121_23957# a_7571_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23822 a_26706_18894# a_12899_10927# a_26310_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23823 vcm_commonmode a_16362_70226# a_33430_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23824 a_4351_26703# a_3301_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23825 VDD a_12901_66665# a_45386_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23826 a_4220_68021# a_3693_68047# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23827 a_38450_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23828 a_35346_11866# a_16362_11500# a_35438_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23829 a_4052_73865# a_2971_73493# a_3705_73461# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2383 a_30561_50639# a_30663_51727# a_30415_50871# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X23830 a_24302_19898# a_11067_67279# a_24794_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23831 VSS a_33155_35839# a_33101_36161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23832 vcm_commonmode a_16362_62194# a_23390_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23833 a_41334_29575# a_41232_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23834 a_18158_47158# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23835 a_28410_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23836 VDD a_12727_58255# a_31330_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23837 a_5462_18365# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23838 VSS a_12877_14441# a_27710_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23839 a_37446_22544# a_16746_22542# a_37354_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2384 a_25744_7638# a_37699_27221# a_37471_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X23840 VDD VDD a_18278_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23841 a_2215_14735# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23842 VDD a_12947_8725# a_35346_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23843 a_18370_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23844 a_8827_29967# a_6649_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23845 VSS a_12983_63151# a_39758_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23846 a_36746_64202# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23847 VDD a_2560_45895# a_2007_45717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23848 a_32334_67214# a_12983_63151# a_32826_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23849 a_43774_65206# a_10975_66407# a_43378_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2385 VDD a_7159_50260# a_6863_49722# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X23850 a_5531_53903# a_5258_54223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23851 a_41766_8854# a_12947_8725# a_41370_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23852 VSS a_2244_18231# a_2021_17973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23853 a_2291_47753# a_1941_47381# a_2196_47741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23854 a_41370_63198# a_16362_63198# a_41462_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23855 a_7183_45199# a_6559_45205# a_7075_45577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23856 a_11491_55535# a_11141_55535# a_11396_55535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23857 a_24067_42583# a_14258_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23858 a_33734_57174# a_10515_22671# a_33338_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23859 a_17670_8854# a_12947_8725# a_17274_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2386 a_24746_31849# a_23119_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23860 a_32730_22910# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23861 VSS a_38454_43983# a_38999_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23862 a_29322_21906# a_16362_21540# a_29414_21540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23863 vcm_commonmode a_16362_68218# a_40458_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23864 VSS a_1643_63125# a_1591_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23865 a_19500_44869# a_18627_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23866 VDD a_2672_18543# a_2847_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23867 a_46786_56170# a_12257_56623# a_46390_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23868 VDD a_12877_16911# a_44382_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23869 a_29718_66210# a_12983_63151# a_29322_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2387 a_38450_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23870 a_36600_49159# a_4351_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23871 VSS a_10299_47607# a_10195_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X23872 a_3410_70589# a_3372_70197# a_2824_70197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23873 a_2250_56989# a_2124_56891# a_1846_56875# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X23874 a_20747_27765# a_10873_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23875 a_15941_31055# a_14097_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23876 a_33264_37601# a_32795_38053# a_33727_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X23877 VSS a_23901_44220# a_23593_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23878 vcm_commonmode a_16362_59182# a_43470_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23879 a_32785_50639# a_26397_51183# a_32370_50871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2388 a_35346_60186# a_16362_60186# a_35438_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23880 vcm_commonmode a_16362_69222# a_26402_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23881 a_48490_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23882 a_7273_56623# a_6835_46823# a_6927_56873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23883 a_30418_67214# a_16746_67216# a_30326_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23884 a_24755_42325# a_12641_43124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23885 VDD a_12516_7093# a_38358_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23886 a_35838_66532# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23887 a_10317_55223# a_7155_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23888 a_43539_29967# a_20267_30503# a_43321_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23889 a_9963_13760# a_9083_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2389 a_6567_25615# a_5211_24759# a_6985_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X23890 a_19374_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23891 a_8957_65103# a_8896_65015# a_8638_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23892 a_38450_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23893 a_35346_56170# a_16362_56170# a_35438_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23894 a_2215_49551# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23895 a_21686_61190# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23896 VDD a_8753_66103# a_7987_64213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X23897 a_20378_59182# a_16746_59184# a_20286_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23898 vcm_commonmode a_16362_58178# a_47486_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23899 a_18278_66210# a_16362_66210# a_18370_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X239 a_38454_43983# a_38277_43983# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2390 a_20378_63198# a_16746_63200# a_20286_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X23900 a_33430_8488# a_16746_8486# a_33338_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23901 VDD VDD a_24302_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23902 VSS VDD a_20682_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23903 a_40366_72234# VDD a_40858_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23904 a_39854_65528# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23905 a_36350_62194# a_12355_15055# a_36842_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23906 a_40858_60508# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23907 a_49402_22910# a_10515_23975# a_49894_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23908 VDD a_30716_51701# a_30663_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X23909 a_6375_64489# a_4119_70741# a_6457_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2391 VSS a_1761_22895# a_33155_40191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X23910 VDD a_17280_48695# a_17095_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23911 a_39362_55166# VSS a_39454_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23912 VSS a_12981_62313# a_28714_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23913 a_25702_60186# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23914 VDD a_3509_58487# a_2695_58951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X23915 a_24394_58178# a_16746_58180# a_24302_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23916 vcm_commonmode VSS a_21382_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23917 a_25702_19898# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23918 a_38450_71230# a_16746_71232# a_38358_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23919 VDD a_11067_63143# a_12723_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2392 a_45478_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23920 VSS a_12381_35836# a_12325_35862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X23921 VSS a_12677_36893# a_12369_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23922 VDD a_12869_2741# a_33338_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23923 a_39362_14878# a_12877_14441# a_39854_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23924 a_1915_11092# a_2007_10901# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23925 VSS a_12985_7663# a_39758_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23926 VSS a_20747_27765# a_20514_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23927 a_9370_58575# a_7210_55081# a_9560_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23928 a_43870_12472# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23929 a_26802_22512# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2393 a_18278_70226# a_16362_70226# a_18370_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X23930 a_31440_32259# a_27535_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23931 a_8143_47919# a_7889_48246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23932 a_2764_33609# a_1849_33237# a_2417_33205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23933 a_30818_71552# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23934 a_16362_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23935 VDD a_11067_67279# a_30326_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23936 VDD a_12355_65103# a_29322_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23937 VDD a_23789_39100# a_23733_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X23938 a_30326_61190# a_16362_61190# a_30418_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23939 a_33734_10862# a_12546_22351# a_33338_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2394 VSS a_2926_15253# a_2867_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X23940 a_17867_32117# a_17672_32259# a_18177_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23941 VDD a_15607_46805# a_40691_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X23942 VSS a_16863_29415# a_39299_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23943 a_77002_39738# a_77098_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X23944 VSS a_2292_43291# a_7337_45565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23945 a_4987_52508# a_4831_52413# a_5132_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23946 vcm_commonmode a_16362_21540# a_40458_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23947 a_43470_24552# VDD a_43378_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23948 a_2781_45577# a_1591_45205# a_2672_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23949 VDD a_10055_58791# a_20286_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2395 vcm_commonmode a_16362_65206# a_34434_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23950 VDD a_12257_56623# a_19282_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23951 a_6453_71855# a_5975_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23952 a_12671_43222# a_12641_43124# a_12599_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23953 a_27314_14878# a_16362_14512# a_27406_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23954 a_33430_16520# a_16746_16518# a_33338_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X23955 VSS a_20351_49525# a_20282_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23956 a_42866_18496# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23957 VSS a_29943_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X23958 a_31422_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23959 a_31726_69222# a_12516_7093# a_31330_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2396 VSS VDD a_28714_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23960 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X23961 a_46482_15516# a_16746_15514# a_46390_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23962 vcm_commonmode a_16362_12504# a_43470_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23963 a_7467_57863# a_6559_59663# a_7634_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23964 a_17274_10862# a_12985_16367# a_17766_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23965 vcm_commonmode a_16362_22544# a_26402_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23966 a_22386_7484# VDD a_22294_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23967 VSS a_76648_40202# a_76461_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23968 VSS a_17682_50095# a_29915_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23969 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2397 a_26020_30199# a_14926_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X23970 a_30418_20536# a_16746_20534# a_30326_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23971 a_45782_57174# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23972 a_5023_13255# a_3983_12879# a_5169_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23973 VSS a_13669_35253# a_14088_35279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23974 a_28714_67214# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23975 a_19374_17524# a_16746_17522# a_19282_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23976 VDD a_9275_15253# a_9963_13760# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23977 VDD a_7195_65564# a_7126_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23978 VSS a_5190_59575# a_11801_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23979 VSS a_12355_65103# a_32730_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2398 a_10526_22057# a_6559_22671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X23980 a_20378_12504# a_16746_12502# a_20286_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23981 a_28157_40747# a_22671_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23982 vcm_commonmode a_16362_11500# a_47486_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23983 a_5825_20175# a_3987_19623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23984 a_30418_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23985 a_42866_9460# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23986 a_1915_45908# a_2007_45717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X23987 a_24279_47753# a_23763_47381# a_24184_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23988 a_2196_47741# a_2079_47546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23989 a_46882_19500# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2399 VDD a_12546_22351# a_38358_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X23990 a_11697_62063# a_11145_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23991 a_45478_62194# a_16746_62196# a_45386_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23992 a_18674_59182# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23993 a_20286_69222# a_16362_69222# a_20378_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23994 VSS a_12257_56623# a_22690_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23995 a_21615_49007# a_21169_49007# a_21519_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23996 VDD a_4119_70741# a_3983_70767# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23997 a_18770_9460# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X23998 a_49798_14878# a_12727_15529# a_49402_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23999 a_28810_63520# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24 a_1923_59583# a_2511_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X240 a_29814_58500# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2400 a_33734_9858# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24000 a_11587_60975# a_11141_60975# a_11491_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24001 a_17867_32117# a_17711_32385# a_18012_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24002 a_34639_37737# a_35033_37692# a_34699_37683# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X24003 a_24394_11500# a_16746_11498# a_24302_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24004 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24005 VDD a_12985_19087# a_28318_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24006 a_35165_52093# a_34895_51727# a_35061_51727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24007 VDD a_10379_66389# a_9914_68279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24008 VDD a_12895_13967# a_23298_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24009 VDD a_4495_35925# a_4985_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2401 vcm_commonmode a_16362_64202# a_47486_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24010 a_36720_49551# a_30928_49007# a_36465_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24011 a_24302_68218# a_16362_68218# a_24394_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24012 a_36442_64202# a_16746_64204# a_36350_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24013 VSS a_2411_26133# a_5037_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24014 VSS a_40737_37692# a_40429_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24015 VSS a_12947_23413# a_41766_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24016 a_38450_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24017 a_5805_74575# a_5599_74549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24018 a_41370_56170# a_12947_56817# a_41862_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24019 a_2319_54684# a_2124_54715# a_2629_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2402 VDD a_4351_26703# a_8215_25071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X24020 a_5309_25853# a_5087_24643# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X24021 a_27806_69544# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24022 VDD a_12727_67753# a_31330_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24023 a_9280_65327# a_2840_66103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24024 a_27314_59182# a_16362_59182# a_27406_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24025 VSS a_5877_54421# a_5336_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24026 a_31422_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24027 VSS a_20505_29967# a_22727_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24028 a_47790_17890# a_12899_11471# a_47394_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24029 a_14293_37455# a_13867_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2403 a_49402_22910# a_16362_22544# a_49494_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24030 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24031 a_32029_38565# a_32611_39141# a_33543_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24032 a_23392_31599# a_5915_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24033 a_26310_9858# a_16362_9492# a_26402_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24034 a_36746_72234# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24035 a_45386_55166# VSS a_45878_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24036 a_31726_22910# a_11067_21583# a_31330_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24037 VSS a_12516_7093# a_40762_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24038 a_1644_62037# a_1591_59343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24039 VSS a_32795_29967# a_33515_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X2404 a_36746_68218# a_12901_66959# a_36350_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24040 VDD a_4758_45369# a_5357_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24041 a_28318_65206# a_12355_65103# a_28810_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24042 a_4642_54991# a_4516_55107# a_4238_55123# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24043 a_28244_31415# a_25313_31599# a_28172_31415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24044 a_8671_22351# a_5531_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24045 vcm_commonmode a_16362_61190# a_44474_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24046 vcm_commonmode a_16362_71230# a_27406_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24047 VSS a_12727_15529# a_48794_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24048 a_45782_10862# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24049 VSS a_15253_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X2405 VSS a_1586_9991# a_5639_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24050 a_18278_57174# a_12257_56623# a_18770_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24051 a_22786_55488# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24052 a_2012_12925# a_1895_12730# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24053 a_28714_20902# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24054 a_32887_44581# a_32121_44545# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X24055 a_32334_12870# a_12877_16911# a_32826_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24056 VDD a_23271_50943# a_23258_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24057 a_21382_61190# a_16746_61192# a_21290_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24058 VSS a_3949_41935# a_5731_40079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24059 a_37354_7850# VDD a_37846_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2406 VSS a_2411_26133# a_3749_37949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X24060 a_18674_12870# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24061 a_17008_49007# a_16891_49220# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24062 a_25702_13874# a_12877_16911# a_25306_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24063 VSS a_12985_16367# a_22690_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24064 a_5381_68345# a_2843_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24065 a_7969_58799# a_7107_58487# a_8060_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24066 vcm_commonmode VSS a_32426_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24067 VSS a_17039_51157# a_21873_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24068 a_47886_7452# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24069 a_43774_7850# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2407 a_31243_35831# a_30311_35877# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X24070 a_45386_72234# VSS a_45478_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24071 VSS a_12727_58255# a_47790_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24072 a_15788_28335# a_13390_29575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24073 VSS a_11067_67279# a_47790_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24074 a_37750_66210# a_12983_63151# a_37354_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24075 VSS a_7464_39215# a_7847_40847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24076 a_19678_7850# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24077 VDD a_10515_23975# a_35346_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24078 vcm_commonmode a_16362_16520# a_22386_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24079 a_31330_18894# a_12895_13967# a_31822_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2408 VSS a_18579_27399# a_17278_28309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24080 a_5913_11169# a_5695_10927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24081 VSS a_34482_29941# a_37553_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24082 a_35346_64202# a_16362_64202# a_35438_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24083 a_28056_44869# a_27183_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24084 VDD a_11067_21583# a_48398_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24085 VSS VDD a_29718_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24086 VDD a_26433_39631# a_29915_41959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24087 a_8071_48246# a_7889_48246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24088 a_22386_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24089 vcm_commonmode a_16362_69222# a_34434_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2409 VSS a_15011_34717# a_14951_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X24090 a_24698_60186# a_12981_59343# a_24302_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24091 a_24698_19898# a_12895_13967# a_24302_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24092 VDD a_27869_50095# a_29715_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24093 VSS a_2345_33749# a_2279_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24094 a_16615_39095# a_16043_38825# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X24095 a_36350_70226# a_12516_7093# a_36842_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24096 VDD a_12727_15529# a_38358_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24097 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24098 a_41636_37601# a_41351_38053# a_42283_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24099 VDD a_1586_18695# a_7571_16917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X241 a_20778_8456# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2410 VSS a_13909_41923# a_40527_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X24100 a_36442_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24101 VDD a_8423_39367# a_8377_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24102 VDD a_3019_13621# a_4075_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24103 a_4627_23439# a_3983_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24104 a_35412_51433# a_35382_51157# a_35069_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24105 a_39362_63198# a_16362_63198# a_39454_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24106 vcm_commonmode a_16362_63198# a_21382_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24107 a_49494_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24108 a_46390_11866# a_16362_11500# a_46482_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24109 a_8162_53609# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2411 vcm_commonmode a_16362_56170# a_37446_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24110 a_9945_73807# a_9353_72399# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24111 a_35438_23548# a_16746_23546# a_35346_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24112 a_1941_47381# a_1775_47381# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24113 a_39854_10464# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24114 a_2125_34863# a_1915_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24115 VDD a_8556_10357# a_8494_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24116 a_4717_45985# a_4499_45743# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24117 VSS a_2283_15797# a_4229_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24118 a_10851_16367# a_10405_16367# a_10755_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24119 a_11372_12381# a_10935_11989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2412 a_49798_67214# a_12727_67753# a_49402_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24120 a_2781_21807# a_1591_21807# a_2672_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24121 a_13891_36189# a_13743_35836# a_13528_36055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24122 a_4798_23759# a_3983_24233# a_4712_23759# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X24123 a_31350_47919# a_26397_51183# a_31031_47919# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u w=650000u l=150000u
X24124 VDD VDD a_29322_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24125 VSS a_12727_67753# a_37750_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24126 a_15315_27791# a_15064_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24127 VDD a_10506_29967# a_14167_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24128 a_26251_30083# a_25263_29981# a_26155_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24129 a_29414_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2413 a_42770_15882# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24130 a_21686_9858# a_12985_19087# a_21290_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24131 vcm_commonmode VSS a_45478_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24132 a_2834_51549# a_1757_51183# a_2672_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24133 a_4345_69679# a_2686_70223# a_4357_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24134 a_28410_67214# a_16746_67216# a_28318_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24135 vcm_commonmode a_16362_64202# a_25398_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24136 a_8205_26159# a_3607_34639# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24137 a_30722_23914# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24138 VSS a_13643_28327# a_39391_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24139 a_27314_22910# a_16362_22544# a_27406_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2414 VSS a_34145_49007# a_36821_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X24140 a_8209_39465# a_8021_39221# a_8127_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24141 VDD a_12355_65103# a_37354_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24142 a_34834_61512# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24143 VSS a_10299_11703# a_9642_10357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24144 a_30125_47919# a_26397_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24145 a_5064_48841# a_4149_48469# a_4717_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24146 a_31422_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24147 a_6619_47607# a_6727_47607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24148 a_42466_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24149 a_44778_57174# a_10515_22671# a_44382_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2415 a_7862_10383# a_7736_10499# a_7458_10515# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X24150 VSS a_10288_17143# a_10239_16911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24151 VSS a_1923_59583# a_1881_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24152 a_4726_20214# a_3247_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X24153 VDD a_2011_34837# a_1887_34863# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24154 a_19678_61190# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24155 a_18370_59182# a_16746_59184# a_18278_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24156 VDD a_1586_40455# a_1591_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24157 a_20682_15882# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24158 VSS a_12895_13967# a_23694_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24159 a_3680_57527# a_1591_57711# a_3608_57527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2416 VSS a_13357_32143# a_25605_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24160 VSS a_4215_51157# a_18335_50645# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24161 a_10747_52854# a_6559_59663# a_10288_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24162 a_6625_29941# a_5993_32687# a_6878_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24163 a_30326_7850# VSS a_30418_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24164 a_38850_60508# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24165 a_11602_25071# a_11163_25321# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X24166 a_46482_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24167 VSS a_3063_9295# a_3247_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X24168 a_30530_51183# a_28881_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24169 a_13123_38231# a_32831_35307# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X2417 a_24394_64202# a_16746_64204# a_24302_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24170 vcm_commonmode VSS a_19374_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24171 VDD a_8540_42167# a_8383_43255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24172 a_2939_31573# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24173 a_24698_14878# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24174 a_22649_27791# a_22562_28023# a_22567_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24175 vcm_commonmode a_16362_22544# a_34434_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24176 a_43378_24918# VSS a_43870_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24177 VSS a_5839_22351# a_6743_23555# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24178 VDD a_16228_28335# a_17415_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24179 VDD a_12516_7093# a_49402_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2418 a_3955_24643# a_2315_24540# a_3883_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24180 a_27797_29423# a_27422_29789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24181 VSS a_9031_54135# a_6236_54421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24182 a_28810_71552# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24183 a_49494_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24184 a_46390_56170# a_16362_56170# a_46482_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24185 VDD a_11455_12157# a_11416_12283# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24186 VDD a_3143_22364# a_3779_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24187 VSS a_38499_37503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24188 a_10480_55107# a_7155_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24189 a_2847_18517# a_2672_18543# a_3026_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2419 a_32612_51727# a_2775_46025# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X24190 VDD a_12899_11471# a_40366_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24191 a_28027_29217# a_25269_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24192 a_49798_66210# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24193 a_17803_44265# a_18197_44220# a_17863_44211# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X24194 a_20778_24520# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24195 a_47394_23914# a_12947_23413# a_47886_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24196 a_40527_41271# a_40921_41245# a_13909_41923# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X24197 a_47394_19898# a_16362_19532# a_47486_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24198 VSS a_26447_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24199 a_1824_61127# a_1768_13103# a_2055_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X242 a_13005_35823# a_12579_35862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2420 VSS a_30127_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24200 a_19743_42359# a_18811_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24201 a_36442_72234# VDD a_36350_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24202 a_7911_21379# a_2339_38129# a_7839_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24203 VSS a_9529_28335# a_15064_27907# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24204 VSS a_12947_56817# a_43774_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24205 a_37354_15882# a_12727_13353# a_37846_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24206 VSS a_11067_21583# a_37750_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24207 a_13097_37455# a_12671_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24208 a_49494_71230# a_16746_71232# a_49402_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24209 VSS a_28680_30057# a_28426_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2421 a_3325_69135# a_2847_69439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24210 a_41862_13476# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24211 VSS a_10975_66407# a_26706_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24212 VSS a_23501_42583# a_18662_43671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24213 a_27379_39095# a_26447_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24214 a_30722_64202# a_12355_65103# a_30326_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24215 VDD VSS a_44382_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24216 a_21290_20902# a_12985_7663# a_21782_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24217 a_24794_23516# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24218 VDD a_6646_50639# a_14291_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24219 a_24394_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2422 a_26402_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24220 a_1761_22895# a_1591_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24221 a_21290_16886# a_16362_16520# a_21382_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24222 a_9289_26703# a_6773_27805# a_9135_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24223 a_3026_44655# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24224 a_12055_62973# a_11053_62607# a_11959_62973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24225 a_28410_20536# a_16746_20534# a_28318_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24226 a_31422_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24227 a_27406_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24228 a_40458_17524# a_16746_17522# a_40366_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24229 a_20682_56170# a_12257_56623# a_20286_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2423 a_10053_69109# a_9835_69513# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X24230 VDD a_12899_10927# a_17274_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24231 a_28670_30663# a_28513_29673# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X24232 a_10191_56445# a_7479_54439# a_9828_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24233 a_2561_28918# a_2011_34837# a_2347_28918# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X24234 a_5241_72765# a_3751_72373# a_5169_72765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24235 a_44778_10862# a_12546_22351# a_44382_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24236 a_10575_62911# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24237 a_7493_12015# a_3327_9308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24238 a_12671_36694# a_12641_36596# a_12599_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24239 VSS a_42188_37149# a_41289_36893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X2424 a_39758_59182# a_12727_58255# a_39362_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24240 a_18370_12504# a_16746_12502# a_18278_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24241 a_27806_14480# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24242 VDD config_1_in[4] a_1591_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X24243 a_28410_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24244 a_25306_15882# a_16362_15516# a_25398_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24245 VDD a_10055_58791# a_31330_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24246 VSS a_30125_47919# a_30633_48829# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24247 a_48890_68540# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24248 a_36442_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24249 a_6817_42255# a_6607_42167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2425 a_6980_42479# a_6863_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X24250 a_12985_19087# a_12815_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24251 a_13107_41317# a_12341_41281# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X24252 a_44474_16520# a_16746_16518# a_44382_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24253 a_2080_59343# a_1643_59317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24254 vcm_commonmode a_16362_13508# a_41462_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24255 a_25295_51183# a_24849_51183# a_25199_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24256 VSS a_26112_30663# a_26063_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X24257 a_28318_10862# a_12985_16367# a_28810_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24258 a_43774_58178# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24259 a_2847_36799# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2426 VDD a_12355_15055# a_33338_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24260 VDD a_12901_66959# a_25306_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24261 a_26706_68218# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24262 a_34337_29967# a_34482_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24263 a_49402_64202# a_11067_13095# a_49894_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24264 VDD a_2606_41079# a_7889_48246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X24265 a_9376_54223# a_9507_53877# a_9186_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24266 a_17366_18528# a_16746_18526# a_17274_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24267 a_7948_38377# a_5631_38127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24268 a_2860_17277# a_2746_16885# a_2788_17277# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24269 a_18551_29451# a_13390_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2427 a_32319_48463# a_28108_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X24270 a_23507_42089# a_23901_42044# a_23567_42035# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X24271 a_33797_29673# a_29927_29199# a_33008_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24272 a_28994_49551# a_28959_49783# a_28691_49783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24273 VDD a_12139_71829# a_12126_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24274 a_9835_62985# a_9319_62613# a_9740_62973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24275 VDD a_1586_45431# a_1591_45205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24276 a_39362_56170# a_12947_56817# a_39854_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24277 VSS a_10515_22671# a_20682_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24278 VSS a_12901_66665# a_34738_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24279 a_26802_64524# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2428 a_7195_27497# a_3301_26703# a_7113_27253# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24280 a_23298_61190# a_12981_59343# a_23790_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24281 a_31330_69222# a_16362_69222# a_31422_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24282 vcm_commonmode a_16362_14512# a_18370_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24283 a_2589_62839# a_2794_62697# a_2752_62723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24284 VDD a_12981_62313# a_30326_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24285 a_17711_32385# a_4191_33449# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24286 a_36459_47919# a_21187_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24287 a_5345_10927# a_5179_10927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24288 a_6362_14441# a_6327_14343# a_6059_14165# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24289 a_35438_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2429 VSS a_12981_59343# a_18674_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X24290 a_10405_16367# a_10239_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24291 a_12651_35645# a_12663_35431# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24292 a_9651_49929# a_9301_49557# a_9556_49917# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24293 VDD a_2686_70223# a_4935_70561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24294 a_3869_16189# a_3391_15797# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24295 VSS a_12516_7093# a_38754_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24296 a_34434_65206# a_16746_65208# a_34342_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24297 a_34738_9858# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24298 a_10131_20175# a_7377_18012# a_9263_24501# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24299 VDD a_26319_38517# a_24892_38237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X243 a_5208_56989# a_4771_56597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2430 VDD a_8268_35381# a_7078_36103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X24300 a_27314_60186# a_12727_58255# a_27806_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24301 a_36442_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24302 a_11711_67325# a_10379_66389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24303 a_47486_64202# a_16746_64204# a_47394_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24304 a_3571_19126# a_3143_22364# a_3112_19319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24305 VSS a_12546_22351# a_44778_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24306 a_49494_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24307 a_24515_36965# a_23749_36929# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X24308 a_32730_60186# a_12981_59343# a_32334_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24309 a_32730_19898# a_12895_13967# a_32334_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2431 a_11335_10076# a_11140_10107# a_11645_9839# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X24310 VSS a_1586_21959# a_1591_23445# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24311 a_41967_31375# a_20359_29199# a_41878_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24312 VSS a_1916_33927# a_1867_32839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24313 a_12671_36367# a_12417_36694# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24314 a_20713_36929# a_20927_35877# a_21800_36165# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X24315 a_37446_56170# a_16746_56172# a_37354_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24316 a_38754_17890# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24317 a_43470_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24318 a_45782_18894# a_12899_10927# a_45386_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24319 VSS a_12727_13353# a_42770_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2432 a_22690_18894# a_12899_10927# a_22294_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24320 VSS a_2376_23047# a_2007_21237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24321 a_2656_70197# a_2824_70197# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24322 VSS a_17983_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24323 a_16928_42919# a_15959_42943# a_16891_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24324 a_2012_19631# a_1867_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24325 a_9869_49525# a_9651_49929# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24326 vcm_commonmode a_16362_62194# a_42466_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24327 a_18674_61190# a_12355_15055# a_18278_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24328 a_43378_58178# a_10515_22671# a_43870_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24329 vcm_commonmode VSS a_25398_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2433 VDD a_11711_12559# a_12174_12381# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X24330 VSS a_12877_14441# a_46786_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24331 a_43774_11866# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24332 a_1757_43029# a_1591_43029# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24333 a_32730_56170# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24334 VDD VDD a_37354_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24335 a_29322_18894# a_12895_13967# a_29814_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24336 a_26706_21906# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24337 VSS VSS a_29718_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24338 a_7800_54223# a_7764_53877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24339 a_41370_8854# a_12985_19087# a_41862_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2434 a_20682_9858# a_12985_19087# a_20286_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24340 a_1642_18231# a_1738_17973# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24341 a_7367_24527# a_5085_23047# a_7285_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24342 a_30326_13874# a_12727_15529# a_30818_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24343 a_1757_12565# a_1591_12565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24344 a_1644_62037# a_1591_59343# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24345 a_2834_23439# a_1757_23445# a_2672_23817# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24346 a_5087_24643# a_5085_24759# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24347 a_2107_44655# a_1591_44655# a_2012_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24348 a_20778_58500# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24349 VSS a_12899_11471# a_19678_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2435 vcm_commonmode VSS a_44474_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24350 a_17274_8854# a_12985_19087# a_17766_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24351 a_23694_14878# a_12727_15529# a_23298_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24352 a_23487_50095# a_23535_50247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24353 VSS a_10055_58791# a_20682_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24354 a_17366_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24355 a_32426_61190# a_16746_61192# a_32334_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24356 a_3104_25321# a_2315_24540# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24357 a_17300_51183# a_16385_51183# a_16953_51425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24358 a_27806_8456# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24359 a_23694_8854# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2436 a_10055_58791# a_9989_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X24360 a_24302_69222# a_12901_66959# a_24794_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24361 a_46482_9492# a_16746_9490# a_46390_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24362 a_35742_67214# a_12727_67753# a_35346_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24363 vcm_commonmode a_16362_63198# a_19374_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24364 a_8015_20175# a_7571_20291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X24365 VSS a_28195_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24366 a_11491_65327# a_11141_65327# a_11396_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24367 VSS a_18627_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24368 a_8059_74746# a_7901_74281# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24369 a_6607_13879# a_5959_13621# a_6841_14013# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2437 a_29718_24918# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24370 a_26495_38517# a_24893_37429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24371 a_48794_66210# a_12983_63151# a_48398_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24372 VDD a_10515_23975# a_46390_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24373 vcm_commonmode a_16362_16520# a_33430_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24374 VSS a_2847_44629# a_2781_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24375 a_18222_47507# a_18500_47491# a_18456_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24376 a_46390_64202# a_16362_64202# a_46482_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24377 a_11959_62973# a_11710_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24378 VDD a_12877_14441# a_36350_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24379 vcm_commonmode a_16362_69222# a_45478_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2438 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24380 a_11794_27791# a_11719_28023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24381 VDD a_4717_45985# a_4607_46109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24382 a_4395_53181# a_1823_53885# a_4032_53047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24383 a_33689_27791# a_15607_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24384 VDD a_2319_59317# a_2250_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24385 VDD a_12727_15529# a_49402_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24386 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24387 a_47486_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24388 a_31453_47919# a_26514_47375# a_31350_47919# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u w=650000u l=150000u
X24389 a_35263_28879# a_33839_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2439 a_37446_9492# a_16746_9490# a_37354_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24390 VDD a_4227_37887# a_4214_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24391 a_40762_61190# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24392 VSS a_31131_35281# a_31077_35307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24393 a_37354_66210# a_16362_66210# a_37446_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24394 a_13867_42134# a_13909_41923# a_13867_41807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24395 a_23694_71230# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24396 a_22386_69222# a_16746_69224# a_22294_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24397 vcm_commonmode a_16362_68218# a_49494_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24398 a_37846_11468# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24399 a_30722_72234# VDD a_30326_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X244 VSS a_10055_58791# a_29718_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2440 VDD a_4127_63669# a_2927_68565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24400 VDD a_17191_32117# a_16917_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24401 a_21290_24918# VSS a_21382_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24402 a_11141_65327# a_10975_65327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24403 a_41046_31055# a_34759_31029# a_40743_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24404 VDD a_2856_47753# a_3031_47679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24405 a_27406_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24406 VDD a_12056_55535# a_12231_55509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24407 vcm_commonmode a_16362_8488# a_25398_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24408 a_44778_60186# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24409 a_43470_58178# a_16746_58180# a_43378_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2441 a_41766_62194# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24410 a_4584_20407# a_3987_19623# a_4726_20214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24411 a_5504_37815# a_4314_40821# a_5735_37699# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24412 vcm_commonmode VSS a_40458_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24413 a_44778_19898# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24414 VDD a_15189_39889# a_15131_39997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24415 VDD a_35033_42044# a_34639_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24416 a_28056_43781# a_27183_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24417 a_27710_70226# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24418 a_26402_68218# a_16746_68220# a_26310_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24419 vcm_commonmode a_16362_65206# a_23390_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2442 a_6066_28309# a_2317_28892# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X24420 VSS a_9455_11079# a_9405_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24421 a_25306_23914# a_16362_23548# a_25398_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24422 VDD a_2008_28487# a_1683_27399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24423 VDD a_10975_66407# a_35346_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24424 a_9006_17277# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24425 VSS a_6514_37191# a_5701_37013# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X24426 a_17670_62194# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24427 VDD a_12355_65103# a_48398_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24428 a_45878_61512# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24429 VSS a_12727_58255# a_21686_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2443 a_31552_43781# a_30679_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X24430 VSS a_11067_67279# a_21686_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24431 VSS a_8933_22583# a_9135_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24432 a_29414_59182# a_16746_59184# a_29322_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24433 vcm_commonmode a_16362_56170# a_26402_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24434 VDD a_1586_9991# a_4075_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24435 VSS a_26319_37429# a_16152_37601# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24436 a_32334_71230# a_16362_71230# a_32426_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24437 a_35742_20902# a_11067_67279# a_35346_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24438 a_31726_15882# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24439 VDD a_12257_56623# a_38358_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2444 a_11909_51727# a_11855_51959# a_9240_53877# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X24440 a_18770_24520# a_18007_27441# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24441 a_22411_38007# a_21479_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24442 a_49402_72234# VDD a_49894_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24443 VDD a_11067_21583# a_22294_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24444 VSS a_23298_28487# a_23303_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24445 a_49894_60508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24446 a_1644_72373# a_1823_72381# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24447 a_29175_28335# a_28902_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24448 vcm_commonmode a_16362_22544# a_45478_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24449 VDD a_13643_28327# a_40233_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2445 a_38358_67214# a_16362_67214# a_38450_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24450 VSS a_22521_37692# a_22213_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24451 a_19282_20902# a_12985_7663# a_19774_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24452 a_3355_25071# a_3104_25321# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24453 a_26802_72556# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24454 a_34738_68218# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24455 a_19282_16886# a_16362_16520# a_19374_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24456 a_5226_48463# a_4149_48469# a_5064_48841# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24457 VDD a_12901_66665# a_30326_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24458 a_23390_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24459 a_20286_11866# a_16362_11500# a_20378_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2446 ctopp a_8583_33551# ctopp VSS sky130_fd_pr__nfet_01v8 ad=2.7645e+12p pd=2.191e+07u as=0p ps=0u w=1.9e+06u l=220000u M=2
X24460 VDD a_12981_59343# a_26310_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24461 a_47790_67214# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24462 VSS a_24515_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24463 a_38450_17524# a_16746_17522# a_38358_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24464 VDD a_51330_39932# a_52590_39198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X24465 VSS a_2011_34837# a_3707_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24466 VSS a_1923_59583# a_1881_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24467 a_22386_22544# a_16746_22542# a_22294_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24468 vcm_commonmode a_16362_21540# a_49494_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24469 VSS a_29791_52436# a_19720_55394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2447 VDD a_12981_59343# a_37354_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X24470 VDD a_10317_67191# a_10010_68021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X24471 a_26221_29423# a_26191_29397# a_25971_29789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24472 a_37750_59182# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24473 VSS a_33385_46805# a_29760_55394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X24474 VSS a_12257_56623# a_41766_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24475 a_35346_16886# a_12899_11471# a_35838_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24476 a_47486_72234# VDD a_47394_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24477 VSS a_12983_63151# a_24698_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24478 a_21686_64202# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24479 vcm_commonmode a_16362_13508# a_39454_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2448 a_10430_17277# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X24480 VDD a_2012_33927# a_2561_28918# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24481 a_48398_15882# a_12727_13353# a_48890_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24482 a_43470_11500# a_16746_11498# a_43378_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24483 a_8753_66103# a_7803_55509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24484 VDD a_12895_13967# a_42374_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24485 a_26402_21540# a_16746_21538# a_26310_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24486 a_2882_64605# a_2124_64507# a_2319_64476# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24487 a_26413_31055# a_26065_31171# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X24488 a_19500_40743# a_18627_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24489 a_5756_69135# a_5682_69367# a_5295_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2449 a_33338_55166# a_12869_2741# a_33830_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X24490 VDD a_2467_67668# a_2263_68218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X24491 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24492 VSS a_35033_38780# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24493 a_31726_56170# a_12257_56623# a_31330_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24494 a_25798_15484# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24495 VDD a_12899_10927# a_28318_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24496 a_13762_42895# a_13716_43047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24497 VDD a_34297_35516# a_33903_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24498 a_7567_64391# a_7445_63695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X24499 a_4149_45743# a_3983_45743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X245 a_1799_29556# a_27267_39605# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2450 VSS a_14049_36341# a_13983_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24500 a_13107_34789# a_12251_39069# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X24501 a_27563_35831# a_26631_35877# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24502 a_46882_69544# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24503 a_43378_66210# a_10975_66407# a_43870_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24504 a_29414_12504# a_16746_12502# a_29322_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24505 vcm_commonmode a_16362_60186# a_38450_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24506 VDD a_23747_31055# a_24746_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24507 a_12993_50345# a_6646_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24508 vcm_commonmode a_16362_19532# a_38450_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24509 VDD a_23447_28853# a_23298_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2451 VSS a_9529_28335# a_24768_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X24510 VDD a_35196_35425# a_34297_35516# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X24511 VSS a_10515_22671# a_18674_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24512 a_2559_24566# a_2223_28617# a_2100_24759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24513 a_29322_69222# a_16362_69222# a_29414_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24514 a_19743_41271# a_18811_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24515 VDD a_12039_69367# a_11943_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24516 VDD a_12985_19087# a_21290_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24517 a_26310_11866# a_10055_58791# a_26802_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24518 VDD a_3325_29967# a_4903_29975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24519 VDD a_12516_7093# a_23298_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2452 VSS a_5211_24759# a_5087_24643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X24520 a_20778_66532# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24521 a_47394_65206# a_12355_65103# a_47886_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24522 a_2467_67668# a_2559_67477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X24523 a_31009_39659# a_28099_42895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24524 VDD a_12727_58255# a_19282_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24525 VSS a_6752_29941# a_7089_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24526 a_28688_50247# a_29147_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24527 VSS a_6459_30511# a_11803_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24528 a_23390_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24529 a_20286_56170# a_16362_56170# a_20378_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2453 a_2203_44655# a_1757_44655# a_2107_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X24530 VDD a_1586_36727# a_1591_38677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24531 a_10575_69439# a_10400_69513# a_10754_69501# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24532 a_34738_21906# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24533 a_3983_30761# a_2216_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24534 a_9943_62607# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24535 vcm_commonmode a_16362_58178# a_32426_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24536 a_6683_37815# a_6377_38133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X24537 a_26671_50095# a_26155_50095# a_26576_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24538 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24539 a_37354_57174# a_12257_56623# a_37846_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2454 VDD a_9184_49159# a_7251_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24540 a_12157_68047# a_11053_69135# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24541 VSS a_6382_61127# a_6177_61127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24542 a_41862_55488# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24543 a_76082_40202# a_76178_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24544 a_47790_20902# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24545 a_2203_12937# a_1757_12565# a_2107_12937# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24546 VDD a_5993_32687# a_6651_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X24547 a_24794_65528# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24548 a_21290_62194# a_12355_15055# a_21782_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24549 VDD a_12947_8725# a_37354_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2455 a_20286_58178# a_10515_22671# a_20778_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24550 VSS a_12985_19087# a_33734_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24551 VSS a_12901_66665# a_45782_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24552 a_35039_51335# a_2959_47113# a_36097_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24553 a_24302_55166# VSS a_24394_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24554 VSS a_23051_28023# a_22991_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24555 a_37750_12870# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24556 a_23390_71230# a_16746_71232# a_23298_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24557 VSS a_6883_37019# a_6514_37191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24558 VSS a_12985_16367# a_41766_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24559 a_43774_8854# a_12947_8725# a_43378_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2456 a_18370_55166# VDD a_18278_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24560 a_2215_26525# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24561 a_27710_23914# a_10515_23975# a_27314_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24562 a_24302_14878# a_12877_14441# a_24794_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24563 VSS a_12985_7663# a_24698_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24564 a_2295_17429# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X24565 a_27806_56492# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24566 VSS a_2283_15797# a_3881_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24567 a_12671_42134# a_12713_41923# a_12671_41807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24568 a_8082_54599# a_7210_55081# a_8296_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24569 VSS a_12516_7093# a_49798_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2457 a_19678_16886# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24570 a_45478_65206# a_16746_65208# a_45386_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24571 a_17670_15882# a_12877_14441# a_17274_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24572 a_24716_31757# a_24632_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X24573 a_47486_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24574 VSS a_8827_17215# a_8761_17289# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24575 VSS a_12355_15055# a_39758_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24576 a_35438_57174# a_16746_57176# a_35346_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24577 a_2781_9839# a_1591_9839# a_2672_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24578 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X24579 a_36746_18894# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2458 a_19311_35823# a_19134_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24580 a_41462_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24581 a_43774_60186# a_12981_59343# a_43378_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24582 VSS a_12899_11471# a_40762_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24583 a_35346_8854# a_16362_8488# a_35438_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24584 a_43774_19898# a_12895_13967# a_43378_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24585 a_12257_56623# a_10055_58791# a_12269_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X24586 a_26706_70226# a_12901_66665# a_26310_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24587 a_18770_58500# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24588 a_8746_71443# a_9024_71427# a_8980_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24589 VSS a_3024_67191# a_9424_60949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2459 VDD a_6224_73095# a_7499_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X24590 VDD a_6473_40277# a_7107_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24591 VSS a_10055_58791# a_18674_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24592 a_45478_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24593 a_5683_18365# a_5535_18012# a_5320_18231# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24594 vcm_commonmode a_16362_17524# a_27406_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24595 a_40858_7452# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24596 a_5345_10927# a_5179_10927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24597 a_31422_15516# a_16746_15514# a_31330_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24598 vcm_commonmode a_16362_63198# a_40458_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24599 a_41370_59182# a_12901_58799# a_41862_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X246 a_42466_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2460 VSS a_18627_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X24600 a_35647_40229# a_33856_40743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X24601 a_16762_7452# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24602 VDD a_15345_34717# a_14951_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24603 a_22595_43177# a_21663_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24604 VSS a_5612_52520# a_5550_52637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24605 a_29718_61190# a_12355_15055# a_29322_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24606 a_30722_57174# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24607 a_14482_27497# a_11866_27791# a_14369_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24608 a_4985_69725# a_3325_69135# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X24609 VSS config_1_in[7] a_1591_4399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2461 VSS a_12877_14441# a_23694_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X24610 a_2126_16911# a_1591_16917# a_2040_17289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24611 VDD VDD a_26310_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24612 VSS VDD a_22690_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24613 a_11215_69679# a_10865_69679# a_11120_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24614 VDD VDD a_48398_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24615 a_5991_21263# a_5547_21379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X24616 VDD a_9863_51420# a_9794_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24617 vcm_commonmode a_16362_11500# a_32426_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24618 a_1895_71482# a_2322_72631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24619 a_42466_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2462 a_23685_50345# a_23631_50069# a_23487_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X24620 a_23749_36929# a_24055_36415# a_24987_36649# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X24621 VSS a_4852_23413# a_4798_23759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24622 VDD a_52778_39936# a_53378_39250# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24623 a_48490_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24624 a_31822_19500# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24625 VDD a_23685_29111# a_23447_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24626 a_30418_62194# a_16746_62196# a_30326_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24627 a_20009_48981# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X24628 VDD a_12546_22351# a_35346_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24629 vcm_commonmode a_16362_64202# a_44474_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2463 VDD a_6646_54135# a_7755_54999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24630 a_4031_50247# a_3325_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24631 VSS a_18662_43671# a_18667_43439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24632 a_7994_49917# a_2595_47653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24633 a_9333_72105# a_7925_72399# a_8539_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24634 VDD a_11067_67279# a_18278_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24635 a_33734_68218# a_12901_66959# a_33338_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24636 a_14088_39631# a_13837_39860# a_13867_39958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24637 a_18278_61190# a_16362_61190# a_18370_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24638 a_46786_67214# a_12727_67753# a_46390_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24639 VSS a_1923_59583# a_1881_59709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2464 a_20682_11866# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24640 vcm_commonmode a_16362_56170# a_34434_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24641 VSS a_32167_29611# a_25971_52263# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24642 vcm_commonmode a_16362_66210# a_17366_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24643 a_4151_28879# a_3707_28995# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X24644 VSS a_14963_39783# a_18949_39958# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24645 a_21382_64202# a_16746_64204# a_21290_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24646 a_2325_19873# a_2107_19631# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24647 a_19282_24918# VSS a_19374_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24648 a_24401_31171# a_2787_30503# a_24305_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24649 a_23390_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2465 a_17274_10862# a_16362_10496# a_17366_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X24650 a_36746_59182# a_12727_58255# a_36350_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24651 a_19374_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24652 a_31186_48169# a_26417_47919# a_31453_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u w=650000u l=150000u
X24653 a_2199_52271# a_1849_52271# a_2104_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24654 VDD a_12727_13353# a_34342_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24655 a_19678_69222# a_12516_7093# a_19282_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24656 a_1761_11471# a_1591_11471# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X24657 a_2944_59893# a_1591_59343# a_2872_59893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24658 a_10233_21379# a_10045_21379# a_10151_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24659 a_35438_10496# a_16746_10494# a_35346_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2466 a_33430_22544# a_16746_22542# a_33338_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24660 a_7676_61493# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24661 VSS a_5839_22351# a_6007_23145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24662 VSS a_2872_44111# a_19439_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X24663 VDD a_22259_48981# a_22246_49373# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24664 VDD a_23901_42044# a_23507_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24665 a_35346_67214# a_16362_67214# a_35438_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24666 VDD a_28446_31375# a_29926_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24667 VSS VSS a_37750_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24668 a_24394_7484# VDD a_24302_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24669 VDD a_12725_44527# a_27247_43047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2467 a_28881_52271# a_28423_52245# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X24670 VDD a_1586_45431# a_6559_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24671 a_30326_55166# VSS a_30818_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24672 a_21686_72234# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24673 a_9639_12015# a_9491_12297# a_9276_12167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24674 a_48398_66210# a_16362_66210# a_48490_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24675 a_4404_65327# a_4287_65540# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24676 a_1846_56875# a_2163_56765# a_2121_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24677 VDD a_10667_60735# a_10654_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24678 a_34342_9858# a_12546_22351# a_34834_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X24679 VSS a_4215_51157# a_23763_47381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2468 vcm_commonmode a_16362_61190# a_32426_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X24680 a_29718_15882# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2469 a_29035_38825# a_28103_38591# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X247 VDD a_4528_26159# a_7821_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2470 a_42866_24520# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2471 a_37520_49783# a_4351_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X2472 a_33734_10862# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2473 VDD a_14983_51157# a_17600_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.955e+12p ps=1.791e+07u w=1e+06u l=150000u M=4
X2474 a_27588_52271# a_8491_57487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2475 a_7161_19631# a_3247_20495# a_6743_19631# VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X2476 VSS a_23685_29111# a_25077_28129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2477 a_15681_27497# a_10964_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X2478 VDD a_12947_71576# a_27314_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2479 a_45478_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X248 a_28931_39679# a_28152_40517# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X2480 VSS a_30835_38695# a_13669_38517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2481 a_2325_29941# a_2107_30345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X2482 a_36336_36391# a_35463_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2483 VSS a_10975_66407# a_48794_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2484 a_20112_49551# a_19675_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2485 a_46882_23516# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2486 a_43378_20902# a_12985_7663# a_43870_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2487 a_43378_16886# a_16362_16520# a_43470_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2488 a_46482_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2489 VDD a_32121_40741# a_33668_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X249 VSS a_23395_32463# a_43623_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X2490 a_20672_51183# a_19946_51157# a_19502_51157# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X2491 a_76082_39738# a_76178_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2492 VSS a_23567_42035# a_23507_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2493 a_18674_63198# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2494 a_23830_49525# a_8531_70543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2495 VDD a_10975_66407# a_49402_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2496 VDD a_3799_20407# a_3799_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2497 a_75199_38962# a_75111_39506# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2498 a_38959_29967# a_37527_29397# a_16863_29415# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2499 a_49494_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X25 a_40366_20902# a_12985_7663# a_40858_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X250 a_42770_71230# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2500 a_42770_56170# a_12257_56623# a_42374_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2501 a_36842_15484# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2502 a_36746_21906# a_12985_7663# a_36350_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2503 a_30104_31849# a_28757_27247# a_14287_51175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=2
X2504 a_33338_72234# VSS a_33430_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2505 VDD a_12877_16911# a_40366_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2506 VSS a_4461_53113# a_4395_53181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2507 a_25702_66210# a_12983_63151# a_25306_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2508 VDD a_10515_22671# a_39362_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2509 a_11709_61217# a_11491_60975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X251 a_26523_28111# a_35907_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X2510 VDD a_14354_32117# a_14298_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X2511 VDD a_26433_39631# a_30007_38695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2512 a_49894_14480# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2513 a_49798_20902# a_11067_67279# a_49402_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2514 VDD a_10515_23975# a_23298_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2515 a_9865_14191# a_9275_15253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X2516 a_20778_20504# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2517 a_20378_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2518 a_47394_15882# a_16362_15516# a_47486_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2519 a_2834_10205# a_1757_9839# a_2672_9839# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X252 a_41462_69222# a_16746_69224# a_41370_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2520 VSS a_11067_23759# a_16362_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X2521 a_5159_43933# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X2522 a_23298_64202# a_16362_64202# a_23390_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2523 a_29679_37737# a_28747_37503# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2524 a_8485_29673# a_6649_25615# a_8485_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2525 a_3978_74183# a_4031_73095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X2526 result_out[0] a_1644_53877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2527 a_39758_12870# a_10055_58791# a_39362_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2528 VSS a_38436_29941# a_38380_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2529 vcm_commonmode a_16362_69222# a_22386_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X253 a_2629_64239# a_2250_64605# a_2557_64239# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2530 a_3305_38671# a_2847_38975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X2531 a_37354_11866# a_10055_58791# a_37846_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2532 VDD a_15607_46805# a_31481_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2533 vcm_commonmode a_16362_23548# a_46482_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2534 VDD a_3305_38671# a_5885_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X2535 VDD a_12727_15529# a_26310_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2536 a_3969_20175# a_3799_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2537 VSS a_36432_42919# a_36395_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2538 a_40218_27247# a_16863_29415# a_40049_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2539 a_24394_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X254 a_8297_31055# a_2235_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=0p ps=0u w=1e+06u l=150000u
X2540 VSS a_15681_27497# a_20685_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X2541 a_21290_12870# a_16362_12504# a_21382_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2542 a_20563_36649# a_20957_36604# a_20623_36595# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2543 a_6095_44807# a_7815_45503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X2544 a_27314_63198# a_16362_63198# a_27406_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2545 VDD a_12901_66959# a_47394_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2546 a_2557_56623# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2547 a_33071_51183# a_33041_51157# a_10687_52553# VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u M=2
X2548 a_48794_68218# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2549 a_4227_73791# a_4052_73865# a_4406_73853# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X255 a_2369_40303# a_2325_40545# a_2203_40303# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2550 vcm_commonmode a_16362_15516# a_36442_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2551 a_39454_18528# a_16746_18526# a_39362_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2552 VSS a_14681_50247# a_14511_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2553 a_7299_59663# a_6559_59663# a_7162_59575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2554 a_40458_13508# a_16746_13506# a_40366_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2555 a_13835_43177# a_27183_43493# a_28056_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X2556 a_2307_33231# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2557 VSS a_24893_37429# a_26495_38517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2558 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2559 VDD a_2899_16367# a_3301_16617# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X256 a_40366_24918# VSS a_40458_24552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2560 a_41232_28879# a_33641_29967# a_41141_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X2561 VDD a_2325_38645# a_2215_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2562 a_12580_15939# a_10055_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2563 a_26933_50095# a_26889_50337# a_26767_50095# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2564 a_27806_10464# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2565 VSS a_10515_22671# a_42770_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2566 VSS a_30609_49159# a_30485_49257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X2567 VDD a_3316_42313# a_3491_42239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2568 VSS a_12727_67753# a_25702_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2569 a_48890_64524# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X257 a_39854_21508# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2570 a_45386_61190# a_12981_59343# a_45878_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2571 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2572 a_8639_15113# a_8289_14741# a_8544_15101# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X2573 VSS a_26413_31055# a_27808_32459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X2574 a_6182_72943# a_6098_73095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X2575 VSS a_1586_69367# a_1591_71317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2576 a_8349_17277# a_8305_16885# a_8183_17289# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2577 a_9161_72737# a_7707_70741# a_9075_72737# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2578 vcm_commonmode a_16362_59182# a_29414_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2579 a_11396_65327# a_8999_61493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X258 VDD a_11803_55311# a_16746_66212# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X2580 a_36350_19898# a_11067_67279# a_36842_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2581 a_42165_36367# a_41999_36367# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2582 VSS a_12713_43011# a_19743_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2583 VDD a_4891_47388# a_27257_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2584 a_14831_50095# a_14445_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2585 a_37569_32143# a_27535_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2586 a_21479_34239# a_19596_34215# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X2587 a_38850_56492# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2588 a_33734_71230# a_12947_71576# a_33338_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2589 a_17613_30287# a_2235_30503# a_17554_30663# VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=2
X259 VSS a_4127_50069# a_4073_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X2590 a_18278_63198# a_12981_62313# a_18770_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2591 a_2834_45021# a_1757_44655# a_2672_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2592 VDD a_12355_65103# a_25306_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2593 a_22786_61512# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2594 a_11771_23671# a_11480_23957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2595 a_49402_60186# a_12727_58255# a_49894_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2596 VSS a_34482_29941# a_21187_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X2597 a_30418_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2598 a_17366_14512# a_16746_14510# a_17274_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2599 a_2721_55329# a_1591_54447# a_2635_55329# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X26 a_40366_16886# a_16362_16520# a_40458_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X260 a_39454_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2600 a_16746_65208# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X2601 a_11214_47919# a_2419_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X2602 a_37750_70226# a_12901_66665# a_37354_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2603 a_2325_12533# a_2107_12937# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X2604 a_8332_38377# a_6372_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.7e+11p pd=5.74e+06u as=0p ps=0u w=1e+06u l=150000u
X2605 a_21859_35831# a_20713_36929# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X2606 a_26802_60508# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2607 a_4149_48469# a_3983_48469# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2608 a_2107_40303# a_1757_40303# a_2012_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X2609 a_22921_52245# a_23193_52245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X261 a_36350_14878# a_16362_14512# a_36442_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2610 a_16746_14510# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X2611 a_40557_29451# a_32970_31145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2612 a_9161_30511# a_9204_30663# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X2613 a_14039_41271# a_13835_41001# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X2614 vcm_commonmode a_16362_22544# a_22386_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2615 a_8169_10749# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2616 a_31330_24918# VSS a_31822_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2617 a_28921_28879# a_28817_29111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2618 a_21290_57174# a_16362_57174# a_21382_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2619 VDD a_7265_56053# a_7201_56079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X262 VDD a_18016_46983# a_17311_46833# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2620 VSS a_12899_10927# a_37750_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2621 a_6895_15253# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2622 vcm_commonmode VSS a_47486_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2623 a_41766_15882# a_12877_14441# a_41370_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2624 a_5987_16733# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X2625 a_3307_18259# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X2626 a_19500_35303# a_18627_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2627 a_24698_67214# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2628 a_11320_16367# a_10405_16367# a_10973_16609# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X2629 a_9759_67869# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X263 a_40458_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2630 a_48794_21906# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2631 a_11049_18543# a_10883_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2632 a_14298_32143# a_12412_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X2633 VSS a_12546_22351# a_43774_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2634 a_9263_24501# a_4792_20443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X2635 a_7733_10749# a_7255_10357# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2636 a_32867_28879# a_32038_29575# a_32649_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2637 VSS a_2235_30503# a_16129_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2638 a_41462_62194# a_16746_62196# a_41370_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2639 a_42866_58500# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X264 a_46482_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2640 a_10589_12879# a_9491_12297# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X2641 a_38754_13874# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2642 a_24394_72234# VDD a_24302_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2643 a_45782_14878# a_12727_15529# a_45386_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2644 VSS a_10055_58791# a_42770_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2645 a_39454_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2646 a_2691_40847# a_2004_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X2647 a_7901_74281# a_7499_74031# a_7737_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X2648 a_9043_24527# a_9263_24501# a_9221_24847# VSS sky130_fd_pr__nfet_01v8 ad=5.07e+11p pd=5.46e+06u as=0p ps=0u w=650000u l=150000u
X2649 VSS a_12947_56817# a_31726_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X265 a_43378_60186# a_16362_60186# a_43470_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2650 a_30816_37253# a_29943_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2651 a_25306_15882# a_12727_13353# a_25798_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2652 a_28810_18496# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2653 VSS a_11067_21583# a_25702_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2654 a_28714_24918# VSS a_28318_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2655 VDD a_4067_15797# a_3998_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2656 a_33727_38825# a_32795_38591# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2657 a_3070_22717# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2658 a_11865_24527# a_7571_26151# a_11711_24847# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X2659 vcm_commonmode a_16362_12504# a_29414_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X266 a_10411_23759# a_9263_24501# a_10073_23439# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X2660 VSS a_41334_29575# a_41335_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2661 VSS a_20713_40193# a_22319_39913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2662 VSS a_4215_51157# a_27627_51733# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2663 a_18674_16886# a_12727_13353# a_18278_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2664 a_24643_28335# a_23685_29111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X2665 a_7183_49551# a_6559_49557# a_7075_49929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X2666 a_19525_28585# a_17222_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X2667 a_5169_13103# a_4429_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2668 a_12907_27023# a_40599_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2669 VSS a_25015_48437# a_24961_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X267 a_27267_39605# a_12641_37684# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2670 a_15211_50959# a_14983_51157# a_15074_50871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2671 a_9740_69501# a_9503_68841# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2672 VDD a_8082_54599# a_7313_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X2673 a_23790_69544# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2674 a_20286_66210# a_10975_66407# a_20778_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2675 inp_analog a_3339_43023# ctopp VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=0p ps=0u w=1.9e+06u l=220000u M=4
X2676 a_40366_8854# a_12985_19087# a_40858_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2677 a_10409_18543# a_9983_18870# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2678 a_18370_63198# a_16746_63200# a_18278_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2679 VDD a_7833_66415# a_7580_61751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X268 a_11299_62215# a_11395_62037# a_11697_62063# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X2680 a_19774_59504# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2681 a_4674_40277# a_5211_24759# a_7161_19631# VSS sky130_fd_pr__nfet_01v8 ad=9.035e+11p pd=9.28e+06u as=0p ps=0u w=650000u l=150000u M=4
X2682 VDD a_22448_37253# a_22352_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2683 VSS a_14293_39631# a_12889_39889# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2684 a_34738_8854# a_12947_8725# a_34342_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2685 a_10825_29688# a_6459_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.58e+11p pd=2.36e+06u as=0p ps=0u w=420000u l=150000u
X2686 VSS a_3031_47679# a_2959_47113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X2687 vcm_commonmode a_16362_18528# a_28410_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2688 a_32426_16520# a_16746_16518# a_32334_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2689 VDD a_32970_31145# a_34895_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X269 a_24302_56170# a_12947_56817# a_24794_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2690 a_32856_48463# a_32319_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X2691 a_2847_51157# a_1923_54591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2692 a_45478_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2693 a_2012_45565# a_1867_45743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2694 a_26802_8456# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2695 a_22690_8854# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2696 VSS a_6619_47607# a_5963_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2697 a_5612_52520# a_6985_52815# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X2698 a_24302_65206# a_12355_65103# a_24794_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2699 a_34943_51335# a_28881_52271# a_35183_51183# VSS sky130_fd_pr__nfet_01v8 ad=3.8025e+11p pd=3.77e+06u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X27 a_43470_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X270 a_33430_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2700 a_22352_42693# a_20897_42917# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X2701 a_45782_71230# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2702 a_31726_58178# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2703 a_44474_69222# a_16746_69224# a_44382_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2704 vcm_commonmode a_16362_66210# a_41462_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2705 a_1824_61127# a_1768_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X2706 VSS a_12985_19087# a_32730_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2707 a_43378_24918# VSS a_43470_24552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2708 a_34098_31849# a_33798_31145# a_34016_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2709 a_24698_20902# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X271 a_12340_29967# a_11803_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X2710 a_49494_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2711 a_46390_60186# a_16362_60186# a_46482_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2712 a_27314_56170# a_12947_56817# a_27806_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2713 a_36442_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2714 VSS a_12901_66665# a_22690_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2715 a_49798_70226# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2716 a_48490_68218# a_16746_68220# a_48398_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2717 VDD a_12985_16367# a_36350_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2718 vcm_commonmode a_16362_65206# a_45478_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2719 VDD a_10659_9813# a_9484_11989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X272 a_20754_37782# a_18127_35797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2720 a_17422_48829# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2721 a_20378_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2722 VDD a_12985_7663# a_19282_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2723 a_47394_23914# a_16362_23548# a_47486_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2724 VDD a_16744_41605# a_16648_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2725 a_11141_60975# a_10975_60975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2726 VDD a_12546_22351# a_49402_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2727 a_19885_50095# a_19715_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2728 a_39758_62194# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2729 vcm_commonmode a_16362_57174# a_35438_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X273 a_30534_49393# a_30525_49551# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2730 a_3297_53153# a_3231_53047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2731 VSS a_12727_58255# a_43774_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2732 a_8468_48841# a_7387_48469# a_8121_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X2733 a_40762_16886# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2734 VSS a_11067_67279# a_43774_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2735 vcm_commonmode a_16362_67214# a_18370_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2736 VDD a_1923_54591# a_2464_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2737 VSS a_16928_35303# a_16891_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2738 VSS a_12516_7093# a_26706_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2739 a_22386_65206# a_16746_65208# a_22294_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X274 a_5345_74031# a_5179_74031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2740 vcm_commonmode a_16362_56170# a_48490_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2741 a_18475_47158# a_12447_29199# a_18016_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X2742 VDD a_4341_62109# a_4441_62327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X2743 a_24394_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2744 a_21290_20902# a_16362_20536# a_21382_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2745 a_12792_51017# a_11877_50645# a_12445_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X2746 VSS a_10975_66407# a_12899_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X2747 a_9735_12342# a_9484_11989# a_9276_12167# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X2748 a_16640_51183# a_8132_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X2749 a_10351_12879# a_10317_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X275 a_26310_70226# a_16362_70226# a_26402_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2750 VDD a_12355_15055# a_44382_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2751 a_20682_60186# a_12981_59343# a_20286_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2752 a_9431_59887# a_9177_60214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2753 a_20682_19898# a_12895_13967# a_20286_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2754 a_22632_42919# a_21663_42943# a_22595_43177# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2755 VDD a_20635_29415# a_41697_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X2756 a_12473_42869# a_32187_40513# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2757 vcm_commonmode a_16362_8488# a_24394_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2758 VSS a_12981_59343# a_29718_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2759 a_25398_56170# a_16746_56172# a_25306_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X276 vcm_commonmode a_16362_65206# a_42466_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2760 a_26706_17890# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2761 a_2781_26159# a_1591_26159# a_2672_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2762 VDD a_9184_13255# a_7999_13083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2763 a_31422_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2764 VSS a_12727_13353# a_30722_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2765 VSS a_11035_47893# a_10969_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X2766 a_3714_56445# a_3668_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2767 VDD a_10257_56377# a_10287_56118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2768 a_36350_68218# a_16362_68218# a_36442_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2769 VDD VSS a_17274_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X277 VDD a_12985_16367# a_33338_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2770 VSS a_1923_54591# a_2369_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2771 VDD config_1_in[0] a_1591_8751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2772 a_48890_72556# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2773 a_11527_28701# a_10873_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X2774 VSS a_31096_38341# a_31059_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2775 result_out[11] a_1644_70197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2776 a_42374_11866# a_16362_11500# a_42466_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2777 a_53570_39250# a_52778_39198# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2778 VDD a_12981_59343# a_48398_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2779 a_34923_32375# a_30788_28487# a_35069_32463# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X278 a_18674_64202# a_12355_65103# a_18278_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2780 VDD a_23540_48981# a_23487_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X2781 vcm_commonmode a_16362_62194# a_30418_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2782 a_7917_13885# a_7917_12265# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X2783 a_31330_58178# a_10515_22671# a_31822_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2784 a_9390_51435# a_9668_51451# a_9624_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2785 a_29414_55166# VDD a_29322_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2786 VSS a_4151_28879# a_4351_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X2787 a_36264_30511# a_35815_31751# a_35959_30485# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X2788 a_31726_11866# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2789 a_28318_10862# a_16362_10496# a_28410_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X279 VDD a_12056_65327# a_12231_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2790 a_44474_22544# a_16746_22542# a_44382_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2791 a_18278_71230# a_12901_66665# a_18770_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2792 a_35601_27497# a_22015_28111# a_35529_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2793 a_18770_20504# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2794 VDD VDD a_25306_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2795 VSS a_12727_67753# a_33734_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2796 a_18370_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2797 VSS a_13669_39605# a_14088_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2798 VSS a_2419_48783# a_2511_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X2799 VSS a_4831_52413# a_4792_52539# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X28 VDD a_19807_28111# a_35079_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X280 a_44382_23914# a_16362_23548# a_44474_23548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2800 a_2387_47753# a_1941_47381# a_2291_47753# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X2801 a_7337_49917# a_7293_49525# a_7171_49929# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2802 VSS config_2_in[9] a_1591_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2803 VSS a_12983_63151# a_46786_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2804 a_43774_64202# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2805 VDD a_42188_37149# a_41289_36893# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X2806 VDD a_37534_51701# a_6467_55527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X2807 a_10679_74397# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X2808 a_41370_21906# a_11067_21583# a_41862_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2809 a_41370_17890# a_16362_17524# a_41462_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X281 VDD a_12546_22351# a_46390_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2810 a_7293_42721# a_7075_42479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X2811 a_10513_48161# a_10295_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X2812 VSS a_24331_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X2813 a_7622_61839# a_2952_66139# a_7812_61839# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X2814 a_19559_35561# a_13909_35395# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X2815 a_15959_36415# a_13097_35279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X2816 VDD a_6921_72943# a_4307_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X2817 VDD a_21829_48161# a_21719_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X2818 a_10216_67503# a_9135_67503# a_9869_67745# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X2819 a_48490_21540# a_16746_21538# a_48398_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X282 a_9971_23439# a_7841_22895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X2820 VSS a_12901_58799# a_36746_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2821 VDD a_6831_63303# a_26218_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X2822 a_19282_12870# a_16362_12504# a_19374_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2823 a_11902_27497# a_11711_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X2824 a_40762_57174# a_10515_22671# a_40366_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2825 VSS a_10515_63143# a_12539_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X2826 a_34834_16488# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2827 VSS a_12901_66959# a_19678_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2828 a_16746_22542# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X2829 a_23694_67214# a_12727_67753# a_23298_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X283 a_19374_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2830 VSS a_11067_13095# a_20682_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2831 a_4630_15823# a_3872_15939# a_4067_15797# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X2832 a_9468_53609# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2833 a_38450_13508# a_16746_13506# a_38358_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2834 vcm_commonmode a_16362_10496# a_35438_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2835 VSS a_9379_15039# a_9313_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X2836 a_47886_15484# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2837 a_19069_50613# a_18851_51017# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X2838 vcm_commonmode a_16362_20536# a_18370_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2839 a_21290_65206# a_16362_65206# a_21382_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X284 VDD a_12907_56399# a_16362_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X2840 a_4330_63827# a_4647_63937# a_4605_64061# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X2841 a_35838_9460# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2842 VDD a_9187_56597# a_9135_56623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X2843 a_2012_69501# a_1775_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2844 a_37750_55166# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2845 a_2107_12937# a_1757_12565# a_2012_12925# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X2846 a_2215_29967# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2847 VSS a_9705_11989# a_9639_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2848 a_5515_60137# a_5333_59343# a_5421_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X2849 a_18278_18894# a_16362_18528# a_18370_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X285 a_11522_23145# a_11574_22869# a_11067_47695# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X2850 vcm_commonmode a_16362_69222# a_33430_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 VDD a_12877_14441# a_24302_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2852 a_4341_62109# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2853 VSS a_2411_18517# a_8901_15101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2854 a_48398_11866# a_10055_58791# a_48890_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2855 a_38358_68218# a_12727_67753# a_38850_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2856 VDD a_12516_7093# a_45386_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2857 a_42866_66532# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2858 a_33338_9858# a_12546_22351# a_33830_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2859 a_37446_60186# a_16746_60188# a_37354_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X286 a_35237_52093# a_8531_70543# a_35165_52093# VSS sky130_fd_pr__nfet_01v8 ad=1.47e+11p pd=1.54e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2860 a_37446_19532# a_16746_19530# a_37354_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2861 a_17670_58178# a_12901_58799# a_17274_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2862 a_6662_33775# a_6372_38279# a_6662_34025# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X2863 a_42374_56170# a_16362_56170# a_42466_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2864 VSS a_2606_41079# a_8364_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2865 a_8157_58255# a_7107_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2866 a_28410_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2867 a_25306_66210# a_16362_66210# a_25398_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2868 a_25798_11468# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2869 a_26694_29473# a_2787_30503# a_26701_29739# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X287 a_20378_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2870 VDD a_32823_29397# a_36507_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2871 VDD a_7841_12167# a_9963_13760# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X2872 a_46882_65528# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2873 a_43378_62194# a_12355_15055# a_43870_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2874 a_7653_31599# a_7565_31751# a_7571_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2875 VSS a_38101_38565# a_39247_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2876 a_32273_40513# a_12357_37999# a_32187_40513# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X2877 VSS a_11067_21583# a_33734_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2878 a_32730_60186# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2879 a_49402_8854# a_12985_19087# a_49894_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X288 a_2292_17179# a_2295_17429# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X2880 a_31422_58178# a_16746_58180# a_31330_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2881 a_32730_19898# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2882 VDD a_24029_39355# a_36520_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X2883 VDD a_28708_52105# a_28883_52031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2884 a_10325_49929# a_9135_49557# a_10216_49929# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2885 a_11759_63927# a_11053_62607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2886 a_4893_33821# a_1915_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2887 a_36842_57496# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2888 VDD a_2830_15431# a_2781_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X2889 VSS a_11719_28023# a_14471_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X289 VDD a_11067_67279# a_29322_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2890 VDD VSS a_40366_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2891 VSS a_12985_7663# a_46786_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2892 a_31280_40517# a_30311_40229# a_31243_40183# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X2893 VDD a_12985_19087# a_20286_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2894 VDD a_4032_49159# a_2467_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2895 a_19774_67536# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2896 a_10717_53113# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2897 a_49894_56492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2898 VDD a_10975_66407# a_23298_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2899 a_20778_62516# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X29 a_20009_48981# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X290 VSS a_9955_20969# a_10521_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X2900 a_29322_24918# VSS a_29814_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2901 a_20672_51183# a_4758_45369# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X2902 a_2315_24540# a_2847_23743# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2903 a_44778_71230# a_12947_71576# a_44382_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2904 a_19282_57174# a_16362_57174# a_19374_57174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2905 VDD a_4227_37887# a_4685_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X2906 a_3523_13967# a_3843_13880# a_3677_13647# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2907 a_23390_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2908 a_26417_47919# a_25879_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2909 VSS a_12877_16911# a_36746_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X291 a_44778_68218# a_12901_66959# a_44382_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2910 VSS a_27250_27791# a_11067_46823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=5.6e+06u w=420000u l=150000u M=8
X2911 a_17891_43805# a_13005_43983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X2912 a_10515_23975# a_12815_6031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2913 a_10509_73193# a_9353_72399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2914 a_18811_34789# a_16928_36391# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X2915 a_32029_41829# a_32611_41317# a_33484_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X2916 a_25971_29423# a_2787_30503# a_26221_29423# VSS sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=2.7965e+11p ps=3.21e+06u w=420000u l=150000u
X2917 a_40762_10862# a_12546_22351# a_40366_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2918 a_5060_67753# a_5024_67885# a_4988_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2919 VSS a_10515_23975# a_19678_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X292 a_19678_72234# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2920 VSS a_7803_55509# a_7749_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2921 a_23790_14480# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2922 a_23694_20902# a_11067_67279# a_23298_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2923 VDD a_12257_56623# a_26310_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2924 a_48794_70226# a_12901_66665# a_48398_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2925 a_10288_17143# a_5535_18012# a_10430_17277# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X2926 a_11872_57711# a_10957_57711# a_11525_57953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X2927 a_7295_60751# a_6737_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2928 vcm_commonmode a_16362_17524# a_49494_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2929 VDD config_2_in[15] a_1591_52815# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X293 VDD a_4987_58229# a_4918_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X2930 vcm_commonmode a_16362_23548# a_20378_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2931 a_2847_23743# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2932 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2933 a_8173_70543# a_2686_70223# a_8531_70543# VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=9.035e+11p ps=9.28e+06u w=650000u l=150000u M=4
X2934 a_38754_62194# a_12981_62313# a_38358_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2935 a_24302_10862# a_12985_16367# a_24794_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2936 a_42770_8854# a_12947_8725# a_42374_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2937 a_36746_7850# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2938 VSS a_12895_13967# a_35742_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2939 VSS config_2_in[1] a_1591_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X294 a_3112_9527# a_1761_8751# a_3254_9661# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2940 vcm_commonmode a_16362_22544# a_33430_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2941 a_39836_38567# a_38867_38591# a_39799_38825# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X2942 VSS a_19780_41605# a_19743_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X2943 a_22436_51005# a_10503_52828# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2944 a_22690_68218# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2945 VDD a_12901_58799# a_17274_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2946 VSS a_36116_44765# a_35217_44509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X2947 a_3031_47679# a_2856_47753# a_3210_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X2948 a_28115_44535# a_27183_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X2949 a_17670_11866# a_12985_16367# a_17274_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X295 a_11067_23759# a_39331_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2950 a_7987_40821# a_7847_39872# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2951 VDD a_11760_46983# a_10407_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2952 a_9370_58575# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X2953 a_26402_17524# a_16746_17522# a_26310_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2954 a_2285_38155# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2955 a_9505_63401# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2956 a_20839_41001# a_21233_40956# a_19245_39747# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X2957 VSS a_15259_46805# a_12355_65103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X2958 a_10969_47919# a_9779_47919# a_10860_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2959 a_2375_29588# a_2467_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X296 VSS a_12516_7093# a_23694_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2960 a_3026_66415# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X2961 a_40858_59504# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2962 a_37354_70226# a_16362_70226# a_37446_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2963 VDD a_28089_31157# a_28446_31375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X2964 a_36746_14878# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2965 a_25702_59182# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2966 a_34342_8854# a_16362_8488# a_34434_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2967 a_23298_16886# a_12899_11471# a_23790_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2968 VDD a_40139_32143# a_35815_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X2969 a_4607_21085# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X297 a_49798_61190# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2970 a_12139_71829# a_11964_71855# a_12318_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X2971 vcm_commonmode a_16362_13508# a_27406_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2972 a_6786_37557# a_4314_40821# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2973 a_44474_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2974 a_31422_11500# a_16746_11498# a_31330_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2975 a_4312_19061# a_1586_18695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2976 a_5600_47919# a_4240_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X2977 VDD a_12895_13967# a_30326_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2978 a_4891_47388# a_5239_48767# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X2979 a_29718_58178# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 a_48490_59182# a_16746_59184# a_48398_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2980 a_36579_42359# a_35647_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2981 vcm_commonmode a_16362_66210# a_39454_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2982 a_29718_16886# a_12727_13353# a_29322_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2983 VSS a_2713_31353# a_2647_31421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2984 a_43470_64202# a_16746_64204# a_43378_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2985 a_4351_67279# a_7637_69679# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X2986 a_41510_29673# a_39727_27765# a_41418_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2987 a_33939_43439# a_33762_43439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2988 VSS a_4685_37583# a_6377_38133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X2989 VDD VDD a_25306_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X299 vcm_commonmode a_16362_56170# a_45478_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2990 VSS VDD a_21686_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2991 a_17366_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2992 a_11759_59575# a_11521_66567# a_11993_59709# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2993 a_31330_66210# a_10975_66407# a_31822_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2994 a_33430_56170# a_16746_56172# a_33338_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2995 a_34738_17890# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2996 a_29414_63198# a_16746_63200# a_29322_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2997 vcm_commonmode a_16362_60186# a_26402_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2998 vcm_commonmode VSS a_38450_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2999 vcm_commonmode a_16362_19532# a_26402_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3 a_30722_10862# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X30 VDD a_2787_32679# a_7544_32937# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X300 VSS a_1761_6031# a_1683_5059# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X3000 a_16362_66210# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3001 VSS a_5441_27791# a_7259_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X3002 a_31726_7850# VDD a_31330_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3003 VDD a_4717_48437# a_4607_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X3004 a_3295_62083# a_3983_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3005 a_18370_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3006 a_6676_69455# a_6921_72943# a_7449_69455# VSS sky130_fd_pr__nfet_01v8 ad=1.27725e+12p pd=1.303e+07u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X3007 a_37277_48169# a_20359_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3008 a_26221_29423# a_27234_29789# a_27422_29789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X3009 a_33668_39655# a_32795_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X301 a_2672_21807# a_1757_21807# a_2325_22049# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3010 a_43774_72234# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3011 VSS a_11395_62037# a_11341_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3012 a_35647_39141# a_33764_38567# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X3013 VDD a_2672_71689# a_2847_71615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3014 a_2122_19087# a_1945_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3015 a_5483_74244# a_2451_72373# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3016 a_9301_49557# a_9135_49557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3017 a_22690_21906# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3018 a_19282_20902# a_16362_20536# a_19374_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3019 VDD a_21948_34973# a_22352_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X302 a_21382_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3020 a_25306_57174# a_12257_56623# a_25798_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3021 a_23298_7850# VSS a_23390_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3022 a_34434_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3023 a_36746_55166# VSS a_36350_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3024 VSS VDD a_20682_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3025 a_19678_65206# a_10975_66407# a_19282_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3026 a_23987_39126# a_19629_39631# a_23915_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X3027 a_47486_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3028 result_out[12] a_1644_71829# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3029 VSS a_12727_13353# a_28714_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 a_5779_75093# a_5441_72399# a_5805_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3030 a_25702_12870# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3031 a_37750_63198# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3032 a_10949_72719# a_10615_72399# a_10865_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X3033 a_5625_37039# a_4887_36495# a_5537_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X3034 VSS a_12907_56399# a_16362_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X3035 VDD a_35815_31751# a_35615_30199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.25e+11p ps=2.85e+06u w=1e+06u l=150000u
X3036 VSS a_32887_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3037 a_4482_57863# a_22259_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3038 vcm_commonmode a_16362_57174# a_46482_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3039 a_23390_7484# VDD a_23298_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X304 vcm_commonmode a_16362_66210# a_28410_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3040 a_16824_28309# a_17278_28309# a_17216_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X3041 a_8189_27497# a_6773_27805# a_8117_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3042 a_77664_40024# a_75475_38962# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3043 a_25307_51549# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3044 a_35346_22910# a_10515_23975# a_35838_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3045 VDD a_10216_67503# a_10391_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3046 a_11212_57711# a_6417_62215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3047 a_29322_58178# a_10515_22671# a_29814_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3048 a_17711_32385# a_4191_33449# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3049 VDD a_10515_23975# a_42374_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X305 VDD a_10055_58791# a_19282_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3050 a_29718_11866# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3051 a_42374_64202# a_16362_64202# a_42466_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3052 VSS a_9260_25045# a_9481_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X3053 VSS a_12355_15055# a_27710_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3054 a_43870_9460# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3055 a_15775_42405# a_14919_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3056 a_31726_60186# a_12981_59343# a_31330_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3057 VDD a_12877_14441# a_32334_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3058 a_5918_27497# a_4248_29967# a_5795_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.65e+11p ps=2.93e+06u w=1e+06u l=150000u
X3059 a_31726_19898# a_12895_13967# a_31330_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X306 VSS a_8197_31599# a_14471_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3060 result_out[7] a_1644_63669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3061 a_39362_21906# a_11067_21583# a_39854_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3062 a_22922_30287# a_7862_34025# a_22753_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X3063 a_11803_55311# a_26267_43983# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3064 a_11619_56615# a_11067_46823# a_13051_46831# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X3065 VDD a_7221_43541# a_7251_43894# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3066 a_43378_70226# a_12516_7093# a_43870_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3067 a_39362_17890# a_16362_17524# a_39454_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3068 VDD a_12727_15529# a_45386_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3069 a_43470_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X307 a_17366_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3070 a_40366_12870# a_16362_12504# a_40458_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3071 a_5825_20495# a_5963_20149# a_5909_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3072 a_11141_60975# a_10975_60975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3073 VDD VSS a_28318_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3074 a_12713_28585# a_9179_22351# a_12631_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3075 VSS a_12901_66959# a_40762_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3076 a_2107_66415# a_1591_66415# a_2012_66415# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X3077 a_5497_63303# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X3078 a_1644_70197# a_1591_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3079 a_33830_11468# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X308 a_32426_64202# a_16746_64204# a_32334_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3080 VSS a_11067_13095# a_18674_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3081 a_10755_16367# a_10405_16367# a_10660_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X3082 a_42466_23548# a_16746_23546# a_42374_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3083 a_16270_72234# VDD a_16762_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3084 a_20778_70548# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3085 a_16362_17524# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X3086 a_46882_10464# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3087 a_19282_65206# a_16362_65206# a_19374_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3088 a_7838_38671# a_4685_37583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3089 a_24959_30503# a_34895_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X309 a_8219_56623# a_7210_55081# a_8082_56775# VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3090 VSS a_16152_37601# a_15253_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X3091 a_23390_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3092 a_20286_60186# a_16362_60186# a_20378_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3093 a_29814_20504# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3094 VSS a_12727_67753# a_44778_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3095 a_29414_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3096 a_17039_51157# a_19439_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3097 a_41766_65206# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3098 VSS a_13909_38659# a_26359_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X3099 a_30418_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X31 a_41596_29423# a_15607_46805# a_41335_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X310 VDD a_2672_69513# a_2847_69439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3100 a_29829_29673# a_28446_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X3101 VSS a_15459_41781# a_15271_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3102 a_10784_31599# a_9405_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3103 a_7812_57711# a_6559_59879# a_7622_57711# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=0p ps=0u w=650000u l=150000u
X3104 VDD a_5475_74895# a_5779_75093# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3105 a_10601_60809# a_9411_60437# a_10492_60809# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X3106 a_19774_12472# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3107 VSS a_2847_66389# a_2781_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X3108 VDD a_5915_30287# a_21101_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3109 a_28721_47081# a_20267_30503# a_13183_52047# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X311 a_37846_63520# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3110 a_17274_13874# a_16362_13508# a_17366_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3111 VDD a_12546_22351# a_23298_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3112 a_41211_28023# a_30052_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3113 vcm_commonmode a_16362_64202# a_32426_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3114 a_35602_34191# a_35425_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3115 a_1757_12565# a_1591_12565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3116 VSS a_19807_28111# a_35383_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3117 VSS a_6883_37019# a_8307_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3118 a_37354_63198# a_12981_62313# a_37846_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3119 a_35183_51183# a_2840_66103# a_35076_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u w=650000u l=150000u
X312 VDD a_5291_56765# a_5252_56891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3120 a_21686_68218# a_12901_66959# a_21290_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3121 VSS a_12901_58799# a_47790_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3122 a_41862_61512# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3123 VDD a_12663_40871# a_12651_41085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3124 VDD a_41289_43421# a_40895_43447# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3125 a_6996_53359# a_3016_60949# a_6516_53511# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3126 a_27314_9858# a_16362_9492# a_27406_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3127 a_36442_14512# a_16746_14510# a_36350_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3128 VDD a_6156_67477# a_6094_67825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.58e+11p ps=2.36e+06u w=420000u l=150000u
X3129 a_45878_16488# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X313 a_8761_17289# a_7571_16917# a_8652_17289# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X3130 a_9557_54991# a_7210_55081# a_9123_55223# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X3131 a_12651_39997# a_12663_39783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3132 a_12805_16911# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3133 a_4951_44330# a_5043_44085# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3134 VDD a_1923_59583# a_4127_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3135 a_7162_60039# a_7210_55081# a_7376_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X3136 vcm_commonmode a_16362_56170# a_22386_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3137 a_19374_24552# VDD a_19282_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3138 a_10931_53942# a_10680_54171# a_10472_54135# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X3139 VSS a_1586_9991# a_1591_9839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X314 VDD a_12355_15055# a_41370_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3140 VSS a_11067_23759# a_16362_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X3141 VDD a_33694_30761# a_42807_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X3142 VSS a_3339_43023# a_6614_21237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3143 a_49494_13508# a_16746_13506# a_49402_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3144 vcm_commonmode a_16362_10496# a_46482_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3145 VDD a_2143_15271# a_10873_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3146 a_25744_7638# a_20635_29415# a_37554_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X3147 VDD a_40323_29967# a_32823_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X3148 a_1757_69141# a_1591_69141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3149 VDD a_12983_63151# a_17274_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X315 a_40895_43447# a_41289_43421# a_39244_41953# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X3150 a_24698_59182# a_12727_58255# a_24302_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3151 a_31169_36395# a_26433_39631# a_31083_36395# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3152 VDD a_26523_29199# a_36350_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X3153 VDD a_4191_33449# a_21003_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3154 VDD a_8005_53333# a_2952_53333# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3155 a_30311_35877# a_29545_35841# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3156 a_9670_24527# a_9043_24527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3157 a_11304_71855# a_10969_71631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3158 a_36350_69222# a_12901_66959# a_36842_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3159 a_40858_67536# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X316 VSS a_4985_69725# a_5091_69685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3160 a_8219_56623# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3161 a_5975_16367# a_5529_16367# a_5879_16367# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X3162 a_12985_7663# a_12815_7663# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3163 a_40366_57174# a_16362_57174# a_40458_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3164 a_3254_19453# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3165 VDD a_12473_37429# a_12417_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3166 a_18770_62516# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3167 a_28714_58178# a_12901_58799# a_28318_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3168 a_23298_67214# a_16362_67214# a_23390_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3169 VDD a_12981_59343# a_22294_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X317 a_24638_49871# a_6835_46823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X3170 VSS VSS a_25702_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3171 a_18811_39141# a_18045_39105# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X3172 a_48890_7452# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3173 a_44778_7850# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3174 VSS a_10515_23975# a_40762_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3175 VSS a_21948_34973# a_21049_34717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X3176 a_37446_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3177 a_6752_29941# a_4248_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3178 a_18084_28111# a_13390_29575# a_17964_28111# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X3179 a_6666_53359# a_3668_56311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 VDD a_7939_30503# a_27323_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3180 VDD a_2327_54135# a_2327_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3181 VSS a_12546_22351# a_37750_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3182 a_20612_37607# a_14293_37455# a_20754_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3183 VDD a_5239_65301# a_5682_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3184 VDD a_6435_47893# a_6559_22671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X3185 a_33734_17890# a_12899_11471# a_33338_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3186 a_3843_13880# a_2873_13879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3187 a_36671_39913# a_36708_39655# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X3188 VDD a_4952_68279# a_4211_67655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3189 a_43470_72234# VDD a_43378_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X319 a_9179_22351# a_8671_22671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.35e+11p pd=2.67e+06u as=0p ps=0u w=1e+06u l=150000u
X3190 a_32401_49871# a_27869_50095# a_32134_49159# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3191 a_30418_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3192 VDD a_1586_51335# a_1683_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3193 a_47790_24918# VSS a_47394_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3194 a_44382_15882# a_12727_13353# a_44874_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3195 VSS a_11067_21583# a_44778_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3196 a_7213_62215# a_7107_65871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3197 a_47886_57496# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3198 VDD a_75475_40594# a_76180_40594# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3199 VSS a_2927_39733# a_1895_38842# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X32 VDD a_10975_66407# a_46390_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X320 a_38450_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3200 a_17274_58178# a_16362_58178# a_17366_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3201 a_31822_23516# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3202 a_31422_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3203 VSS a_29667_31055# a_30203_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3204 VSS a_6095_44807# a_11345_53359# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3205 VSS a_6625_29941# a_6039_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X3206 a_15064_27907# a_14471_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3207 a_37750_16886# a_12727_13353# a_37354_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3208 VSS a_12727_15529# a_34738_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3209 VSS a_2143_15271# a_10883_11177# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X321 VSS a_12981_59343# a_26706_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3210 a_20897_42917# a_21479_42405# a_22352_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3211 VDD a_4758_45369# a_19894_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3212 VDD a_8121_48437# a_8011_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X3213 a_2345_33749# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3214 a_17274_17890# a_12899_10927# a_17766_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3215 VSS a_12947_23413# a_17670_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3216 a_2007_39978# a_2052_38377# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3217 VSS a_12877_16911# a_47790_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3218 a_21782_15484# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3219 a_21686_21906# a_12985_7663# a_21290_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X322 a_22386_56170# a_16746_56172# a_22294_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3220 a_20635_27247# a_10873_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X3221 a_9431_60214# a_6559_59879# a_9431_59887# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X3222 VDD a_26319_41781# a_13576_42589# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3223 a_9313_15113# a_8123_14741# a_9204_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X3224 a_22230_32259# a_20905_32143# a_22148_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3225 VDD a_10515_22671# a_24302_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3226 VSS a_4495_35925# a_6883_37019# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3227 VDD a_26350_28585# a_26523_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X3228 vcm_commonmode a_16362_60186# a_34434_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3229 vcm_commonmode a_16362_19532# a_34434_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 a_23694_17890# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3230 a_38850_59504# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3231 a_32334_15882# a_16362_15516# a_32426_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3232 VSS a_1761_52815# a_30591_37455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3233 vcm_commonmode a_16362_70226# a_17366_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3234 a_4157_32259# a_1915_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3235 a_19069_50613# a_18851_51017# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X3236 VSS a_11067_13095# a_12727_13353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X3237 vcm_commonmode a_16362_18528# a_47486_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3238 a_6069_30761# a_6039_30663# a_5997_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3239 VSS a_37076_37253# a_37039_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X324 vcm_commonmode VSS a_49494_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3240 a_41872_29423# a_41335_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X3241 a_7444_34025# a_5691_36727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3242 a_24698_12870# a_10055_58791# a_24302_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3243 a_36746_63198# a_15439_49525# a_36350_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3244 a_8424_58255# a_7773_63927# a_7963_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X3245 a_22690_9858# a_12985_19087# a_22294_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3246 a_12024_30199# a_11710_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3247 a_2177_53359# a_1899_53387# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3248 a_22294_11866# a_10055_58791# a_22786_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3249 VSS a_2787_30503# a_26191_29397# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X325 a_13984_43781# a_13015_43493# a_13947_43447# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X3250 a_16648_41605# a_15775_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3251 vcm_commonmode a_16362_23548# a_31422_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3252 VDD a_38784_42589# a_39372_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X3253 a_39454_9492# a_16746_9490# a_39362_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3254 a_49798_62194# a_12981_62313# a_49402_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3255 a_13743_35836# a_18811_34789# a_19743_34743# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X3256 a_19715_52271# a_19478_51959# a_19621_52271# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X3257 a_33430_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3258 a_3521_57283# a_1591_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X3259 a_33734_68218# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X326 a_30722_18894# a_12899_10927# a_30326_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3260 a_23626_31573# a_22151_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3261 a_1823_54973# a_2847_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3262 a_9513_65301# a_11521_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3263 VDD a_38784_42589# a_37885_42333# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X3264 VDD a_12901_58799# a_28318_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3265 vcm_commonmode a_16362_15516# a_21382_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3266 a_24394_18528# a_16746_18526# a_24302_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3267 VDD a_11067_21583# a_34342_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3268 a_4149_24527# a_3801_24643# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3269 VSS a_12473_37429# a_12417_37782# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X327 VSS a_51714_39886# a_51330_39932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X3270 a_28714_11866# a_12985_16367# a_28318_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3271 VDD a_26433_39631# a_30835_38695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3272 a_4528_62069# a_4341_62109# a_4441_62327# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X3273 a_8377_39465# a_7948_38377# a_8304_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.281e+11p pd=1.45e+06u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X3274 a_9217_29423# a_9367_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X3275 a_48398_70226# a_16362_70226# a_48490_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3276 VSS a_12901_66665# a_41766_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3277 a_29322_66210# a_10975_66407# a_29814_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3278 a_7571_26151# a_11035_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3279 a_3145_34319# a_2216_28309# a_3063_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X328 VDD a_7862_34025# a_20103_30287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3280 a_6818_50959# a_6795_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X3281 a_30326_61190# a_12981_59343# a_30818_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3282 VDD a_17311_46833# a_17171_46859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3283 vcm_commonmode a_16362_14512# a_25398_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3284 VDD a_12985_7663# a_38358_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3285 VSS a_41289_36893# a_40981_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3286 a_35438_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3287 VDD a_9275_15253# a_7987_15431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3288 VSS a_23193_52245# a_22951_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X3289 VDD a_6637_20407# a_4839_21495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X329 VSS a_8636_63669# a_7891_64213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X3290 a_32611_41317# a_31004_40743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3291 a_38358_62194# a_16362_62194# a_38450_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3292 a_21290_19898# a_11067_67279# a_21782_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3293 a_42466_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3294 a_23790_56492# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3295 VDD a_22084_49007# a_22259_48981# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3296 a_7019_50639# a_6795_51157# a_6646_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u M=2
X3297 a_25398_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3298 vcm_commonmode a_16362_67214# a_37446_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3299 VSS a_39449_39868# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X33 a_5098_41391# a_4960_40847# a_5098_41641# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X330 a_33486_34191# a_33309_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3300 ctopp a_3339_43023# ctopp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u M=2
X3301 a_27183_34789# a_23567_35507# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3302 a_41462_65206# a_16746_65208# a_41370_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3303 a_4685_37583# a_4227_37887# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X3304 a_40366_20902# a_16362_20536# a_40458_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3305 a_43470_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3306 a_30845_51727# a_29361_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X3307 a_8271_74953# a_7755_74581# a_8176_74941# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X3308 a_39454_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3309 VDD a_76365_40202# a_76178_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X331 a_2307_33231# a_1683_33237# a_2199_33609# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3310 VSS a_4495_35925# a_9135_27023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3311 VSS a_22132_44129# a_21233_44220# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X3312 a_41159_28585# a_28817_29111# a_41261_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3313 a_36328_49525# a_34145_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X3314 VDD a_37761_44759# a_37706_44135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3315 vcm_commonmode a_16362_8488# a_18370_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3316 VSS a_32143_35281# a_32089_35307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3317 VSS a_1586_69367# a_4719_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3318 VSS a_2099_59861# a_2511_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3319 VSS VDD a_18674_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X332 a_7807_69455# a_7571_68047# a_4307_67477# VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X3320 a_1915_51946# a_2007_51701# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3321 a_10651_17277# a_5671_21495# a_10288_17143# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3322 VSS a_9240_53877# a_9186_54223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3323 VDD a_22151_29941# a_20946_30669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3324 a_22690_70226# a_12901_66665# a_22294_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3325 VSS a_12981_59343# a_48794_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3326 a_44474_56170# a_16746_56172# a_44382_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3327 a_45782_17890# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3328 a_1881_64239# a_1846_64491# a_1643_64213# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3329 a_19807_27247# a_20027_27221# a_19889_27497# VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X333 VDD a_35616_27765# a_35550_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3330 a_27406_66210# a_16746_66212# a_27314_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3331 VSS a_27393_47919# a_28524_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3332 a_12967_50943# a_12792_51017# a_13146_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3333 a_29414_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3334 a_26310_21906# a_16362_21540# a_26402_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3335 VDD a_15439_49525# a_36350_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3336 a_5363_25321# a_4149_24527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3337 a_76346_40594# a_76180_40594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3338 VSS a_35647_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3339 a_7126_65693# a_7000_65595# a_6722_65579# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X334 a_46390_67214# a_16362_67214# a_46482_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3340 a_25702_61190# a_12355_15055# a_25306_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3341 VSS a_12899_10927# a_22690_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3342 VDD a_10964_25615# a_16865_27511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3343 a_49798_16886# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3344 vcm_commonmode VSS a_32426_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3345 a_5913_48161# a_5695_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X3346 a_47394_10862# a_16362_10496# a_47486_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3347 VSS a_15775_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3348 a_37354_71230# a_12901_66665# a_37846_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3349 a_33734_21906# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X335 VDD a_12981_59343# a_45386_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3350 a_17422_48502# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3351 a_36579_41271# a_35647_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3352 a_14445_50095# a_14511_50069# a_14291_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X3353 a_5529_16367# a_5363_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3354 a_9637_30511# a_9161_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.34e+11p pd=2.02e+06u as=0p ps=0u w=650000u l=150000u
X3355 a_45478_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3356 a_15829_30287# a_15799_29941# a_15745_30287# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3357 a_27535_30503# a_37287_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3358 a_9626_61635# a_9526_61751# a_9544_61635# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3359 a_30757_37455# a_30591_37455# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X336 a_18285_30511# a_14926_31849# a_7295_44647# VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=1.105e+12p ps=1.12e+07u w=650000u l=150000u M=4
X3360 a_4529_40553# a_1689_10396# a_4446_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X3361 VSS a_4035_11989# a_3983_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3362 VSS a_12899_11471# a_26706_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3363 a_23694_13874# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3364 VDD a_31741_30485# a_30891_28309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3365 a_30722_14878# a_12727_15529# a_30326_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3366 a_24394_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3367 a_35438_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3368 a_48794_63198# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3369 a_25493_29967# a_25145_30083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X337 a_26402_55166# VDD a_26310_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3370 VSS a_12901_66959# a_38754_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3371 a_35742_66210# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3372 a_42770_67214# a_12727_67753# a_42374_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3373 a_27314_59182# a_12901_58799# a_27806_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3374 VDD a_2592_43023# a_3162_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3375 a_2583_68047# a_1959_68053# a_2475_68425# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3376 a_4443_36611# a_3305_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X3377 a_3325_49551# a_2847_49855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3378 VSS a_12489_47919# a_10515_63143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X3379 VSS a_12039_69367# a_11985_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X338 a_27710_16886# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3380 vcm_commonmode a_16362_20536# a_37446_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3381 a_32371_32117# a_31964_30485# a_32589_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X3382 a_40366_65206# a_16362_65206# a_40458_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3383 a_46390_22910# a_10515_23975# a_46882_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3384 a_2656_42301# a_2539_42106# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X3385 VSS a_20899_44211# a_20839_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X3386 a_18770_70548# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3387 a_39454_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3388 a_36350_55166# VSS a_36442_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3389 a_32730_59182# a_12727_58255# a_32334_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X339 VSS a_1586_18695# a_10883_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3390 VSS a_12981_62313# a_25702_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3391 a_35438_71230# a_16746_71232# a_35346_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3392 a_2203_69513# a_1757_69141# a_2107_69513# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X3393 VSS a_6821_26311# a_6773_27805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3394 a_39758_65206# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3395 a_39854_17492# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3396 a_39758_23914# a_10515_23975# a_39362_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3397 a_36350_14878# a_12877_14441# a_36842_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3398 a_28410_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3399 a_16441_41781# a_15459_41781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X34 a_28714_62194# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X340 a_12546_22351# a_10515_22671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X3400 VDD a_12877_14441# a_43378_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3401 a_40858_12472# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3402 a_37354_18894# a_16362_18528# a_37446_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3403 VSS a_12869_2741# a_33734_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X3404 VDD a_4960_40847# a_5098_41641# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3405 a_39454_70226# a_16746_70228# a_39362_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3406 a_30418_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3407 a_12283_42359# a_12343_42333# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X3408 a_12899_2767# a_12869_2741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3409 a_40458_24552# VDD a_40366_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X341 VSS a_2375_13268# a_1895_12730# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3410 a_24201_39126# a_24029_39355# a_23987_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3411 a_44382_66210# a_16362_66210# a_44474_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3412 a_16746_60188# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3413 VDD a_1925_18231# a_1738_17973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3414 VSS a_4528_26159# a_7841_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=2
X3415 a_3026_15101# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X3416 a_30722_71230# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3417 a_44874_11468# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3418 a_33264_37601# a_32795_38053# a_33668_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3419 a_14031_38007# a_13909_37571# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X342 VSS a_12877_14441# a_31726_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3420 VSS a_11067_13095# a_29718_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3421 a_33784_50101# a_33597_50141# a_33697_50359# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X3422 a_34834_68540# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3423 a_27806_21508# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3424 a_6435_47893# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3425 a_27406_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3426 a_1757_19631# a_1591_19631# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3427 a_1586_36727# a_4035_33205# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X3428 VDD a_10475_14165# a_9083_13879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3429 a_31330_60186# a_16362_60186# a_31422_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X343 VDD a_13484_39325# a_12585_39069# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X3430 VSS a_12947_56817# a_19678_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3431 a_3763_10761# a_3247_10389# a_3668_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X3432 a_3529_25731# a_3578_25625# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X3433 a_21382_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3434 a_17766_13476# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3435 VDD a_4891_47388# a_23847_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3436 VDD a_12985_16367# a_21290_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3437 vcm_commonmode a_16362_65206# a_30418_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3438 a_38850_67536# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3439 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X344 a_25306_10862# a_16362_10496# a_25398_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3440 a_35346_64202# a_11067_13095# a_35838_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3441 a_32334_23914# a_16362_23548# a_32426_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3442 a_15775_41317# a_13097_40719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3443 VDD a_10975_66407# a_42374_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3444 a_28318_13874# a_16362_13508# a_28410_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3445 a_48398_63198# a_12981_62313# a_48890_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3446 a_24698_62194# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3447 a_3247_20495# a_5052_14709# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u M=4
X3448 vcm_commonmode a_16362_57174# a_20378_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3449 VDD a_12189_46805# a_12219_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X345 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3450 a_47486_14512# a_16746_14510# a_47394_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3451 a_17589_30761# a_17554_30663# a_17507_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=1.87e+12p ps=1.774e+07u w=1e+06u l=150000u
X3452 a_10471_65002# a_10501_65871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3453 VDD a_10515_22671# a_32334_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3454 a_35932_38689# a_35647_39141# a_36579_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3455 VSS a_10515_23975# a_38754_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3456 vcm_commonmode a_16362_56170# a_33430_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3457 a_42770_20902# a_11067_67279# a_42374_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3458 VDD a_27901_52513# a_27791_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X3459 VDD a_5098_41641# a_5039_42167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X346 a_41462_22544# a_16746_22542# a_41370_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3460 VDD a_5239_20693# a_5226_21085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3461 a_11320_16367# a_10239_16367# a_10973_16609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X3462 VDD a_12257_56623# a_45386_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3463 VSS a_12251_39069# a_12191_39095# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X3464 VSS a_9972_69831# a_9314_69367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3465 VDD a_10665_58487# a_10478_58229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3466 VSS a_22448_38341# a_22411_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X3467 a_42374_8854# a_12985_19087# a_42866_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3468 a_7267_27497# a_4427_30511# a_7195_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3469 VDD a_12983_63151# a_28318_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X347 a_36350_59182# a_16362_59182# a_36442_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3470 a_25798_63520# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3471 VSS a_3123_53047# a_2559_52789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3472 VSS a_1923_73087# a_2737_68413# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3473 a_32730_12870# a_10055_58791# a_32334_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3474 VSS a_5671_21495# a_10338_19631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3475 a_28410_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3476 a_9278_57487# a_7155_55509# a_9468_57487# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X3477 a_33856_42693# a_32887_42405# a_33819_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3478 a_36746_8854# a_12947_8725# a_36350_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3479 VSS a_1642_22583# a_1591_22351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X348 a_5879_16367# a_5363_16367# a_5784_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X3480 VDD a_2959_47113# a_30845_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3481 VDD a_5211_24759# a_9551_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3482 a_2847_18517# a_2411_18517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3483 a_21290_68218# a_16362_68218# a_21382_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3484 VSS a_6467_55527# a_7299_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3485 a_17763_35797# a_17939_36129# a_17891_36189# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X3486 a_28810_8456# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3487 a_24698_8854# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3488 VDD a_27415_36341# a_27239_36341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X3489 a_29814_62516# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X349 a_2503_34319# a_2473_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3490 VDD a_8753_19319# a_8104_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X3491 a_35438_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3492 VSS config_2_in[7] a_1591_40847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3493 a_10515_23975# a_12815_6031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3494 VSS a_2689_65103# a_6721_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X3495 VDD a_22989_48437# a_23685_50345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3496 a_11297_49257# a_7000_43541# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.36e+12p pd=1.272e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X3497 a_5905_57961# a_1823_65853# a_5823_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X3498 VDD a_5052_14709# a_3247_20495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X3499 VSS a_15683_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X35 a_46482_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X350 a_8773_63695# a_4339_64521# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X3500 a_15871_27247# a_11430_26159# a_15681_27497# VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X3501 VSS a_1952_60431# a_2813_56417# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3502 a_38013_47919# a_20359_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3503 VSS config_1_in[0] a_1591_8751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3504 a_3291_22717# a_3143_22364# a_2928_22583# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X3505 a_44778_59182# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3506 a_4311_58229# a_4514_58387# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3507 a_19520_52047# a_19478_51959# a_19217_51701# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3508 a_38754_24918# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3509 a_21371_52263# a_30790_30663# a_30748_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X351 a_19807_28111# a_32319_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X3510 VSS a_32823_29397# a_39771_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X3511 a_2742_42997# a_2592_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X3512 a_44778_17890# a_12899_11471# a_44382_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3513 a_42374_16886# a_12899_11471# a_42866_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3514 a_13716_43047# a_33015_40513# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3515 VDD a_3751_72373# a_2747_72007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3516 a_27710_69222# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3517 VSS a_12983_63151# a_31726_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3518 a_6251_15279# a_5805_15279# a_6155_15279# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X3519 VDD a_32029_38565# a_33484_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X352 a_18756_51005# a_6559_59879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3520 a_33430_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3521 vcm_commonmode a_16362_23548# a_29414_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3522 vcm_commonmode a_16362_61190# a_41462_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3523 VSS a_12120_29941# a_12064_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3524 a_35382_51157# a_35061_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3525 a_28318_58178# a_16362_58178# a_28410_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3526 VSS a_12677_40157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3527 VSS a_12901_58799# a_21686_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3528 a_12757_9295# a_12479_9633# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3529 a_5915_30287# a_14679_31288# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X353 VDD VDD a_22294_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3530 a_48794_16886# a_12727_13353# a_48398_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3531 VSS a_12727_15529# a_45782_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3532 a_28756_55394# a_22843_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X3533 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3534 vcm_commonmode a_16362_15516# a_19374_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3535 a_15103_49525# a_15439_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3536 VDD a_12947_71576# a_36350_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3537 a_28318_17890# a_12899_10927# a_28810_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3538 VDD VDD a_19282_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3539 a_23390_13508# a_16746_13506# a_23298_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X354 a_40458_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3540 vcm_commonmode a_16362_10496# a_20378_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3541 a_31330_7850# VDD a_31822_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3542 a_32826_15484# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3543 a_36890_34191# a_36713_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3544 a_36442_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3545 a_5087_72512# a_3751_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X3546 VDD a_2748_68565# result_out[10] VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3547 a_48490_63198# a_16746_63200# a_48398_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3548 a_19374_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3549 vcm_commonmode a_16362_60186# a_45478_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X355 a_2295_31599# a_1849_31599# a_2199_31599# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X3550 a_3704_61839# a_3016_60949# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3551 a_49894_59504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3552 vcm_commonmode a_16362_19532# a_45478_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3553 a_22690_55166# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3554 VDD a_23395_32463# a_43455_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X3555 vcm_commonmode a_16362_70226# a_28410_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3556 VDD a_10239_16911# a_10423_17455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3557 a_7102_39465# a_7244_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X3558 a_1952_60431# a_1775_60439# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3559 VSS a_2319_73180# a_2250_73309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X356 VDD a_12981_62313# a_18278_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3560 a_34342_21906# a_16362_21540# a_34434_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3561 a_6725_49557# a_6559_49557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3562 VSS a_2411_18517# a_2369_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3563 a_4761_20719# a_4717_20961# a_4595_20719# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3564 a_33338_11866# a_10055_58791# a_33830_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3565 a_30005_48463# a_29651_48576# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3566 a_19282_19898# a_11067_67279# a_19774_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3567 a_24067_42583# a_14258_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3568 a_23298_68218# a_12727_67753# a_23790_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3569 a_34738_66210# a_12983_63151# a_34342_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X357 a_25019_47679# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3570 vcm_commonmode a_16362_62194# a_18370_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3571 a_2284_36103# a_2473_34293# a_2426_35951# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X3572 VDD a_28883_52031# a_29361_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3573 VDD a_12516_7093# a_30326_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3574 a_11872_57711# a_10791_57711# a_11525_57953# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X3575 a_12989_31421# a_12935_31287# a_12883_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3576 a_22386_60186# a_16746_60188# a_22294_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3577 a_22386_19532# a_16746_19530# a_22294_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3578 VDD a_12727_58255# a_26310_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3579 VDD a_17763_43413# a_17711_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X358 VDD a_3843_13880# a_3801_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X3580 a_11943_69367# a_12135_69109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3581 a_25447_34743# a_24515_34789# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3582 a_44382_57174# a_12257_56623# a_44874_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3583 VDD a_32823_29397# a_33689_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.95e+11p ps=5.19e+06u w=1e+06u l=150000u
X3584 a_27314_67214# a_12983_63151# a_27806_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3585 a_7293_42721# a_7075_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3586 a_38754_65206# a_10975_66407# a_38358_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3587 a_31822_65528# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3588 VSS a_2847_15039# a_2781_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X3589 a_20741_41605# a_21049_41245# a_20715_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X359 a_39758_69222# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3590 a_30790_30663# a_4811_34855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3591 a_36350_63198# a_16362_63198# a_36442_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3592 a_44778_12870# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3593 a_6177_61127# a_2952_66139# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3594 VDD a_12985_7663# a_49402_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3595 a_21782_57496# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3596 a_27710_22910# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3597 vcm_commonmode a_16362_68218# a_35438_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3598 a_17366_7484# VDD a_17274_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3599 VSS a_12985_7663# a_31726_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 VDD a_11179_9981# a_11140_10107# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X360 VSS a_4211_67655# a_3668_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.053e+12p ps=1.104e+07u w=650000u l=150000u M=4
X3600 VDD a_4812_13879# a_5199_11791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3601 a_17803_36649# a_17863_36595# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X3602 a_11067_46823# a_27250_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=0p ps=0u w=1e+06u l=150000u M=8
X3603 a_18829_29423# a_18551_29451# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X3604 VSS a_3162_43023# a_3339_43023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u M=5
X3605 a_4625_50613# a_4407_51017# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X3606 vcm_commonmode a_16362_67214# a_48490_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3607 a_16746_58180# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X3608 VDD a_12877_16911# a_39362_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3609 a_9652_59887# a_6417_62215# a_9431_60214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X361 VSS a_12983_63151# a_43774_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3610 a_19005_47741# a_18626_47375# a_18933_47741# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3611 VSS a_8197_31599# a_15207_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3612 a_21424_49007# a_20161_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3613 a_28699_48169# a_27869_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X3614 VSS a_12877_16911# a_21686_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3615 VSS a_12981_62313# a_33734_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3616 a_10341_10703# a_9642_10357# a_10259_10703# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3617 a_36448_47375# a_22291_29415# a_36357_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X3618 vcm_commonmode a_16362_59182# a_38450_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3619 a_37846_9460# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X362 a_40762_64202# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3620 a_10901_52245# a_4339_64521# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3621 VSS a_12355_15055# a_46786_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3622 a_30991_29397# a_30790_30663# a_31209_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X3623 a_33101_40513# a_12357_37999# a_33015_40513# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3624 VDD a_12680_53511# a_11303_53511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X3625 a_42466_57174# a_16746_57176# a_42374_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3626 a_43774_18894# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3627 VSS VDD a_29718_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3628 a_23467_41237# a_19629_39631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3629 a_25398_67214# a_16746_67216# a_25306_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X363 a_5823_57961# a_4119_70741# a_5905_57711# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X3630 a_14983_51157# a_17475_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3631 a_2787_30503# a_13143_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3632 a_12987_52271# a_12755_53030# a_12818_52521# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3633 a_27245_41829# a_26815_42405# a_27747_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3634 VDD a_12355_65103# a_34342_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3635 VSS a_20957_36604# a_20649_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3636 a_2163_63293# a_1586_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3637 a_26137_29789# a_26063_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X3638 VDD VSS a_47394_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3639 a_17280_48695# a_7050_53333# a_17422_48502# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X364 a_22448_37253# a_21479_36965# a_22411_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X3640 VSS a_35463_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3641 a_18611_52047# a_28963_28853# a_28921_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3642 a_34482_29941# a_37503_31393# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3643 a_20535_51727# a_19877_52245# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X3644 VDD a_38454_34191# a_39331_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3645 a_23694_62194# a_12981_62313# a_23298_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3646 VSS a_12895_13967# a_20682_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3647 a_6457_64489# a_6095_44807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3648 a_11067_13095# a_15103_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3649 VDD a_4803_63669# a_4734_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X365 a_7921_74581# a_7755_74581# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3650 a_7890_54223# a_7519_59575# a_7800_54223# VSS sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X3651 a_35346_72234# VDD a_35838_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3652 VSS a_3339_32463# a_18162_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3653 VDD a_9599_57141# a_9557_57167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3654 VDD a_11521_66567# a_11763_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.646e+11p ps=2.94e+06u w=420000u l=150000u
X3655 a_35838_60508# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3656 a_48398_71230# a_12901_66665# a_48890_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3657 VSS a_1775_60663# a_1775_60439# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3658 a_48890_20504# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3659 a_48490_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X366 a_7387_66781# a_2952_66139# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3660 a_25368_28995# a_9529_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3661 a_12335_50639# a_11711_50645# a_12227_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X3662 a_8635_61751# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X3663 a_19374_58178# a_16746_58180# a_19282_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3664 vcm_commonmode VSS a_16362_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3665 a_2672_26159# a_1757_26159# a_2325_26401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3666 a_4831_58497# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3667 a_22294_70226# a_16362_70226# a_22386_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3668 a_37307_29423# a_30788_28487# a_22843_29415# VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X3669 a_21686_14878# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X367 a_10570_25625# a_9669_26703# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3670 VDD a_1586_69367# a_4719_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3671 a_2040_17289# a_1757_16917# a_1945_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.499e+11p ps=2.35e+06u w=420000u l=150000u
X3672 a_38850_12472# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3673 VDD a_2467_53034# a_1987_52484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3674 VDD a_12546_22351# a_42374_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3675 a_22352_39429# a_21479_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X3676 a_25798_71552# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3677 VDD a_5309_25853# a_5405_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X3678 VDD a_12985_19087# a_22294_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3679 VDD a_11067_67279# a_25306_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X368 a_20754_37455# a_18127_35797# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3680 a_40762_68218# a_12901_66959# a_40366_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3681 a_1881_63151# a_1846_63403# a_1643_63125# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3682 VDD a_2596_16911# a_3166_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3683 a_49402_12870# a_16362_12504# a_49494_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3684 VSS a_38067_47349# a_16955_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3685 a_28410_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3686 a_25306_61190# a_16362_61190# a_25398_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3687 VSS a_12901_66959# a_49798_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3688 a_46786_66210# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3689 a_7457_56053# a_6927_56873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X369 VDD a_9865_14441# a_10589_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X3690 vcm_commonmode a_16362_21540# a_35438_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3691 a_38450_24552# VDD a_38358_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3692 VDD a_7755_26703# a_8123_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3693 a_4427_25071# a_3983_25321# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3694 vcm_commonmode a_16362_66210# a_24394_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3695 a_2672_15113# a_1591_14741# a_2325_14709# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X3696 a_16648_44869# a_15193_44005# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X3697 a_37733_37477# a_38315_38053# a_39247_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3698 a_1925_22583# a_2021_22325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3699 vcm_commonmode a_16362_20536# a_48490_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X37 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u M=1397
X370 a_19282_70226# a_12516_7093# a_19774_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3700 a_18695_47349# a_18500_47491# a_19005_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X3701 a_33830_63520# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3702 a_29814_70548# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3703 VDD a_19780_37253# a_19684_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X3704 a_7650_35951# a_7598_36103# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=0p ps=0u w=650000u l=150000u M=4
X3705 a_43774_59182# a_12727_58255# a_43378_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3706 VSS a_12947_56817# a_40762_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3707 a_37846_18496# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3708 a_26402_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3709 a_24387_47375# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X371 VSS a_12901_58799# a_33734_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3710 a_19877_41972# a_19967_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3711 VDD a_12727_13353# a_41370_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3712 a_8902_36469# a_8017_36495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3713 a_26706_69222# a_12516_7093# a_26310_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3714 a_29322_60186# a_16362_60186# a_29414_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3715 VDD a_23789_39100# a_24201_39126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3716 VDD a_5515_32661# a_5502_33053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3717 vcm_commonmode a_16362_12504# a_38450_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3718 a_2467_53034# a_2559_52789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3719 a_2981_16367# a_2283_15797# a_2899_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X372 a_26706_63198# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3720 a_48398_18894# a_16362_18528# a_48490_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3721 a_42466_10496# a_16746_10494# a_42374_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3722 a_4687_18543# a_4241_18543# a_4591_18543# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X3723 VDD a_11320_16367# a_11495_16341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3724 a_19028_35823# a_18851_35823# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3725 a_25398_20536# a_16746_20534# a_25306_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3726 a_20286_9858# a_16362_9492# a_20378_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3727 a_15285_52245# a_15557_52245# a_15956_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X3728 a_38754_7850# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3729 a_42374_67214# a_16362_67214# a_42466_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X373 VDD a_4685_37583# a_8570_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X3730 a_47790_58178# a_12901_58799# a_47394_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3731 VSS VSS a_44778_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3732 VDD a_8583_33551# a_33479_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3733 VSS a_12355_65103# a_27710_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3734 a_30418_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3735 a_49876_37608# a_49984_39288# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=3.32e+06u as=0p ps=0u w=500000u l=150000u M=4
X3736 a_4951_44330# a_5043_44085# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3737 a_25398_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3738 a_29943_36965# a_27600_36165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3739 a_45878_68540# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X374 vcm_commonmode a_16362_71230# a_36442_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3740 a_11339_24233# a_11480_23957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X3741 a_16080_28111# a_10873_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.2575e+11p pd=3.91e+06u as=0p ps=0u w=650000u l=150000u
X3742 VSS a_12257_56623# a_17670_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3743 VDD a_9955_21807# a_10665_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3744 VDD a_37557_32463# a_39113_32204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3745 a_21686_55166# VSS a_21290_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3746 a_19591_50943# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3747 VDD a_12355_15055# a_27314_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3748 a_32426_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3749 a_19374_11500# a_16746_11498# a_19282_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X375 a_7844_68367# a_6224_73095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3750 a_2012_68565# a_2191_68565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3751 VSS a_2223_28617# a_3983_25321# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3752 a_10754_69501# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X3753 VDD a_12895_13967# a_18278_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3754 a_2672_49929# a_1591_49557# a_2325_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X3755 a_49894_67536# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3756 a_46390_64202# a_11067_13095# a_46882_64524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3757 a_22690_63198# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3758 a_46482_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3759 a_7925_72399# a_7571_72512# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X376 VSS a_29927_29199# a_36487_46859# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3760 VSS a_41351_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3761 a_19282_68218# a_16362_68218# a_19374_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3762 a_41862_7452# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3763 a_49402_57174# a_16362_57174# a_49494_57174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3764 a_17187_31287# a_17459_31145# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X3765 a_23193_52245# a_23487_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3766 a_12073_18543# a_10883_18543# a_11964_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X3767 VSS a_12947_23413# a_36746_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3768 vcm_commonmode a_16362_57174# a_31422_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3769 a_40762_21906# a_12985_7663# a_40366_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X377 a_20682_67214# a_12727_67753# a_20286_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3770 VDD a_18445_46805# a_18475_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3771 a_36350_56170# a_12947_56817# a_36842_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3772 VSS a_40743_31287# a_31659_31751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3773 VDD a_10515_22671# a_43378_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3774 VSS a_10515_23975# a_49798_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3775 a_20286_22910# a_10515_23975# a_20778_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3776 a_7201_56079# a_7169_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3777 VDD a_40383_29575# a_28841_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X3778 a_42283_39095# a_41351_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3779 VDD a_12727_67753# a_26310_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X378 VDD a_2847_71615# a_2834_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3780 a_24849_51183# a_24683_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X3781 VDD VDD a_27314_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3782 VSS VDD a_23694_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3783 a_10216_49929# a_9301_49557# a_9869_49525# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3784 a_26402_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3785 a_31280_40517# a_30311_40229# a_31184_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3786 a_4968_13647# a_3019_13621# a_4866_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X3787 a_20341_30287# a_7862_34025# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X3788 a_43774_12870# a_10055_58791# a_43378_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3789 a_6625_29941# a_5449_25071# a_6782_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X379 a_24961_48783# a_24209_48463# a_24683_48463# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X3790 a_5451_14735# a_4629_13647# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.195e+12p pd=1.039e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X3791 a_1887_34863# a_1915_35015# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3792 a_40981_37253# a_25133_37571# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X3793 a_26706_22910# a_11067_21583# a_26310_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3794 VSS a_12516_7093# a_35742_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3795 a_24302_21906# a_11067_21583# a_24794_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3796 a_24302_17890# a_16362_17524# a_24394_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3797 VDD a_12727_15529# a_30326_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3798 a_26321_50095# a_26155_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3799 vcm_commonmode a_16362_61190# a_39454_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_33830_15484# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X380 a_29322_11866# a_16362_11500# a_29414_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3800 a_43455_31055# a_12907_27023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3801 a_49984_39288# a_49750_39288# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X3802 a_43470_18528# a_16746_18526# a_43378_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3803 a_26505_31599# a_26157_31605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X3804 VDD a_12901_58799# a_47394_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3805 vcm_commonmode a_16362_15516# a_40458_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3806 a_12579_43983# a_12325_44310# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3807 a_47790_11866# a_12985_16367# a_47394_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3808 VSS a_10901_54201# a_10835_54269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3809 a_17766_55488# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X381 a_19780_37253# a_18811_36965# a_19684_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X3810 a_27314_12870# a_12877_16911# a_27806_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3811 VDD a_8201_62839# a_7619_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X3812 a_40458_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3813 a_31822_10464# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3814 a_25306_7850# VSS a_25398_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3815 a_23774_49871# a_6835_46823# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=0p ps=0u w=650000u l=150000u M=4
X3816 a_16362_61190# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X3817 vcm_commonmode a_16362_14512# a_44474_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3818 a_22441_28879# a_13357_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X3819 VSS a_12985_16367# a_17670_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X382 VDD a_12899_10927# a_47394_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3820 a_6825_20969# a_3339_43023# a_6743_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3821 VSS config_1_in[9] a_1591_7119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3822 a_5081_50095# a_2840_66103# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3823 a_40366_19898# a_11067_67279# a_40858_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3824 vcm_commonmode VSS a_27406_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3825 a_7499_74031# a_6098_73095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3826 a_23685_29111# a_23734_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3827 VDD a_1952_60431# a_3123_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3828 a_18307_27791# a_17774_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3829 a_44474_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X383 a_44874_15484# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3830 a_22294_63198# a_12981_62313# a_22786_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3831 VSS a_35217_44509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X3832 a_25077_28129# a_23195_29967# a_24991_28129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3833 VSS a_12901_58799# a_32730_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3834 vcm_commonmode a_16362_16520# a_17366_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3835 VDD VDD a_34342_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3836 a_26310_18894# a_12895_13967# a_26802_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3837 a_21382_14512# a_16746_14510# a_21290_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3838 VSS a_5682_69367# a_10239_57167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3839 a_30818_16488# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X384 a_41370_12870# a_12877_16911# a_41862_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3840 a_34434_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3841 vcm_commonmode a_16362_9492# a_30418_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3842 vcm_commonmode a_16362_10496# a_31422_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3843 a_17366_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3844 a_19678_60186# a_12981_59343# a_19282_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3845 a_7634_61519# a_7580_61751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3846 VSS a_1644_58773# result_out[4] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X3847 a_19678_19898# a_12895_13967# a_19282_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3848 a_33430_67214# a_16746_67216# a_33338_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3849 a_47486_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X385 a_44778_21906# a_12985_7663# a_44382_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3850 VDD config_2_in[5] a_1591_37039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3851 a_11921_59709# a_11710_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X3852 VSS a_9355_32117# a_9318_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3853 a_2107_39049# a_1591_38677# a_2012_39037# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X3854 VSS a_1586_69367# a_5179_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3855 a_46482_66210# a_16746_66212# a_46390_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3856 a_1881_59709# a_1846_59475# a_1643_59317# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3857 a_12800_36189# a_12549_35836# a_12579_35862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X3858 a_45386_21906# a_16362_21540# a_45478_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3859 a_33313_51157# a_33697_50359# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X386 VSS a_29545_28023# a_11619_3303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3860 a_21290_69222# a_12901_66959# a_21782_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3861 VSS a_12907_56399# a_16362_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X3862 a_3143_22364# a_2847_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X3863 a_12687_34191# a_12510_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3864 VSS a_12899_10927# a_41766_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3865 a_5173_69929# a_4985_69725# a_5091_69685# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3866 a_10280_31171# a_4903_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3867 VSS a_6327_72917# a_6271_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3868 a_27710_71230# a_12947_71576# a_27314_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3869 a_10526_22057# a_10073_23439# a_10526_21807# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X387 a_9278_55311# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X3870 a_22386_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3871 a_49402_20902# a_16362_20536# a_49494_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3872 VDD a_37885_42333# a_37491_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3873 a_8531_70543# a_2689_65103# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X3874 a_23727_28335# a_17869_28585# a_23593_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X3875 a_10786_19881# a_5671_21495# a_8933_22583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X3876 a_24042_30083# a_20881_28111# a_23946_30083# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3877 a_49798_65206# a_10975_66407# a_49402_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3878 VDD a_4995_13103# a_4681_13621# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X3879 a_32887_44581# a_32121_44545# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X388 a_18370_23548# a_16746_23546# a_18278_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3880 VSS a_6519_65301# a_1823_76181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3881 a_42770_13874# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3882 a_17613_30287# a_16228_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X3883 VDD a_75162_39738# a_75111_39506# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3884 a_43470_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3885 a_33830_71552# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3886 a_4187_60673# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3887 a_25702_23914# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3888 a_28056_37253# a_27981_37477# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3889 VDD a_1775_60663# a_2141_61635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X389 a_29545_40193# a_28931_39679# a_29804_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X3890 VSS a_2292_17179# a_4025_10749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3891 a_26402_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3892 a_37446_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3893 a_39758_57174# a_10515_22671# a_39362_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3894 a_21663_35327# a_17863_36595# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X3895 a_32826_57496# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3896 vcm_commonmode a_16362_68218# a_46482_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3897 a_9019_30287# a_6649_25615# a_8923_30287# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X3898 a_39305_32463# a_39113_32204# a_39223_32463# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3899 a_19722_49334# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X39 a_33734_21906# a_12985_7663# a_33338_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X390 a_48490_12504# a_16746_12502# a_48398_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3900 VSS a_12895_13967# a_18674_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3901 VDD a_5682_69367# a_6749_66959# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3902 a_29322_9858# a_16362_9492# a_29414_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3903 a_22690_16886# a_12727_13353# a_22294_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3904 a_30485_49257# a_30534_49393# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3905 a_34251_52263# a_35263_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3906 a_2873_13879# a_3023_16341# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3907 VSS a_3280_70501# a_3372_70197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3908 a_25296_40517# a_25221_41281# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X3909 a_18851_51017# a_18335_50645# a_18756_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X391 a_17366_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3910 a_23774_49551# a_6835_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X3911 VSS a_12877_16911# a_32730_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3912 VDD a_31691_32143# a_32371_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3913 VSS a_17039_51157# a_24541_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3914 VSS a_12981_62313# a_44778_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3915 a_41766_60186# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3916 a_40458_58178# a_16746_58180# a_40366_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3917 a_41766_19898# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3918 a_27257_47375# a_22989_48437# a_27175_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3919 a_11709_55777# a_11491_55535# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X392 VSS a_12546_22351# a_46786_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3920 a_23790_59504# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3921 a_5013_20473# a_3247_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X3922 a_19678_14878# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3923 a_38358_24918# VSS a_38850_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3924 VSS a_35196_35425# a_34297_35516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X3925 a_33430_20536# a_16746_20534# a_33338_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3926 vcm_commonmode a_16362_18528# a_32426_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3927 a_42866_22512# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3928 a_3024_67191# a_8675_68047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X3929 a_21686_63198# a_15439_49525# a_21290_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X393 VDD a_10515_23975# a_31330_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3930 a_9041_13763# a_1929_12131# a_8950_13763# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X3931 a_32121_44545# a_32795_44031# a_33727_44265# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3932 VDD a_12899_11471# a_35346_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3933 a_2913_54991# a_2635_55329# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X3934 VDD a_2319_56860# a_2250_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X3935 a_33430_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3936 VSS a_11067_13095# a_48794_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3937 a_46390_72234# VDD a_46882_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3938 a_46882_21508# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3939 a_46482_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X394 VSS a_9314_69367# a_9319_69141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3940 a_26694_29473# a_27234_29789# a_27422_29789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X3941 a_2012_71677# a_1895_71482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3942 a_43378_14878# a_16362_14512# a_43470_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3943 VSS a_12546_22351# a_39758_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3944 a_49402_65206# a_16362_65206# a_49494_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3945 a_43321_29941# a_20267_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X3946 VDD a_36607_34191# a_36713_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3947 a_30577_27497# a_18979_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3948 VSS a_12947_56817# a_38754_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3949 VDD a_18979_30287# a_43530_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X395 a_6782_29967# a_6752_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=9.65e+11p pd=7.93e+06u as=0p ps=0u w=1e+06u l=150000u
X3950 a_28103_38591# a_27337_38565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X3951 VSS a_7210_55081# a_7005_55223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3952 a_49798_9858# a_12985_19087# a_49402_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3953 a_33338_70226# a_16362_70226# a_33430_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3954 a_36842_13476# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3955 a_6608_19319# a_6816_19355# a_6750_19453# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3956 VDD a_12985_16367# a_40366_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3957 a_25702_64202# a_12355_65103# a_25306_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3958 VDD VSS a_39362_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3959 a_2781_15113# a_1591_14741# a_2672_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X396 a_1846_73195# a_2124_73211# a_2080_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3960 a_19774_23516# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3961 a_19374_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3962 VDD a_11067_23759# a_16362_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X3963 VDD a_6559_22671# a_11308_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X3964 a_49894_12472# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3965 a_9417_31849# a_8117_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3966 VDD a_12985_7663# a_23298_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3967 a_20378_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3968 VSS a_36328_49525# a_35403_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X3969 a_47394_13874# a_16362_13508# a_47486_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X397 a_34738_55166# a_8295_47388# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X3970 a_26402_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3971 a_23298_62194# a_16362_62194# a_23390_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3972 a_35438_17524# a_16746_17522# a_35346_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3973 VSS a_19780_37253# a_19743_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X3974 a_39758_10862# a_12546_22351# a_39362_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3975 a_16129_31599# a_16087_31751# a_5595_33205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X3976 vcm_commonmode a_16362_67214# a_22386_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3977 a_7992_17277# a_7649_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X3978 a_26162_49007# a_26662_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X3979 a_6459_30511# a_5915_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X398 VDD a_2099_59861# a_17191_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3980 VDD a_3143_22364# a_4995_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3981 a_49494_24552# VDD a_49402_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3982 vcm_commonmode a_16362_21540# a_46482_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3983 VDD a_12907_27023# a_28902_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X3984 a_19722_49007# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3985 VDD a_10055_58791# a_26310_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3986 VSS a_7862_34025# a_25145_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3987 a_36350_8854# a_12985_19087# a_36842_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3988 a_24394_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3989 VDD a_12983_63151# a_47394_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X399 a_8143_48246# a_6863_42692# a_8071_48246# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3990 a_44874_63520# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3991 a_39454_16520# a_16746_16518# a_39362_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3992 vcm_commonmode a_16362_13508# a_36442_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3993 a_3475_19453# a_3325_18543# a_3112_19319# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X3994 a_11711_24847# a_9955_20969# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3995 a_26319_37429# a_26495_37429# a_26447_37455# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X3996 a_41597_29967# a_41243_30080# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3997 a_10492_60809# a_9577_60437# a_10145_60405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3998 a_11057_25077# a_9669_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3999 a_40458_11500# a_16746_11498# a_40366_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 a_44874_9460# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X40 a_30326_72234# VSS a_30418_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X400 a_31330_64202# a_16362_64202# a_31422_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4000 a_12489_51005# a_12445_50613# a_12323_51017# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X4001 VDD a_17869_28585# a_22762_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.55e+11p ps=5.31e+06u w=1e+06u l=150000u
X4002 a_3981_10357# a_3763_10761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X4003 a_30722_17890# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4004 a_17507_52047# a_16863_29415# a_37277_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X4005 a_38754_58178# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4006 VSS a_11619_3303# a_12171_3311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4007 a_35431_31751# a_35815_31751# a_35581_31599# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X4008 a_18674_8854# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4009 VDD a_39449_39868# a_39055_39913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X401 a_34738_13874# a_12877_16911# a_34342_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4010 a_40366_68218# a_16362_68218# a_40458_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4011 VDD a_15439_49525# a_21290_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4012 a_48890_62516# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4013 a_11667_63303# a_11943_63125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X4014 a_3325_18543# a_2847_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X4015 VDD a_11525_57953# a_11415_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4016 a_22352_38341# a_21479_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4017 VDD a_5877_70197# a_5208_70063# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4018 a_8297_31375# a_2787_32679# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X4019 a_9218_25321# a_5449_25071# a_9135_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X402 a_5962_41391# a_5490_41365# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X4020 a_25263_39913# a_24331_39679# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4021 vcm_commonmode a_16362_57174# a_29414_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4022 VSS a_7155_55509# a_9544_61635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4023 a_9794_51549# a_9668_51451# a_9390_51435# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X4024 a_2199_31599# a_1849_31599# a_2104_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4025 a_12889_39889# a_19703_38695# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4026 VDD a_1591_16367# a_1768_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4027 a_32334_10862# a_16362_10496# a_32426_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4028 a_22294_71230# a_12901_66665# a_22786_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4029 a_43378_59182# a_16362_59182# a_43470_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X403 a_2203_40303# a_1757_40303# a_2107_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X4030 a_5445_63151# a_5595_63125# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4031 a_16640_51183# a_8132_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4032 a_18278_61190# a_12981_59343# a_18770_61512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4033 VSS a_3668_56311# a_6743_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4034 VDD a_22989_48437# a_27425_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X4035 a_26310_69222# a_16362_69222# a_26402_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4036 VDD a_12981_62313# a_25306_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4037 a_3275_73658# a_3978_74183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4038 a_30418_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4039 VDD a_2606_41079# a_8357_48246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X404 a_17670_65206# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4040 a_8332_59049# a_8199_58229# a_7871_59049# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X4041 VSS a_8082_56775# a_7169_56311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4042 a_21782_8456# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4043 a_20378_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4044 VDD a_12895_13967# a_29322_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4045 a_47394_58178# a_16362_58178# a_47486_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4046 a_10680_54171# a_11127_53544# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=0p ps=0u w=650000u l=150000u
X4047 a_15661_29967# a_14926_31849# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4048 a_33734_63198# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4049 a_5274_62313# a_4797_62063# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X405 a_27320_39429# a_26447_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4050 a_34342_18894# a_12895_13967# a_34834_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4051 VSS a_12899_3311# a_34738_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4052 a_15829_28879# a_6459_30511# a_15661_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4053 vcm_commonmode a_16362_71230# a_43470_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4054 VSS a_37699_27221# a_38524_28585# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4055 VSS a_12901_66959# a_23694_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4056 a_23946_30083# a_7939_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4057 a_20682_66210# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4058 VDD a_12947_8725# a_31330_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4059 a_2322_72631# a_2571_72040# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=0p ps=0u w=650000u l=150000u
X406 a_6473_40277# a_6607_42167# a_6909_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4060 a_16746_12502# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4061 a_47394_17890# a_12899_10927# a_47886_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4062 VSS a_12947_23413# a_47790_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4063 VSS a_4191_33449# a_21003_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4064 a_6671_40630# a_5885_39759# a_6671_40303# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4065 VDD a_26495_41781# a_26319_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4066 vcm_commonmode a_16362_20536# a_22386_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4067 a_31330_22910# a_10515_23975# a_31822_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4068 VSS a_1586_51335# a_10975_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4069 VDD a_34923_32375# a_17599_52263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X407 vcm_commonmode VSS a_41462_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4070 a_24394_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4071 a_21290_55166# VSS a_21382_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4072 a_38450_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4073 VSS a_12727_13353# a_37750_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4074 a_35568_49525# a_2959_47113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X4075 a_2834_71311# a_1757_71317# a_2672_71689# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X4076 a_20378_71230# a_16746_71232# a_20286_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4077 vcm_commonmode a_16362_70226# a_47486_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4078 a_41766_13874# a_12877_16911# a_41370_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4079 VSS a_1761_39215# a_31223_36369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X408 a_17766_17492# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4080 a_15871_39913# a_15931_39859# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X4081 a_24698_65206# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4082 a_12901_66415# a_11067_66191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4083 a_24794_17492# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4084 a_24698_23914# a_10515_23975# a_24302_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4085 a_21290_14878# a_12877_14441# a_21782_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4086 VSS a_6243_30662# a_6194_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4087 a_42807_31849# a_41842_27221# a_20267_30503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X4088 a_22294_18894# a_16362_18528# a_22386_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4089 a_10791_27247# a_8935_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=0p ps=0u w=650000u l=150000u M=2
X409 a_20161_48463# a_19991_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4090 a_42374_68218# a_12727_67753# a_42866_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4091 VDD a_41597_29967# a_18703_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X4092 vcm_commonmode a_16362_62194# a_37446_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4093 VDD a_11719_28023# a_12713_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4094 a_38358_58178# a_10515_22671# a_38850_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4095 a_41462_60186# a_16746_60188# a_41370_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4096 VDD a_2111_38279# a_2052_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X4097 a_41462_19532# a_16746_19530# a_41370_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4098 VSS a_17867_32117# a_17798_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X4099 VDD a_12727_58255# a_45386_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X41 VSS a_12727_58255# a_32730_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X410 VDD a_12877_14441# a_21290_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4100 a_1761_25615# a_1591_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4101 a_38754_11866# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4102 a_24394_70226# a_16746_70228# a_24302_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4103 a_9204_15113# a_8289_14741# a_8857_14709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X4104 a_27710_56170# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4105 VDD a_10717_17209# a_10747_16950# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4106 VSS a_10147_71855# a_8575_74853# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X4107 a_29119_34473# a_29513_34428# a_27560_34337# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X4108 a_28810_16488# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4109 VSS a_41351_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X411 vcm_commonmode a_16362_69222# a_30418_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4110 a_25306_13874# a_12727_15529# a_25798_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4111 a_20185_30287# a_14625_30761# a_20103_30287# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4112 a_15193_44005# a_15775_44581# a_16707_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X4113 a_5043_19306# a_5135_19061# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4114 VSS a_16917_31573# a_18063_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X4115 vcm_commonmode a_16362_10496# a_29414_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4116 VDD a_2847_12863# a_1929_12131# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4117 a_1644_53877# a_1823_53885# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4118 VDD a_7571_29199# a_11527_28701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4119 VDD a_7439_64213# a_7387_64239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X412 a_45386_11866# a_10055_58791# a_45878_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4120 a_18674_14878# a_12727_15529# a_18278_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4121 VDD a_11617_72097# a_11507_72221# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4122 a_30035_44581# a_29269_44545# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X4123 VSS a_11495_16341# a_5671_21495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X4124 a_27406_61190# a_16746_61192# a_27314_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4125 a_10103_48682# a_10195_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4126 VDD a_12907_27023# a_28721_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4127 a_19282_69222# a_12901_66959# a_19774_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4128 a_23790_67536# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4129 a_20286_64202# a_11067_13095# a_20778_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X413 VSS a_11455_12157# a_11416_12283# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4130 VSS a_2686_70223# a_5091_69685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4131 a_2295_52271# a_1849_52271# a_2199_52271# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X4132 a_33338_63198# a_12981_62313# a_33830_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4133 a_12877_16911# a_11251_59879# a_12805_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X4134 a_7381_35407# a_3305_38671# a_7381_35727# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4135 vcm_commonmode a_16362_16520# a_28410_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4136 a_76365_39738# a_76461_39480# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4137 VDD a_2840_66103# a_19946_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=2
X4138 a_32426_14512# a_16746_14510# a_32334_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4139 a_29942_30663# a_30052_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X414 a_17092_50959# a_7050_53333# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=0p ps=0u w=650000u l=150000u
X4140 VDD a_2325_14709# a_2215_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4141 VSS a_10515_23975# a_23694_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4142 a_45478_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4143 a_3595_73487# a_2971_73493# a_3487_73865# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4144 a_5611_59887# a_2840_53511# a_5421_60137# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X4145 VDD a_12257_56623# a_30326_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4146 a_24683_48463# a_24743_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4147 VSS VDD a_48794_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4148 a_44474_67214# a_16746_67216# a_44382_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4149 VDD a_22843_29415# a_30991_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X415 a_35346_68218# a_12727_67753# a_35838_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4150 vcm_commonmode a_16362_64202# a_41462_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4151 a_6930_37583# a_3305_38671# a_6816_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=4.2e+11p ps=2.84e+06u w=1e+06u l=150000u
X4152 a_43378_22910# a_16362_22544# a_43470_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4153 a_8539_18231# a_7377_18012# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4154 VSS a_3417_33231# a_3805_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X4155 VDD a_4771_56597# a_1823_66941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4156 VDD a_6607_39991# a_6559_39759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4157 VSS a_2939_33535# a_2873_33609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X4158 a_33819_42359# a_33856_42693# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4159 VSS a_7295_44647# a_38837_46983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X416 VDD a_12516_7093# a_42374_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4160 a_26065_31171# a_25263_29981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4161 VSS a_36107_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4162 a_35742_61190# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4163 a_34434_59182# a_16746_59184# a_34342_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4164 a_6373_15521# a_6155_15279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X4165 a_42770_62194# a_12981_62313# a_42374_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4166 a_18674_71230# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4167 a_17366_69222# a_16746_69224# a_17274_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4168 a_25702_72234# VDD a_25306_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4169 a_2215_22173# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X417 a_28318_21906# a_11067_21583# a_28810_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4170 a_16270_24918# VSS a_16362_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4171 VSS a_3987_19623# a_6743_20969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4172 a_20378_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4173 VDD a_33694_30761# a_36001_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X4174 a_9209_24527# a_5449_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4175 a_9307_30663# a_7461_27247# a_9509_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4176 VSS a_32121_40741# a_33727_39913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X4177 a_36600_49159# a_35568_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4178 VSS a_42188_43677# a_41289_43421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X4179 a_39758_60186# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 VSS a_2847_40277# a_2339_38129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4180 a_38450_58178# a_16746_58180# a_38358_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4181 a_42188_43677# a_41351_42405# a_42224_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4182 vcm_commonmode VSS a_35438_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4183 a_39758_19898# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4184 VSS a_24067_42583# a_23880_42325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4185 a_9751_25071# a_9218_25321# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4186 VDD a_2319_73180# a_2250_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X4187 a_40762_14878# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4188 VDD a_21856_36513# a_20957_36604# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X4189 vcm_commonmode a_16362_65206# a_18370_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X419 a_14258_44527# a_14081_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4190 a_19580_49159# a_14985_51701# a_19722_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X4191 a_35665_31849# a_33694_30761# a_35581_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4192 VSS a_18045_39105# a_18731_38825# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X4193 VSS a_7803_55509# a_8941_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4194 VSS a_7457_56053# a_7072_56053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X4195 a_38288_32143# a_38239_32375# a_38197_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X4196 VDD a_7901_13077# a_7797_13885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4197 a_23694_24918# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4198 a_44874_71552# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4199 a_6722_65579# a_7039_65469# a_6997_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X42 a_5147_43567# a_4701_43567# a_5051_43567# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X420 a_34434_60186# a_16746_60188# a_34342_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4200 a_24632_32259# a_22399_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4201 VDD a_2325_49525# a_2215_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4202 a_44382_61190# a_16362_61190# a_44474_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4203 a_7901_61519# a_2952_66139# a_7467_61751# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X4204 a_14273_27791# a_13919_27904# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4205 a_10603_25731# a_10570_25625# a_10521_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4206 a_27314_71230# a_16362_71230# a_27406_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4207 a_6733_69135# a_6008_69679# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X4208 a_26706_15882# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4209 VSS a_12895_13967# a_29718_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X421 a_28318_17890# a_16362_17524# a_28410_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4210 a_36520_41605# a_35647_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4211 a_35299_32375# a_28446_31375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4212 VSS a_12727_15529# a_30722_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4213 VDD a_1950_59887# a_10147_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X4214 a_19629_39631# a_19203_39958# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4215 a_3751_72373# a_4227_73791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X4216 VDD a_11067_21583# a_17274_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4217 VDD a_13239_29575# a_13173_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4218 VDD a_12947_71576# a_21290_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4219 a_48890_70548# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X422 a_34434_19532# a_16746_19530# a_34342_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4220 a_31741_30485# a_27535_30503# a_31994_30511# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X4221 a_20635_29415# a_35539_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X4222 a_2107_49929# a_1591_49557# a_2012_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X4223 a_21382_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4224 a_45782_69222# a_12516_7093# a_45386_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4225 a_2012_66415# a_1895_66628# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4226 VSS a_10975_66407# a_42770_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4227 a_44382_8854# a_12985_19087# a_44874_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4228 VSS a_4571_26677# a_7841_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X4229 a_28959_49783# a_28855_48801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X423 VDD a_12727_58255# a_38358_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4230 vcm_commonmode a_16362_60186# a_30418_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4231 vcm_commonmode a_16362_19532# a_30418_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4232 a_40858_23516# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4233 a_40458_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4234 VDD a_11902_27497# a_13059_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4235 a_3020_54135# a_3228_54171# a_3162_54269# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4236 VSS a_7479_17607# a_7479_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4237 a_3677_13647# a_1929_10651# a_3523_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4238 VDD a_7580_61751# a_8424_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4239 a_6559_22671# a_6435_47893# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X424 a_32426_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4240 a_38754_8854# a_12947_8725# a_38358_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4241 a_44474_20536# a_16746_20534# a_44382_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4242 VDD a_2099_59861# a_2511_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4243 VDD a_12901_66665# a_25306_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4244 a_18370_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4245 a_7749_55535# a_7213_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4246 VDD a_12899_10927# a_33338_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4247 a_30264_44007# a_29391_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4248 a_2859_41935# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X4249 VSS a_12355_65103# a_46786_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X425 a_10045_30287# a_3339_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X4250 a_7994_45565# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X4251 a_34434_12504# a_16746_12502# a_34342_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4252 VDD a_12899_11471# a_46390_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4253 a_5529_16367# a_5363_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4254 a_44474_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4255 a_6733_53903# a_6646_54135# a_4240_53083# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4256 a_41370_15882# a_16362_15516# a_41462_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4257 a_17366_22544# a_16746_22542# a_17274_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4258 a_2325_23413# a_2107_23817# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X4259 a_2107_51183# a_1757_51183# a_2012_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X426 VDD a_27983_40871# a_12663_39783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X4260 a_11955_69653# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4261 a_34342_69222# a_16362_69222# a_34434_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4262 VSS a_6417_62215# a_7295_60751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4263 VDD a_11763_20407# a_10275_21495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X4264 VSS a_23567_35507# a_23507_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4265 VSS a_12257_56623# a_36746_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4266 VDD a_75199_40594# a_75628_40594# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4267 a_19203_39958# a_19245_39747# a_19203_39631# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4268 a_40762_55166# VSS a_40366_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4269 a_15941_31849# a_15911_31784# a_5595_33205# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X427 a_17366_70226# a_16746_70228# a_17274_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4270 a_16746_20534# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4271 a_23933_50095# a_22989_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X4272 VSS a_12983_63151# a_19678_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4273 VSS a_8675_68047# a_3024_67191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X4274 VSS a_12947_56817# a_49798_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4275 a_23694_65206# a_10975_66407# a_23298_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4276 a_12671_42895# a_12417_43222# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4277 a_7649_17455# a_7479_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4278 a_38450_11500# a_16746_11498# a_38358_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4279 a_47886_13476# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X428 a_47486_18528# a_16746_18526# a_47394_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4280 VDD a_5682_69367# a_9821_55862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X4281 VDD a_12895_13967# a_37354_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4282 VDD a_1929_12131# a_8167_11561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4283 VDD a_12901_66959# a_41370_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4284 a_21290_63198# a_16362_63198# a_21382_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4285 a_35838_7452# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4286 a_4083_22351# a_3325_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4287 a_35061_51727# a_29361_51727# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.297e+11p pd=3.25e+06u as=0p ps=0u w=420000u l=150000u
X4288 VDD a_6978_58487# a_6782_58951# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X4289 VDD a_7467_57863# a_6880_58773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X429 a_22294_66210# a_16362_66210# a_22386_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4290 VDD a_2375_49172# a_1895_49722# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4291 VSS a_9215_58487# a_4674_57685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4292 VSS a_2928_67191# a_2559_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4293 VSS a_27937_27247# a_28589_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4294 a_36350_30761# a_29927_29199# a_35959_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X4295 vcm_commonmode a_16362_68218# a_20378_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4296 a_18045_38017# a_18351_37503# a_19283_37737# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4297 a_26706_56170# a_12257_56623# a_26310_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4298 VDD a_9271_52789# a_7217_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4299 a_4812_13879# a_6435_10901# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X43 VSS a_11067_67279# a_32730_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X430 a_27710_57174# a_10515_22671# a_27314_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4300 VSS a_19217_51701# a_12755_53030# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4301 vcm_commonmode a_16362_67214# a_33430_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4302 VDD a_12877_16911# a_24302_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4303 a_15959_44031# a_15193_44005# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X4304 a_53906_40254# a_52778_39936# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4305 a_38358_66210# a_10975_66407# a_38850_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4306 a_7097_63151# a_6559_63401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4307 VSS VDD a_17670_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4308 VDD a_12727_67753# a_45386_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4309 a_42866_64524# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X431 a_76971_38925# a_75794_40594# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=4.74e+06u as=0p ps=0u w=500000u l=500000u M=2
X4310 a_33338_7850# VDD a_33830_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4311 a_23593_28335# a_22577_29111# a_23303_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8025e+11p ps=3.77e+06u w=650000u l=150000u
X4312 VSS a_18811_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4313 VSS a_32795_44031# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4314 vcm_commonmode a_16362_59182# a_23390_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4315 a_12174_12381# a_11455_12157# a_11611_12252# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X4316 a_32730_23914# a_10515_23975# a_32334_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4317 VSS a_12355_15055# a_31726_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4318 a_28410_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4319 a_5713_31849# a_4495_35925# a_5629_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X432 a_18278_13874# a_12727_15529# a_18770_13476# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4320 VSS a_12815_16519# a_12815_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4321 a_45782_22910# a_11067_21583# a_45386_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4322 a_2325_22049# a_2107_21807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X4323 VDD a_12516_7093# a_18278_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4324 a_43378_60186# a_12727_58255# a_43870_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4325 a_18370_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4326 VSS a_10501_55535# a_10317_55223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4327 a_26662_48981# a_28648_50101# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4328 a_7578_47158# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X4329 a_5694_32687# a_2411_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X433 VDD a_11619_56615# a_12479_9633# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4330 vcm_commonmode a_16362_58178# a_27406_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4331 a_12047_57685# a_11872_57711# a_12226_57711# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4332 a_36842_55488# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4333 a_28931_39679# a_28152_40517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X4334 VSS a_38436_29941# a_37699_27221# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4335 a_20286_72234# VDD a_20778_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4336 VDD VDD a_20286_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4337 a_19774_65528# a_19720_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4338 a_20778_60508# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4339 a_29322_22910# a_10515_23975# a_29814_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X434 VDD a_5039_42167# a_15457_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X4340 a_1761_41935# a_1591_41935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4341 a_33338_71230# a_12901_66665# a_33830_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4342 a_19282_55166# VSS a_19374_55166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4343 a_5449_25071# a_5085_23047# a_6143_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X4344 VDD a_7155_55509# a_9626_61635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4345 a_1761_39215# a_1591_39215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4346 a_22132_44129# a_24331_44581# a_25263_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4347 VSS a_34482_29941# a_34423_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X4348 VDD a_19807_28111# a_35539_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X4349 a_18370_71230# a_16746_71232# a_18278_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X435 a_22786_11468# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4350 VSS a_12985_16367# a_36746_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4351 VSS a_6372_38279# a_6835_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8025e+11p ps=3.77e+06u w=650000u l=150000u
X4352 a_19282_14878# a_12877_14441# a_19774_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4353 VSS a_12985_7663# a_19678_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4354 a_4889_55535# a_4533_55799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4355 a_5087_23145# a_5085_23047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X4356 a_34738_61190# a_12355_15055# a_34342_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4357 a_23790_12472# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4358 VDD a_1586_45431# a_9135_49557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4359 a_5418_20719# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X436 a_5378_56989# a_5252_56891# a_4974_56875# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X4360 a_4461_53113# a_3668_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X4361 vcm_commonmode VSS a_41462_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4362 VSS a_5682_69367# a_9821_55862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4363 a_19374_7484# VDD a_19282_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4364 a_10426_51549# a_9707_51325# a_9863_51420# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X4365 a_45386_18894# a_12895_13967# a_45878_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4366 VSS VSS a_45782_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4367 VDD a_2959_47113# a_35061_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4368 VSS a_19807_28111# a_31440_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4369 a_31726_66210# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X437 a_39362_67214# a_12983_63151# a_39854_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4370 VDD a_32695_43455# a_32555_43777# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4371 vcm_commonmode a_16362_15516# a_49494_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4372 vcm_commonmode a_16362_21540# a_20378_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4373 a_23390_24552# VDD a_23298_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4374 a_5331_71855# a_4885_71855# a_5235_71855# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X4375 a_9011_74879# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4376 a_36442_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4377 a_38754_60186# a_12981_59343# a_38358_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4378 VSS a_12899_11471# a_35742_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4379 a_38754_19898# a_12895_13967# a_38358_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X438 a_43378_8854# a_12985_19087# a_43870_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4380 vcm_commonmode a_16362_20536# a_33430_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4381 a_19621_52271# a_19576_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4382 a_6997_65327# a_6519_65301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4383 VDD a_1923_59583# a_1643_64213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4384 a_39854_9460# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4385 a_9528_25071# a_6162_28487# a_9408_25071# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X4386 a_6180_54447# a_6138_54599# a_5877_54421# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4387 a_25417_51425# a_25199_51183# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4388 a_49494_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4389 a_13107_34789# a_12251_39069# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X439 a_43870_65528# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4390 a_19703_38695# a_19919_38695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4391 a_22786_18496# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4392 VDD a_8999_61493# a_8938_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X4393 VSS a_7159_50260# a_6863_49722# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4394 VDD a_12985_19087# a_49402_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4395 a_40366_69222# a_12901_66959# a_40858_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4396 a_26402_15516# a_16746_15514# a_26310_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4397 vcm_commonmode a_16362_12504# a_23390_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4398 vcm_commonmode a_16362_63198# a_35438_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4399 a_36350_59182# a_12901_58799# a_36842_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X44 a_22690_66210# a_12983_63151# a_22294_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X440 a_40366_62194# a_12355_15055# a_40858_62516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4400 a_33338_18894# a_16362_18528# a_33430_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4401 VSS a_17711_32385# a_17672_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4402 VDD a_41820_41501# a_42316_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4403 VDD a_8263_45908# a_7644_46805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4404 a_9943_62607# a_9319_62613# a_9835_62985# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4405 a_49402_19898# a_11067_67279# a_49894_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4406 a_4417_22671# a_3325_18543# a_4333_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4407 VDD a_33963_35507# a_33989_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4408 a_11215_69679# a_10699_69679# a_11120_69679# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X4409 vcm_commonmode a_16362_62194# a_48490_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X441 VSS a_2419_48783# a_10557_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4410 VDD a_5441_27791# a_7030_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4411 a_28757_27247# a_28589_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=6
X4412 a_30943_38695# a_1761_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4413 a_25702_57174# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4414 VSS a_15775_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4415 a_3479_53942# a_3228_54171# a_3020_54135# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4416 a_33856_50101# a_33826_50075# a_33784_50101# VSS sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X4417 a_41462_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4418 vcm_commonmode a_16362_11500# a_27406_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4419 a_37446_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X442 a_19282_8854# a_12985_19087# a_19774_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4420 VSS a_19410_43439# a_26267_43983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4421 VSS a_37885_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4422 a_12157_52047# a_5190_59575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X4423 a_26802_19500# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4424 VSS a_13528_36055# a_12641_36596# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4425 a_30818_68540# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4426 a_25398_62194# a_16746_62196# a_25306_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4427 a_22411_44535# a_21479_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X4428 VSS a_7815_45503# a_7749_45577# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X4429 a_5909_20175# a_4792_20443# a_5825_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X443 vcm_commonmode a_16362_14512# a_48490_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4430 VDD a_1586_51335# a_10975_60975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4431 a_7731_64015# a_2840_53511# a_7635_64015# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X4432 a_5964_67655# a_6094_67825# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.344e+11p pd=1.48e+06u as=0p ps=0u w=420000u l=150000u
X4433 vcm_commonmode a_16362_64202# a_39454_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4434 a_29643_49667# a_28959_49783# a_29561_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4435 a_29718_14878# a_12727_15529# a_29322_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4436 a_44778_23914# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4437 VDD a_20964_31029# a_20911_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X4438 VSS a_11955_69653# a_11889_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4439 a_4515_50639# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X444 a_33830_57496# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4440 VDD a_26417_40193# a_26860_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4441 a_31330_64202# a_11067_13095# a_31822_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4442 a_10400_62985# a_9319_62613# a_10053_62581# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4443 a_34738_15882# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4444 a_16746_69224# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4445 a_2787_30503# a_13239_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X4446 a_16362_64202# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X4447 VSS a_29915_41959# a_18127_35797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4448 VSS a_12947_23413# a_21686_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4449 a_29055_49525# a_28108_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X445 a_39758_22910# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4450 a_18370_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4451 VSS a_24515_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4452 VSS a_1643_54421# a_1591_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4453 a_9955_21807# a_3987_19623# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X4454 a_21290_56170# a_12947_56817# a_21782_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4455 a_3803_35523# a_3697_35523# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4456 a_43774_70226# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4457 a_42466_68218# a_16746_68220# a_42374_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4458 a_2012_39037# a_1895_38842# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X4459 VDD a_9557_64757# a_8896_65015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X446 a_11389_14191# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4460 VDD a_2143_15271# a_10197_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X4461 a_41370_23914# a_16362_23548# a_41462_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4462 a_23628_35823# a_23451_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4463 a_2672_26159# a_1591_26159# a_2325_26401# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4464 a_27710_17890# a_12899_11471# a_27314_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4465 a_4983_66959# a_4351_67279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X4466 a_40762_63198# a_15439_49525# a_40366_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4467 a_2773_4943# a_2603_4943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4468 a_35196_35425# a_35463_36415# a_36395_36649# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X4469 a_4525_36611# a_4242_35407# a_4443_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X447 VSS a_12985_7663# a_43774_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4470 a_22026_27497# a_19889_27497# a_22026_27247# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X4471 a_25306_55166# VSS a_25798_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4472 a_53410_40254# a_52778_39198# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4473 VSS a_1644_72373# result_out[13] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4474 a_16666_72234# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X4475 VDD a_3019_13621# a_2830_15431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4476 VSS a_12516_7093# a_20682_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4477 a_46786_61190# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4478 a_22294_9858# a_16362_9492# a_22386_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4479 a_45478_59182# a_16746_59184# a_45386_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X448 a_29814_8456# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4480 a_2361_74575# a_2083_74913# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X4481 VDD a_6775_53877# a_7519_59575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4482 a_6607_13879# a_5959_13621# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X4483 vcm_commonmode a_16362_61190# a_24394_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4484 a_34834_24520# a_12899_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4485 a_11141_55535# a_10975_55535# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4486 VDD a_5877_70197# a_10697_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4487 VDD a_28670_30663# a_28680_30057# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4488 a_32426_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4489 a_19596_34215# a_18627_34239# a_19500_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X449 a_25702_8854# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4490 VDD a_4906_67509# a_5254_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4491 a_2107_23817# a_1757_23445# a_2012_23805# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4492 VSS a_5607_44343# a_5043_44085# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4493 VSS a_12727_15529# a_28714_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4494 a_25702_10862# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4495 VDD config_2_in[11] a_1591_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4496 a_2203_71689# a_1757_71317# a_2107_71689# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X4497 a_37446_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4498 VSS a_5515_32661# a_5449_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4499 a_13620_36519# a_13349_37973# a_13762_36367# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X45 VDD a_5504_37815# a_5449_37191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X450 VDD a_20715_41245# a_20741_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4500 VDD a_7071_62581# a_5428_63669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4501 a_49494_58178# a_16746_58180# a_49402_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4502 vcm_commonmode VSS a_46482_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4503 a_28295_31287# a_28618_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4504 a_34145_49007# a_33681_49373# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4505 a_4503_10687# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4506 a_38850_23516# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4507 a_7097_67655# a_6224_73095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4508 a_35346_20902# a_12985_7663# a_35838_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4509 a_42866_72556# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X451 VDD a_10975_66407# a_20286_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4510 a_35346_16886# a_16362_16520# a_35438_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4511 a_38450_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4512 VDD a_17039_51157# a_18840_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4513 VDD a_12985_7663# a_42374_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4514 VDD a_3417_31599# a_3799_31063# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4515 a_77451_38925# a_76346_40594# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=4.74e+06u as=0p ps=0u w=500000u l=500000u M=2
X4516 a_42374_62194# a_16362_62194# a_42466_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4517 VDD a_10649_58947# a_10607_58799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X4518 a_12412_32143# a_11711_32143# a_12244_32463# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X4519 a_1985_53387# a_1823_54973# a_1899_53387# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X452 a_46882_56492# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4520 a_7393_58255# a_7210_55081# a_6978_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X4521 a_25306_72234# VSS a_25398_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4522 a_48490_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4523 VSS a_12727_58255# a_27710_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4524 VSS a_30415_50871# a_28968_50871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4525 VSS a_11067_67279# a_27710_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4526 a_43870_7452# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4527 a_22319_38825# a_20713_39105# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4528 VDD a_12877_16911# a_32334_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4529 a_17670_66210# a_12983_63151# a_17274_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X453 a_13643_29199# a_13239_29575# a_14061_29199# VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=8.71e+11p ps=9.18e+06u w=650000u l=150000u M=4
X4530 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4531 VDD a_8643_48767# a_6835_46823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X4532 a_6885_40630# a_5885_39759# a_6671_40630# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4533 a_36116_44765# a_35463_44031# a_36336_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4534 VSS a_9529_28335# a_15788_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X4535 a_2781_19631# a_1591_19631# a_2672_19631# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X4536 a_39362_15882# a_16362_15516# a_39454_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4537 a_8017_36495# a_7479_36495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4538 VDD a_1761_25071# a_32695_43455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4539 VDD a_10055_58791# a_45386_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X454 VSS a_4482_57863# a_33515_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4540 VSS a_5239_20693# a_5173_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X4541 VDD a_12663_35431# a_12651_35645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4542 a_12869_2741# a_22026_27497# a_22890_27247# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u M=4
X4543 a_43470_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4544 a_36746_69222# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4545 VDD a_11067_21583# a_28318_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4546 VSS a_12983_63151# a_40762_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4547 a_9869_67745# a_9651_67503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X4548 VSS a_2787_32679# a_7725_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.6475e+11p ps=4.03e+06u w=650000u l=150000u
X4549 a_32426_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X455 VSS a_3751_72373# a_6921_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u M=4
X4550 vcm_commonmode a_16362_23548# a_38450_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4551 a_18674_9858# a_12985_19087# a_18278_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4552 VSS a_3799_20407# a_3799_20175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4553 a_42466_21540# a_16746_21538# a_42374_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4554 VDD a_12727_15529# a_18278_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4555 a_30722_9858# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4556 a_16362_15516# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4557 a_38171_43983# a_37994_43983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4558 a_31422_66210# a_16746_66212# a_31330_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4559 a_6089_23145# a_5991_21263# a_6007_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X456 a_41766_71230# a_12947_71576# a_41370_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4560 VSS a_2143_15271# a_10204_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4561 VSS a_2411_19605# a_4761_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4562 a_19282_63198# a_16362_63198# a_19374_63198# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4563 a_2847_9813# a_2672_9839# a_3026_9839# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4564 a_3856_70589# a_3588_70589# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.341e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4565 a_19435_51727# a_4758_45369# a_19217_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4566 VSS a_1923_59583# a_6757_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4567 a_30326_21906# a_16362_21540# a_30418_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4568 a_7737_16917# a_7571_16917# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4569 a_10570_49917# a_2419_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X457 a_29814_66532# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4570 a_15261_51433# a_13925_51727# a_15189_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4571 VDD a_15439_49525# a_40366_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4572 VDD a_4903_23983# a_4571_26677# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X4573 VDD a_14258_34191# a_18851_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4574 a_29414_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4575 a_26310_11866# a_16362_11500# a_26402_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4576 a_7833_66415# a_7567_66781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4577 VDD a_12899_10927# a_44382_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4578 VSS a_2319_56860# a_2250_56989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X4579 a_4595_65327# a_4149_65327# a_4499_65327# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X458 a_48490_9492# a_16746_9490# a_48398_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4580 a_16441_41781# a_15459_41781# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X4581 a_45478_12504# a_16746_12502# a_45386_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4582 a_19774_10464# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4583 a_35910_50959# a_30928_49007# a_35683_50613# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=1.9825e+11p ps=1.91e+06u w=650000u l=150000u
X4584 VSS a_10515_22671# a_34738_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4585 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4586 VDD a_1915_24148# a_1867_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4587 a_3019_13621# a_2847_15039# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4588 VSS a_12727_67753# a_17670_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4589 a_37354_61190# a_12981_59343# a_37846_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X459 a_26310_63198# a_12981_62313# a_26802_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4590 a_2289_35113# a_1887_34863# a_2125_34863# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4591 VSS a_21267_52047# a_21831_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.085e+11p ps=7.38e+06u w=650000u l=150000u M=2
X4592 a_45386_69222# a_16362_69222# a_45478_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4593 VSS a_12257_56623# a_47790_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4594 a_11138_12267# a_11416_12283# a_11372_12381# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4595 a_5271_34435# a_2473_34293# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4596 VDD a_2375_13268# a_1895_12730# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4597 a_27314_7850# VSS a_27406_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4598 a_4065_12879# a_1929_10651# a_3983_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4599 a_3969_20175# a_3799_20175# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X46 a_1761_46287# a_1591_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X460 a_12892_36367# a_12641_36596# a_12671_36694# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X4600 a_49494_11500# a_16746_11498# a_49402_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4601 a_17682_50095# a_17493_50639# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=0p ps=0u w=650000u l=150000u M=4
X4602 a_34434_9492# a_16746_9490# a_34342_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4603 VDD a_12895_13967# a_48398_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4604 a_4073_72943# a_4031_73095# a_3978_74183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X4605 VDD a_1586_51335# a_9411_60437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4606 VDD a_12355_65103# a_17274_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4607 a_22386_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4608 a_24698_57174# a_10515_22671# a_24302_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4609 a_49402_68218# a_16362_68218# a_49494_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X461 VSS a_12473_42869# a_12417_43222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4610 vcm_commonmode a_16362_68218# a_31422_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4611 a_40691_30511# a_12447_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4612 VDD a_4443_46607# a_6619_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4613 a_30845_51727# a_28881_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4614 a_36350_67214# a_12983_63151# a_36842_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4615 a_26319_35253# a_12549_35836# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X4616 a_40858_65528# a_39222_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4617 a_1757_40303# a_1591_40303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4618 a_17171_46859# a_4443_46607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4619 VDD a_2479_50899# a_1923_54591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X462 VSS a_2004_42453# a_1948_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4620 a_43470_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4621 vcm_commonmode a_16362_9492# a_32426_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4622 a_40366_55166# VSS a_40458_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4623 VSS a_1586_36727# a_1591_38677# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4624 a_18770_60508# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4625 a_11921_12015# a_11542_12381# a_11849_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4626 a_26402_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4627 a_36746_22910# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4628 a_8662_28111# a_4495_35925# a_8493_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X4629 VDD a_26319_36341# a_19096_36513# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X463 a_30818_61512# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4630 a_22026_27497# a_17222_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X4631 VSS a_1761_34319# a_33155_35839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4632 a_43870_17492# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4633 a_40366_14878# a_12877_14441# a_40858_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4634 VSS a_12985_7663# a_40762_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4635 a_43774_23914# a_10515_23975# a_43378_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4636 VDD a_25493_29967# a_26867_29739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.8025e+11p ps=1.99e+06u w=420000u l=150000u
X4637 a_23298_24918# VSS a_23790_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4638 a_32135_28335# a_22291_29415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4639 VSS a_1761_32143# a_31959_34751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X464 VSS a_12877_16911# a_33734_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4640 VSS a_32970_31145# a_38378_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4641 VDD a_12516_7093# a_29322_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4642 a_2689_65103# a_1768_13103# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4643 a_40276_28335# a_38210_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=0p ps=0u w=650000u l=150000u
X4644 VSS a_2595_47653# a_2553_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4645 vcm_commonmode VSS a_39454_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4646 a_33734_15882# a_12877_14441# a_33338_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4647 a_5550_52637# a_4792_52539# a_4987_52508# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4648 a_6743_23555# a_4571_26677# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X4649 a_29414_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X465 a_25398_14512# a_16746_14510# a_25306_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4650 a_43470_70226# a_16746_70228# a_43378_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4651 a_26310_56170# a_16362_56170# a_26402_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4652 a_33727_44265# a_32121_44545# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X4653 a_32089_35307# a_30757_37455# a_32003_35307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X4654 a_2847_69439# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4655 VDD a_12725_44527# a_27155_40871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4656 a_39222_48169# a_37557_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X4657 VDD a_12899_11471# a_20286_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4658 a_9186_54223# a_6515_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4659 a_44382_13874# a_12727_15529# a_44874_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X466 a_40981_37253# a_41289_36893# a_25133_37571# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4660 a_2347_29245# a_2093_28918# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4661 a_20946_30669# a_14646_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4662 a_29718_66210# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4663 VDD a_2283_15797# a_4075_14191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X4664 a_47886_55488# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4665 a_27314_23914# a_12947_23413# a_27806_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4666 VSS a_19877_41972# a_13349_37973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4667 VDD a_12447_29199# a_28027_29217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4668 a_31330_72234# VDD a_31822_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4669 a_33430_62194# a_16746_62196# a_33338_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X467 a_5713_74895# a_5599_74549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X4670 a_27314_19898# a_16362_19532# a_27406_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4671 a_34834_58500# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4672 a_31822_21508# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4673 a_4307_67477# a_7755_68591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X4674 a_31422_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4675 a_16362_72234# VDD a_16270_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4676 a_37750_14878# a_12727_15529# a_37354_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4677 VSS a_10055_58791# a_34738_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4678 a_15959_42943# a_15193_42917# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X4679 a_46482_61190# a_16746_61192# a_46390_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X468 a_8638_64783# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X4680 vcm_commonmode a_16362_17524# a_43470_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4681 a_19684_39429# a_18811_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4682 VSS a_12947_56817# a_23694_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4683 a_17274_15882# a_12727_13353# a_17766_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4684 VSS a_11067_21583# a_17670_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4685 a_29414_71230# a_16746_71232# a_29322_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4686 a_21782_13476# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4687 VSS a_12985_16367# a_47790_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4688 VDD VSS a_24302_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4689 a_34759_31029# a_39035_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X469 a_29322_56170# a_16362_56170# a_29414_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4690 a_2360_43389# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4691 a_8011_48463# a_2595_47653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4692 a_32334_13874# a_16362_13508# a_32426_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4693 a_14291_50345# a_9963_50959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4694 a_11145_60431# a_10667_60735# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4695 a_20378_17524# a_16746_17522# a_20286_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4696 vcm_commonmode a_16362_16520# a_47486_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4697 a_9135_27023# a_7461_27247# a_9289_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4698 a_6169_44655# a_6095_44807# a_5823_44905# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X4699 a_24698_10862# a_12546_22351# a_24302_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X47 VDD a_10515_22671# a_36350_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X470 VSS a_17358_31069# a_18285_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4700 VSS a_5671_21495# a_6614_21237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4701 vcm_commonmode a_16362_21540# a_31422_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4702 VDD a_10400_62985# a_10575_62911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4703 a_47486_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4704 a_49798_60186# a_12981_59343# a_49402_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4705 a_5021_55357# a_4642_54991# a_4949_55357# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4706 a_49798_19898# a_12895_13967# a_49402_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4707 a_28810_68540# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4708 a_18430_32143# a_17672_32259# a_17867_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4709 VDD a_16917_31573# a_11719_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X471 a_41842_27221# a_42941_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X4710 a_75475_40594# a_75199_40594# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4711 VSS a_14421_49007# a_12516_7093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X4712 a_24394_16520# a_16746_16518# a_24302_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4713 VDD a_11067_67279# a_34342_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4714 vcm_commonmode a_16362_13508# a_21382_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4715 a_38382_31375# a_28446_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X4716 a_23736_7638# a_20635_29415# a_31022_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X4717 a_37446_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4718 a_8021_39221# a_7187_37583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4719 a_1846_59475# a_2124_59459# a_2080_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X472 a_7939_30503# a_8123_34319# a_8656_34639# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=5.4925e+11p ps=5.59e+06u w=650000u l=150000u M=2
X4720 VDD a_4220_68021# a_3143_66972# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X4721 vcm_commonmode a_16362_63198# a_46482_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4722 a_39188_39429# a_38101_38565# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X4723 a_23694_58178# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4724 a_37750_71230# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4725 a_36442_69222# a_16746_69224# a_36350_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4726 a_2250_64605# a_2124_64507# a_1846_64491# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X4727 a_29322_64202# a_11067_13095# a_29814_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4728 a_35346_24918# VSS a_35438_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4729 a_23736_7638# a_30155_32375# a_30939_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X473 a_3212_14441# a_3019_13621# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4730 a_14361_29967# a_14013_30083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X4731 VDD a_17003_49770# a_16891_49220# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4732 VDD a_32121_42369# a_33668_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4733 a_35438_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4734 VSS a_15683_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4735 a_12599_43222# a_12417_43222# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X4736 a_38358_60186# a_16362_60186# a_38450_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4737 a_6641_63151# a_2927_68565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X4738 a_19282_56170# a_12947_56817# a_19774_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4739 a_22562_28023# a_22441_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X474 a_10953_14191# a_10475_14165# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4740 vcm_commonmode a_16362_65206# a_37446_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4741 a_1757_45205# a_1591_45205# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X4742 a_42770_24918# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4743 a_39362_23914# a_16362_23548# a_39454_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4744 a_36579_35831# a_35647_35877# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4745 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4746 a_7933_51183# a_7073_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4747 a_39758_68218# a_12901_66959# a_39362_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4748 VDD a_34943_51335# a_34411_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.85e+11p ps=2.57e+06u w=1e+06u l=150000u
X4749 VSS a_12516_7093# a_18674_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X475 a_20682_20902# a_11067_67279# a_20286_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4750 a_32334_58178# a_16362_58178# a_32426_58178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4751 VSS a_12895_13967# a_48794_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4752 a_45782_15882# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4753 a_16362_23548# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X4754 a_27406_64202# a_16746_64204# a_27314_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4755 VSS a_10515_22671# a_12546_22351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X4756 a_12584_25935# a_11430_26159# a_12484_25935# VSS sky130_fd_pr__nfet_01v8 ad=4.55e+11p pd=4e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X4757 VDD a_12947_71576# a_40366_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4758 a_32334_17890# a_12899_10927# a_32826_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4759 VSS a_12947_23413# a_32730_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X476 a_5515_32661# a_5340_32687# a_5694_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4760 a_29414_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4761 VDD a_12355_15055# a_36350_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4762 a_5975_71829# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X4763 a_16746_15514# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X4764 a_38358_8854# a_12985_19087# a_38850_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4765 a_2672_19631# a_1591_19631# a_2325_19873# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X4766 a_5253_29673# a_2011_34837# a_5169_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4767 a_17366_56170# a_16746_56172# a_17274_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4768 a_18674_17890# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4769 VDD a_8815_13879# a_8026_13885# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X477 VSS a_7939_30503# a_26065_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4770 a_2107_30345# a_1591_29973# a_2012_30333# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X4771 VSS a_12473_41781# a_26495_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4772 a_23390_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4773 a_1757_23445# a_1591_23445# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4774 a_25702_18894# a_12899_10927# a_25306_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4775 a_5639_37699# a_3949_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4776 VSS a_12727_13353# a_22690_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4777 a_49798_14878# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4778 vcm_commonmode a_16362_70226# a_32426_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4779 a_7295_25321# a_5085_24759# a_6162_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X478 a_9382_61225# a_7580_61751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4780 a_34342_11866# a_16362_11500# a_34434_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4781 VSS a_24800_44129# a_25447_43447# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X4782 a_8569_24527# a_8031_24527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4783 vcm_commonmode a_16362_62194# a_22386_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4784 a_6156_67477# a_6224_73095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=700000u l=150000u
X4785 a_5226_21085# a_4149_20719# a_5064_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X4786 a_23298_58178# a_10515_22671# a_23790_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4787 VDD a_12727_58255# a_30326_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4788 VSS a_12877_14441# a_26706_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4789 a_23694_11866# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X479 VDD a_12257_56623# a_23298_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4790 a_21371_52263# a_31084_30485# a_30665_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X4791 a_36442_22544# a_16746_22542# a_36350_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4792 a_12981_62313# a_12712_62313# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X4793 a_45878_24520# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4794 VDD VDD a_17274_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4795 a_35438_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4796 a_12283_36919# a_12343_36893# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X4797 a_75728_39738# a_75824_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4798 a_24667_31055# a_24223_31171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X4799 a_16707_44535# a_15193_44005# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X48 a_10665_58487# a_6417_62215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X480 a_5616_43567# a_4535_43567# a_5269_43809# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4800 a_25204_34215# a_24331_34239# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X4801 a_18627_34239# a_16928_35303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X4802 a_27417_32509# a_28430_32143# a_28618_32143# VSS sky130_fd_pr__nfet_01v8 ad=2.7965e+11p pd=3.21e+06u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X4803 VSS a_2099_59861# a_17429_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4804 VSS a_12983_63151# a_38754_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4805 VSS a_5682_69367# a_5024_67885# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u M=2
X4806 a_35742_64202# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4807 a_30211_48169# a_6831_63303# a_29956_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X4808 a_42770_65206# a_10975_66407# a_42374_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4809 a_8772_63927# a_3024_67191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X481 a_37446_67214# a_16746_67216# a_37354_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4810 VDD a_6473_40277# a_6885_40630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4811 a_30875_41271# a_29943_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X4812 a_40366_63198# a_16362_63198# a_40458_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4813 a_46390_20902# a_12985_7663# a_46882_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4814 a_49894_23516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4815 a_49494_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4816 a_46390_16886# a_16362_16520# a_46482_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4817 a_32730_57174# a_10515_22671# a_32334_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4818 VSS a_2223_28617# a_3104_25321# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4819 a_13867_39958# a_13909_39747# a_13867_39631# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X482 a_8383_27247# a_7939_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4820 a_23790_8456# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4821 VSS a_5595_12167# a_5399_13255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X4822 a_7295_44647# a_17651_30485# a_17771_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.8e+11p pd=5.16e+06u as=5.5e+11p ps=5.1e+06u w=1e+06u l=150000u M=2
X4823 a_45782_56170# a_12257_56623# a_45386_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4824 a_39854_15484# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4825 a_36350_12870# a_12877_16911# a_36842_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4826 a_39758_21906# a_12985_7663# a_39362_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4827 VDD a_12877_16911# a_43378_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4828 a_40858_10464# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4829 a_4065_24233# a_2315_24540# a_3983_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X483 VDD a_14425_37981# a_14031_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4830 a_28714_66210# a_12983_63151# a_28318_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4831 a_12587_51335# a_12683_51329# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X4832 VSS a_2451_72373# a_8059_74746# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4833 a_2747_72007# a_2686_70223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4834 VDD a_10515_23975# a_26310_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4835 vcm_commonmode a_16362_8488# a_46482_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4836 a_7102_39465# a_6473_40277# a_7010_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X4837 VDD a_34699_42035# a_34725_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4838 a_26310_64202# a_16362_64202# a_26402_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4839 a_30418_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X484 a_45782_70226# a_12901_66665# a_45386_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4840 vcm_commonmode a_16362_59182# a_42466_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4841 a_9953_62313# a_9643_63125# a_9424_60949# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4842 a_11993_59709# a_11521_58951# a_11921_59709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4843 a_2672_15113# a_1757_14741# a_2325_14709# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X4844 vcm_commonmode VSS a_36442_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4845 a_18977_27791# a_13390_29575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X4846 VSS a_3327_9308# a_5595_12167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4847 VDD a_7815_19319# a_7756_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X4848 vcm_commonmode a_16362_69222# a_25398_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4849 VDD a_29175_28335# a_40049_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X485 a_36350_22910# a_16362_22544# a_36442_22544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4850 VDD a_12516_7093# a_37354_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4851 a_13762_40719# a_13067_38517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4852 VSS a_23901_44220# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4853 a_36013_50959# a_8531_70543# a_35910_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4854 a_34834_66532# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4855 a_9031_54135# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4856 VDD a_12727_15529# a_29322_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4857 a_27333_52271# a_27167_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4858 a_27406_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4859 a_27305_44011# a_12357_37999# a_27219_44011# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X486 a_30375_51335# a_30947_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X4860 a_34342_56170# a_16362_56170# a_34434_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4861 a_35676_49525# a_29361_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X4862 a_20682_61190# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4863 a_17274_66210# a_16362_66210# a_17366_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4864 VSS a_1761_43567# a_30115_38695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4865 VSS a_19580_49159# a_19531_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4866 VDD a_2686_70223# a_5087_72512# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4867 a_5245_69929# a_5208_70063# a_5173_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X4868 VDD a_7755_11471# a_7917_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.2e+11p ps=3.04e+06u w=1e+06u l=150000u
X4869 VDD a_22351_47893# a_7571_29199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X487 a_7640_49929# a_6559_49557# a_7293_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X4870 a_9759_49551# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X4871 vcm_commonmode a_16362_68218# a_29414_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4872 a_17766_11468# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4873 a_31330_8854# a_16362_8488# a_31422_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4874 VDD a_16928_42919# a_16832_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X4875 VDD a_4758_45369# a_19502_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X4876 a_38850_65528# a_38557_32143# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4877 a_35346_62194# a_12355_15055# a_35838_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4878 VSS a_10515_22671# a_45782_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4879 VSS config_2_in[4] a_1591_35407# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X488 a_3668_56311# a_4351_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4880 VSS a_38077_29941# a_31084_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4881 a_48398_61190# a_12981_59343# a_48890_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4882 a_24698_60186# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4883 a_23390_58178# a_16746_58180# a_23298_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4884 vcm_commonmode VSS a_20378_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4885 a_24698_19898# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4886 a_22291_29415# a_36401_46859# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X4887 a_9955_20969# a_6816_19355# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.4495e+12p pd=1.486e+07u as=0p ps=0u w=650000u l=150000u M=4
X4888 a_37747_27791# a_30788_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X4889 VDD a_2656_70197# a_2686_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X489 a_40458_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4890 VDD a_11067_47695# a_32334_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4891 a_6607_42167# a_6559_27907# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4892 VSS a_12985_7663# a_38754_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4893 a_1761_49007# a_1591_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4894 a_31422_8488# a_16746_8486# a_31330_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4895 a_36746_71230# a_12947_71576# a_36350_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4896 VSS a_6473_40277# a_6892_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4897 VDD a_1586_36727# a_1683_33237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4898 a_42316_41831# a_41443_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4899 a_3452_70537# a_3280_70501# a_3856_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.89e+11p ps=1.74e+06u w=420000u l=150000u
X49 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u M=394
X490 a_7921_64239# a_7891_64213# a_7825_64239# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X4900 VDD a_12355_65103# a_28318_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4901 a_25798_61512# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4902 a_1642_22583# a_1738_22325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4903 VDD a_22132_40865# a_22352_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X4904 a_11053_69135# a_10575_69439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4905 a_33689_27791# a_28757_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4906 a_35765_30287# a_32970_31145# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.9e+11p pd=3.8e+06u as=0p ps=0u w=650000u l=150000u
X4907 a_24279_47753# a_23929_47381# a_24184_47741# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X4908 a_7561_36495# a_7001_36495# a_7479_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X4909 a_9390_51435# a_9707_51325# a_9665_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X491 VSS a_4555_55233# a_4516_55107# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4910 a_4229_14191# a_3023_16341# a_4157_14191# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4911 a_32730_10862# a_12546_22351# a_32334_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4912 VDD a_10053_62581# a_9943_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4913 VDD a_2375_76372# a_1823_77821# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4914 a_10862_10091# a_11179_9981# a_11137_9839# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X4915 a_5445_63151# a_5274_62313# a_2944_64488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4916 VDD a_12257_56623# a_18278_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4917 VSS a_30599_28023# a_19720_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4918 a_29322_72234# VDD a_29814_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4919 a_43353_27791# a_41597_29967# a_43270_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X492 VSS a_1644_58229# result_out[3] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X4920 a_41862_18496# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4921 a_41766_24918# VSS a_41370_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4922 a_29814_60508# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4923 a_35438_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4924 a_30912_39429# a_29943_39141# a_30875_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X4925 a_5199_11791# a_4429_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4926 a_30722_69222# a_12516_7093# a_30326_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4927 VSS a_6831_63303# a_26162_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4928 VDD a_6066_28309# a_5823_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X4929 VSS a_38784_42589# a_37885_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X493 a_12895_13967# a_10515_63143# a_12806_13967# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X4930 vcm_commonmode a_16362_12504# a_42466_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4931 VSS a_31543_51335# a_30947_51157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4932 a_2847_36799# a_2672_36873# a_3026_36861# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4933 VDD a_13390_29575# a_17869_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4934 a_2375_29588# a_2467_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4935 VDD a_2325_26401# a_2215_26525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X4936 a_43445_28879# a_43495_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4937 VDD a_1586_66567# a_9319_62613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4938 vcm_commonmode a_16362_22544# a_25398_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4939 VSS a_30625_52245# a_30573_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X494 VSS a_6467_55527# a_7363_62063# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X4940 a_35224_49871# a_34145_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4941 VSS a_2295_17429# a_2292_17179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X4942 a_7285_24527# a_7111_22351# a_7203_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4943 a_44778_57174# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4944 a_3387_66998# a_1770_14441# a_2928_67191# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X4945 a_3608_57527# a_3421_57167# a_3521_57283# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X4946 a_44778_15882# a_12877_14441# a_44382_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4947 a_27710_67214# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4948 VDD a_33641_29967# a_34895_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4949 a_18370_17524# a_16746_17522# a_18278_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X495 a_35742_62194# a_12981_62313# a_35346_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4950 VDD a_34763_47349# a_34711_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4951 VSS a_12355_65103# a_31726_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4952 VDD a_12899_11471# a_31330_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4953 a_3707_28995# a_2216_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4954 vcm_commonmode a_16362_21540# a_29414_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4955 a_32057_37479# a_32365_37692# a_32031_37683# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X4956 VSS a_13107_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4957 a_17670_59182# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4958 a_44474_62194# a_16746_62196# a_44382_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4959 vcm_commonmode a_16362_18528# a_41462_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X496 VSS a_28881_52271# a_36600_49159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4960 a_17712_7638# a_30565_30199# a_30577_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4961 VSS a_32795_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X4962 a_45878_58500# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4963 VSS a_12257_56623# a_21686_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4964 VDD a_7637_69679# a_4351_67279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X4965 a_6611_14967# a_5399_13255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X4966 a_27406_72234# VDD a_27314_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4967 a_26137_29789# a_2787_30503# a_26221_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X4968 a_48794_14878# a_12727_15529# a_48398_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4969 VSS a_10055_58791# a_45782_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X497 a_10661_10383# a_9642_10357# a_10589_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4970 vcm_commonmode a_16362_13508# a_19374_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4971 a_22577_29111# a_9529_28335# a_22757_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4972 a_28318_15882# a_12727_13353# a_28810_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4973 a_23390_11500# a_16746_11498# a_23298_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4974 a_4674_40277# a_7756_19087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X4975 a_32826_13476# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4976 a_9405_31599# a_4903_31849# a_9417_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4977 a_14039_41271# a_13107_41317# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4978 a_4699_18909# a_4075_18543# a_4591_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X4979 VDD a_12985_19087# a_18278_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X498 vcm_commonmode a_16362_22544# a_30418_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4980 VDD a_7939_30503# a_22995_30663# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4981 a_49402_69222# a_12901_66959# a_49894_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4982 a_30326_9858# a_12546_22351# a_30818_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4983 VDD a_12895_13967# a_22294_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4984 VDD a_20592_46983# a_20543_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4985 a_21707_47919# a_21261_47919# a_21611_47919# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X4986 a_4242_35407# a_3803_35523# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X4987 VSS a_4831_58497# a_4792_58371# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4988 a_33597_27247# a_19807_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X4989 a_27234_29789# a_5363_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X499 a_27183_40229# a_26417_40193# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X4990 result_out[6] a_1644_62581# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X4991 a_40366_56170# a_12947_56817# a_40858_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4992 a_5993_32687# a_5515_32661# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4993 VSS a_1586_40455# a_1591_49557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4994 a_26802_69544# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4995 a_23298_66210# a_10975_66407# a_23790_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4996 a_34738_64202# a_12355_65103# a_34342_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4997 vcm_commonmode a_16362_60186# a_18370_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4998 vcm_commonmode a_16362_19532# a_18370_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4999 VDD a_12727_67753# a_30326_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5 a_32765_31287# a_32970_31145# a_32928_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X50 a_46882_14480# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X500 a_18674_72234# VDD a_18278_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5000 VDD a_2473_40821# a_1895_40516# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5001 VSS a_35932_37601# a_35033_37692# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X5002 a_35438_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5003 a_5024_67885# a_5682_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X5004 a_20039_49334# a_19788_48981# a_19580_49159# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5005 a_4314_40821# a_4495_35925# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X5006 VSS a_10901_52245# a_10835_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5007 a_44382_55166# VSS a_44874_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5008 VDD a_11067_23759# a_16362_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X5009 a_35742_72234# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X501 a_7449_60431# a_6559_59879# a_7295_60751# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X5010 a_30722_22910# a_11067_21583# a_30326_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5011 a_19684_38341# a_18811_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X5012 VDD a_12412_32143# a_15080_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X5013 a_27314_65206# a_12355_65103# a_27806_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5014 a_2843_71829# a_2847_71615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5015 a_5169_72765# a_2686_70223# a_5087_72512# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5016 a_48794_71230# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5017 a_47486_69222# a_16746_69224# a_47394_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5018 a_12599_36694# a_12417_36694# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5019 VSS a_2327_54135# a_2327_53903# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X502 VDD VSS a_27314_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5020 VSS a_5691_36727# a_6662_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5021 a_46390_24918# VSS a_46482_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5022 a_44778_10862# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5023 VDD a_15253_43421# a_14859_43447# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X5024 a_17274_57174# a_12257_56623# a_17766_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5025 a_1757_38677# a_1591_38677# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5026 a_2107_18543# a_1757_18543# a_2012_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5027 VDD a_10526_22057# a_8295_47388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X5028 a_21782_55488# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5029 VSS a_29545_35841# a_30139_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X503 VDD a_14831_50095# a_29651_48576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X5030 a_27710_20902# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5031 a_21479_39141# a_20713_39105# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5032 VSS a_12981_59343# a_42770_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5033 a_5453_72097# a_5235_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X5034 a_39454_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5035 VSS a_12901_66665# a_25702_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5036 a_5105_47673# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5037 a_15956_52271# a_7050_53333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5038 VDD a_12985_16367# a_39362_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5039 a_27271_37455# a_1761_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X504 VSS a_2451_72373# a_10239_74575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5040 vcm_commonmode a_16362_65206# a_48490_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5041 a_16746_56172# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X5042 a_2283_15797# a_3166_16911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5043 a_42801_27497# a_41334_29575# a_42718_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X5044 a_17670_12870# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5045 VDD a_9187_51157# a_6795_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5046 a_10216_49929# a_9135_49557# a_9869_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X5047 VSS a_12985_16367# a_21686_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5048 a_2960_60975# a_2775_46025# a_2657_60949# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X5049 a_2847_26133# a_2672_26159# a_3026_26159# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X505 VDD a_28589_27247# a_28757_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=6
X5050 a_37846_7452# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5051 a_6737_60431# a_5024_67885# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5052 vcm_commonmode a_16362_57174# a_38450_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5053 a_2788_17277# a_1591_16917# a_2596_16911# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5054 a_44382_72234# VSS a_44474_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5055 VSS a_12727_58255# a_46786_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5056 a_8079_43732# a_8171_43541# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5057 a_42466_55166# VDD a_42374_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5058 VSS a_11067_67279# a_46786_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5059 VSS a_3016_60949# a_5091_60981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 a_48794_61190# a_12355_15055# a_48398_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5060 a_43774_16886# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5061 a_4503_10687# a_4328_10761# a_4682_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5062 a_12340_29967# a_11803_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X5063 VSS a_12516_7093# a_29718_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5064 VDD a_12755_51562# a_13735_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X5065 a_25398_65206# a_16746_65208# a_25306_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5066 a_41370_10862# a_16362_10496# a_41462_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5067 a_39188_38341# a_37733_37477# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X5068 a_30326_18894# a_12895_13967# a_30818_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5069 VSS VSS a_30722_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X507 VSS a_12899_10927# a_45782_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5070 a_3217_34319# a_2289_35113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=0p ps=0u w=1e+06u l=150000u
X5071 a_6008_69679# a_5682_69367# a_5925_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X5072 a_27406_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5073 a_1881_57711# a_1846_57963# a_1643_57685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5074 VDD a_12981_62313# a_34342_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5075 a_34342_64202# a_16362_64202# a_34434_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5076 a_2250_63517# a_2124_63419# a_1846_63403# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5077 VSS a_3449_54201# a_3383_54269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5078 VDD a_11067_21583# a_47394_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5079 VSS a_12355_15055# a_19678_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X508 a_36579_42359# a_36392_43677# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X5080 VSS VDD a_19678_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5081 a_11151_14428# a_10995_14333# a_11296_14557# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X5082 a_21382_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5083 a_23694_60186# a_12981_59343# a_23298_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5084 VDD a_33764_41831# a_33668_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5085 VSS a_12899_11471# a_20682_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5086 a_23694_19898# a_12895_13967# a_23298_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5087 VSS a_34699_37683# a_34639_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X5088 a_4031_56118# a_3780_56347# a_3572_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X5089 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X509 a_10317_55223# a_10501_55535# a_10480_55107# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5090 a_29718_7850# VDD a_29322_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5091 a_35346_70226# a_12516_7093# a_35838_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5092 VDD a_12727_15529# a_37354_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5093 a_18162_31055# a_13353_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X5094 a_5997_30761# a_5547_31599# a_5915_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5095 a_7464_39215# a_6927_39215# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X5096 a_35069_32463# a_34267_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5097 a_9260_25045# a_9167_24011# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X5098 a_41462_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5099 vcm_commonmode a_16362_63198# a_20378_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 a_46786_20902# a_11067_67279# a_46390_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X510 a_2606_41079# a_3983_44655# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X5100 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5101 VDD a_4685_37583# a_5691_36727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X5102 a_48490_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5103 VSS a_15959_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5104 VSS a_20009_48981# a_19943_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5105 a_21290_59182# a_12901_58799# a_21782_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5106 a_45386_11866# a_16362_11500# a_45478_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5107 a_13848_44135# a_13944_43957# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5108 a_27999_41495# a_1761_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X5109 a_8916_65987# a_7803_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X511 a_2764_33609# a_1683_33237# a_2417_33205# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X5110 a_34434_23548# a_16746_23546# a_34342_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5111 vcm_commonmode a_16362_62194# a_33430_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5112 a_7067_30663# a_5441_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X5113 a_38850_10464# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5114 a_12892_42895# a_12641_43124# a_12671_43222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X5115 a_47486_22544# a_16746_22542# a_47394_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5116 a_7808_48829# a_7557_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X5117 VSS a_7862_34025# a_20185_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5118 a_40981_43781# a_41289_43421# a_39244_41953# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5119 VDD VDD a_28318_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X512 a_21479_39141# a_20713_39105# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X5120 VSS a_12727_67753# a_36746_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5121 a_11793_24527# a_9751_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5122 VDD a_5755_14709# a_5451_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5123 VDD VDD a_22294_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5124 a_22386_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5125 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5126 a_27263_40871# a_1761_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5127 a_28410_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5128 VSS a_8263_45908# a_7644_46805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5129 VSS a_1923_54591# a_1881_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X513 a_5239_20693# a_5064_20719# a_5418_20719# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5130 VSS a_12983_63151# a_49798_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5131 a_46786_64202# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5132 vcm_commonmode VSS a_35438_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5133 VSS a_2663_43541# a_2419_48783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X5134 a_8162_53609# a_8132_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5135 VDD a_23192_27791# a_28733_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5136 vcm_commonmode a_16362_64202# a_24394_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5137 a_45478_7484# VDD a_45386_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5138 VDD a_19096_44129# a_19500_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5139 VSS a_12901_58799# a_39758_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 VDD a_29361_51727# a_31669_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X5140 a_36746_56170# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5141 a_33830_61512# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5142 a_41462_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5143 a_43774_57174# a_10515_22671# a_43378_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5144 a_37846_16488# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5145 a_26706_67214# a_12727_67753# a_26310_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5146 a_9370_60975# a_7210_55081# a_9560_60975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5147 vcm_commonmode a_16362_10496# a_38450_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5148 a_20741_35077# a_21049_34717# a_20715_34717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5149 a_6978_58487# a_6467_55527# a_7192_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X515 a_32730_67214# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5150 vcm_commonmode a_16362_9492# a_26402_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5151 a_43439_28111# a_20359_29199# a_43270_27791# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5152 a_10200_47919# a_9392_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X5153 a_20286_7850# VSS a_20378_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5154 a_3123_53047# a_3231_53047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5155 a_31033_28111# a_30975_28023# a_30599_28023# VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X5156 VDD a_2122_20719# a_2228_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5157 a_19224_37479# a_18351_37503# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X5158 a_30418_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5159 VDD a_1586_45431# a_6559_45205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X516 a_23390_17524# a_16746_17522# a_23298_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5160 a_19559_35561# a_18627_35327# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5161 a_42374_24918# VSS a_42866_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5162 a_29072_38567# a_28103_38591# a_29035_38825# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5163 VDD a_12516_7093# a_48398_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5164 a_45878_66532# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5165 VSS a_9735_63669# a_7676_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5166 VSS VSS a_17670_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5167 a_3327_9308# a_4503_10687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5168 a_48490_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5169 a_25269_27791# a_24991_28129# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X517 a_13947_43447# a_13015_43493# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5170 VDD a_11759_59575# a_11019_59575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5171 a_45386_56170# a_16362_56170# a_45478_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5172 a_31726_61190# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5173 VDD a_10351_12879# a_10753_12559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5174 VDD a_2847_21781# a_2317_28892# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5175 a_30418_59182# a_16746_59184# a_30326_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5176 a_21879_30663# a_20881_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5177 a_8206_29199# a_6649_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X5178 a_28318_66210# a_16362_66210# a_28410_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5179 VSS a_1929_12131# a_4211_11989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X518 VSS a_4067_15797# a_3998_15823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X5180 VSS a_2971_48463# a_2595_47653# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u M=2
X5181 a_9318_32509# a_3339_32463# a_9234_32509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5182 a_35196_35425# a_35463_36415# a_36336_36391# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5183 a_12786_30761# a_12340_29967# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=5.72e+06u as=0p ps=0u w=1e+06u l=150000u
X5184 a_41351_38053# a_39468_37479# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5185 VDD a_3987_19623# a_7821_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5186 VSS a_33963_35507# a_33903_35561# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X5187 VSS a_1644_76181# result_out[15] VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5188 a_49894_65528# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5189 a_46390_62194# a_12355_15055# a_46882_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X519 VDD a_7987_40821# a_8017_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X5190 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5191 a_22386_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5192 VSS a_3143_22364# a_3983_25321# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5193 a_49402_55166# VSS a_49494_55166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5194 a_36507_31573# a_32823_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X5195 a_7457_71017# a_7707_70741# a_7651_71017# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5196 VSS a_11067_21583# a_36746_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5197 a_26247_30761# a_7862_34025# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5198 vcm_commonmode VSS a_31422_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5199 a_48490_71230# a_16746_71232# a_48398_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X52 VDD a_10515_23975# a_20286_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X520 a_27710_10862# a_12546_22351# a_27314_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5200 a_1761_9295# a_1591_9295# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5201 a_39854_57496# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5202 a_34738_72234# VDD a_34342_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5203 VDD VSS a_43378_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5204 a_49402_14878# a_12877_14441# a_49894_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5205 VSS a_12985_7663# a_49798_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5206 a_23790_23516# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5207 a_20286_20902# a_12985_7663# a_20778_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5208 a_20286_16886# a_16362_16520# a_20378_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5209 a_23390_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X521 a_34342_70226# a_16362_70226# a_34434_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5210 VDD a_7862_34025# a_20905_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5211 VDD a_10975_66407# a_26310_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5212 a_10433_12879# a_10317_13647# a_10351_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5213 a_29361_38017# a_28747_37503# a_29679_37737# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5214 a_12245_31599# a_12215_31573# a_12161_31599# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5215 VDD a_4052_37961# a_4227_37887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5216 VSS a_13510_44759# a_13515_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5217 a_4181_73193# a_3751_72373# a_3978_74183# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5218 a_26402_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5219 VDD a_7829_60431# a_7901_61519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X522 VSS a_10515_63143# a_14809_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5220 VSS a_12877_16911# a_39758_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5221 a_9183_72007# a_7707_70741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5222 a_43774_10862# a_12546_22351# a_43378_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5223 a_33668_42919# a_32795_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5224 a_5600_74031# a_5483_74244# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5225 a_23747_31055# a_23303_31171# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5226 a_26802_14480# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5227 a_26706_20902# a_11067_67279# a_26310_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5228 a_2875_61225# a_3016_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5229 a_24302_15882# a_16362_15516# a_24394_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X523 VSS a_35568_49525# a_35487_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.355e+11p ps=3.94e+06u w=650000u l=150000u
X5230 VDD a_10055_58791# a_30326_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5231 VDD a_12257_56623# a_29322_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5232 a_35647_42405# a_34699_42035# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5233 VSS a_26465_48463# a_27009_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X5234 a_9253_30511# a_9204_30663# a_9161_30511# VSS sky130_fd_pr__nfet_01v8 ad=3.9e+11p pd=3.8e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X5235 a_21686_69222# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5236 vcm_commonmode a_16362_18528# a_39454_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5237 VDD a_18979_30287# a_30657_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X5238 a_37922_47695# a_18703_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X5239 VDD a_2325_19873# a_2215_19997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X524 a_22690_59182# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5240 a_43470_16520# a_16746_16518# a_43378_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5241 vcm_commonmode a_16362_13508# a_40458_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5242 vcm_commonmode a_16362_23548# a_23390_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5243 a_36350_71230# a_16362_71230# a_36442_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5244 a_27314_10862# a_12985_16367# a_27806_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5245 a_42770_58178# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5246 VDD a_16152_37601# a_15253_37692# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X5247 a_2824_70197# a_3372_70197# a_3330_70223# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.73e+11p pd=2.98e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5248 a_16746_64204# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X5249 a_25702_68218# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X525 a_10405_16367# a_10239_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5250 a_24302_9858# a_16362_9492# a_24394_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5251 a_5074_41935# a_5039_42167# a_4771_42167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5252 a_16362_18528# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X5253 VSS a_13107_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5254 a_29414_17524# a_16746_17522# a_29322_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5255 a_5725_43567# a_4535_43567# a_5616_43567# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5256 a_30418_12504# a_16746_12502# a_30326_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5257 a_42466_63198# a_16746_63200# a_42374_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5258 a_8123_34639# a_6372_38279# a_8123_34319# VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5259 a_20925_44007# a_20899_44211# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X526 vcm_commonmode a_16362_8488# a_27406_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5260 VSS a_12901_66665# a_33734_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5261 a_7299_59663# a_3143_66972# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5262 VDD a_2284_31287# a_2235_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5263 a_28714_59182# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5264 a_1761_30511# a_1591_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5265 a_22294_61190# a_12981_59343# a_22786_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5266 a_30326_69222# a_16362_69222# a_30418_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5267 VSS a_12257_56623# a_32730_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5268 vcm_commonmode a_16362_14512# a_17366_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5269 VDD a_12901_66665# a_34342_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X527 a_16666_24918# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5270 a_26310_16886# a_12899_11471# a_26802_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5271 a_8152_58575# a_7107_58487# a_8061_58575# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X5272 a_35849_29967# a_7295_44647# a_35765_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5273 a_2163_73085# a_1586_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5274 a_34434_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5275 VDD a_6816_19355# a_8338_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5276 a_17409_51183# a_16219_51183# a_17300_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5277 a_3137_27023# a_2223_28617# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X5278 a_17366_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5279 VSS a_1915_24148# a_1867_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X528 a_8945_74953# a_7755_74581# a_8836_74953# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5280 VDD a_3949_41935# a_4259_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.25e+11p ps=7.65e+06u w=1e+06u l=150000u M=2
X5281 a_33430_65206# a_16746_65208# a_33338_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5282 a_7749_22057# a_7187_20719# a_7653_22057# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5283 VSS a_12889_40977# a_12921_40719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X5284 a_4339_64521# a_10239_57167# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X5285 a_9959_20175# a_4792_20443# a_9872_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=8.65e+11p ps=7.73e+06u w=1e+06u l=150000u
X5286 a_3983_16617# a_3301_16617# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5287 a_19517_31751# a_19626_31751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5288 VDD a_10216_49929# a_10391_49855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5289 VDD a_15661_29199# a_5915_35943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.65e+12p ps=1.53e+07u w=1e+06u l=150000u M=4
X529 VSS a_5085_24759# a_6821_26311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5290 VSS a_17003_49770# a_16891_49220# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5291 a_46482_64202# a_16746_64204# a_46390_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5292 a_5147_19605# a_4839_21495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X5293 a_27659_27275# a_23928_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5294 a_7005_55223# a_6467_55527# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5295 a_8781_71677# a_8746_71443# a_8459_71285# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5296 VSS a_12546_22351# a_34738_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5297 a_48490_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5298 a_21290_67214# a_12983_63151# a_21782_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5299 VSS a_10472_26159# a_12584_25935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X53 VDD a_12727_67753# a_19282_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X530 a_18627_44581# a_16928_44007# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5300 a_37287_51433# a_37423_51335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X5301 a_23192_27791# a_22567_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5302 a_7201_56079# a_3295_62083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5303 a_36442_56170# a_16746_56172# a_36350_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5304 a_37750_17890# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5305 a_44778_9858# a_12985_19087# a_44382_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5306 VSS a_12727_13353# a_41766_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5307 a_19374_66210# a_16746_66212# a_19282_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5308 a_34221_47695# a_33802_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5309 a_7311_60975# a_7060_61225# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X531 VSS a_12899_11471# a_49798_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5310 a_4721_45199# a_4458_45565# a_4308_45431# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5311 a_21686_22910# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5312 a_18278_21906# a_16362_21540# a_18370_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5313 a_21675_43447# a_21712_43781# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X5314 VDD a_1950_59887# a_2511_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5315 a_32730_9858# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5316 VSS a_8251_39367# a_8127_39465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X5317 a_9219_71285# a_9024_71427# a_9529_71677# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X5318 a_46786_72234# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5319 a_17670_61190# a_12355_15055# a_17274_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X532 a_20286_16886# a_12899_11471# a_20778_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5320 a_42374_58178# a_10515_22671# a_42866_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5321 vcm_commonmode VSS a_24394_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5322 a_42770_11866# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5323 a_39362_10862# a_16362_10496# a_39454_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5324 a_27652_38237# a_29943_36965# a_30816_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5325 VSS VSS a_28714_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5326 a_25702_21906# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5327 a_33764_38567# a_32795_38591# a_33727_38825# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5328 VSS a_12355_15055# a_40762_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5329 a_28318_57174# a_12257_56623# a_28810_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X533 a_46786_13874# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5330 a_37446_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5331 a_39758_55166# VSS a_39362_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5332 a_32826_55488# a_11067_47695# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5333 VSS a_12899_11471# a_18674_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5334 a_29322_7850# VSS a_29414_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5335 a_12039_69367# a_11803_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5336 a_22690_14878# a_12727_15529# a_22294_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5337 VDD a_12082_25077# a_12349_25847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5338 VSS a_5691_36727# a_7526_33775# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5339 a_16362_10496# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X534 a_32426_72234# VDD a_32334_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5340 a_31422_61190# a_16746_61192# a_31330_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5341 VDD a_11053_62607# a_11667_63303# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5342 VDD VSS a_41370_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5343 VDD a_2100_24759# a_2007_23957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5344 a_28714_12870# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5345 vcm_commonmode a_16362_58178# a_36442_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5346 a_17766_8456# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5347 a_4425_32687# a_4259_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5348 VSS a_12985_16367# a_32730_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5349 VSS a_5915_30287# a_8480_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X535 a_30875_36919# a_27652_38237# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X5350 VDD a_2695_58951# a_2695_58799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5351 a_36442_9492# a_16746_9490# a_36350_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5352 VSS a_6059_14165# a_5943_15492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5353 a_29847_48734# a_27869_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X5354 a_19282_59182# a_12901_58799# a_19774_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5355 a_10299_20969# a_10590_21263# a_10665_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X5356 a_11323_70045# a_10699_69679# a_11215_69679# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5357 a_33760_44869# a_32887_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X5358 a_37478_52047# a_35568_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5359 a_47790_66210# a_12983_63151# a_47394_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X536 a_47486_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5360 a_12821_20175# a_7377_18012# a_12166_21501# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.48e+11p ps=2.78e+06u w=1e+06u l=150000u
X5361 a_38358_22910# a_10515_23975# a_38850_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5362 VSS a_22259_48981# a_4482_57863# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5363 a_42866_20504# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5364 VDD a_10515_23975# a_45386_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5365 vcm_commonmode a_16362_16520# a_32426_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5366 a_42466_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5367 VSS a_12981_62313# a_17670_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5368 VSS a_3143_22364# a_4897_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X5369 a_18627_40767# a_15397_39631# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X537 a_14945_43781# a_15253_43421# a_14919_43421# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5370 a_7799_12265# a_1929_12131# a_7691_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.4e+11p pd=2.88e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X5371 a_45386_64202# a_16362_64202# a_45478_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5372 VDD a_2012_68565# a_1586_69367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5373 a_15095_41781# a_15271_41781# a_15223_41807# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X5374 a_18811_42405# a_16928_42919# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5375 a_11130_22869# a_11574_22869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5376 a_32426_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5377 vcm_commonmode a_16362_69222# a_44474_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5378 VDD a_12877_14441# a_35346_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5379 VDD a_5915_30287# a_22753_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X538 a_37846_71552# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5380 a_8815_13879# a_9179_13737# a_9114_13763# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X5381 a_30745_27791# a_30975_28023# a_30599_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X5382 VDD a_12727_15529# a_48398_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5383 VDD a_28423_52245# a_28410_52637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5384 a_46390_70226# a_12516_7093# a_46882_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5385 a_46482_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5386 a_43378_12870# a_16362_12504# a_43470_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5387 a_22386_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5388 a_11141_55535# a_10975_55535# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5389 a_49402_63198# a_16362_63198# a_49494_63198# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X539 a_33360_51701# a_34579_50613# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X5390 vcm_commonmode a_16362_63198# a_31422_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5391 a_27009_47919# a_26514_47375# a_26917_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X5392 a_2672_19631# a_1757_19631# a_2325_19873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5393 a_22690_71230# a_17599_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5394 a_21382_69222# a_16746_69224# a_21290_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5395 a_2143_15271# a_5147_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5396 a_36842_11468# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5397 VDD a_14289_29687# a_14646_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5398 a_45478_23548# a_16746_23546# a_45386_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5399 a_13357_32143# a_7695_31573# a_13275_32463# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X54 a_1644_65845# a_1823_65853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X540 vcm_commonmode a_16362_13508# a_24394_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5400 a_2307_52637# a_1683_52271# a_2199_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5401 a_20286_24918# VSS a_20378_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5402 a_19774_21508# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5403 a_19374_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5404 VDD a_11067_23759# a_16362_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X5405 a_49894_10464# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5406 a_12269_56873# a_11619_56615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5407 a_20378_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5408 a_26402_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5409 a_23298_60186# a_16362_60186# a_23390_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X541 VDD a_11067_67279# a_37354_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5410 a_27890_32459# a_28430_32143# a_28618_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X5411 VSS a_26753_37981# a_26445_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X5412 VSS a_12727_67753# a_47790_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5413 VSS a_2787_30503# a_12631_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.6875e+11p ps=4.35e+06u w=650000u l=150000u
X5414 a_35438_15516# a_16746_15514# a_35346_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5415 VSS a_39836_38567# a_39799_38825# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X5416 a_40585_42369# a_41167_42943# a_42040_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5417 VDD a_8509_47673# a_8539_47414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5418 vcm_commonmode a_16362_65206# a_22386_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5419 a_31953_51183# a_28881_52271# a_31543_51335# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=5.07e+11p ps=5.46e+06u w=650000u l=150000u
X542 a_7407_46529# a_1586_45431# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5420 a_36425_28879# a_28305_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5421 a_25398_8488# a_16746_8486# a_25306_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5422 a_24302_23914# a_16362_23548# a_24394_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5423 VDD a_4211_11989# a_4035_11989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5424 VDD a_12546_22351# a_26310_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5425 a_41766_58178# a_12901_58799# a_41370_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5426 a_3026_51183# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X5427 VSS a_2843_71829# a_2789_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5428 a_24698_68218# a_12901_66959# a_24302_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5429 VDD a_12355_65103# a_47394_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X543 a_33338_15882# a_12727_13353# a_33830_15484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5430 a_10501_55535# a_10075_55862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5431 a_21424_49007# a_20161_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5432 a_44874_61512# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5433 VSS a_26523_29199# a_33449_30305# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5434 a_39454_14512# a_16746_14510# a_39362_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5435 vcm_commonmode a_16362_11500# a_36442_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5436 VSS a_23271_50943# a_22989_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5437 VDD a_2865_58799# a_2882_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5438 a_1644_62581# a_1823_62589# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5439 a_11396_60975# a_7773_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X544 a_9653_69831# a_9314_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5440 a_12710_63151# a_11067_13095# a_12541_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5441 a_29718_61190# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5442 a_28410_59182# a_16746_59184# a_28318_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5443 vcm_commonmode a_16362_56170# a_25398_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5444 a_25419_50959# a_28671_30539# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5445 a_35838_19500# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5446 a_30722_15882# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5447 a_3572_56311# a_3780_56347# a_3714_56445# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X5448 a_10257_56377# a_5682_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5449 a_5803_11293# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X545 VSS a_2021_22325# a_37939_43455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5450 VDD a_12257_56623# a_37354_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5451 a_11049_20719# a_9955_21807# a_9955_20969# VSS sky130_fd_pr__nfet_01v8 ad=9.62e+11p pd=9.46e+06u as=0p ps=0u w=650000u l=150000u M=4
X5452 a_40086_28335# a_38436_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=0p ps=0u w=1e+06u l=150000u
X5453 a_17766_63520# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5454 VDD a_32031_37683# a_32057_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X5455 a_18061_29967# a_17358_31069# a_17696_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u M=2
X5456 VDD a_12355_15055# a_21290_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5457 a_6559_50959# a_3325_49551# a_6646_50639# VSS sky130_fd_pr__nfet_01v8 ad=5.525e+11p pd=5.6e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X5458 a_48890_60508# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5459 a_3487_37961# a_2971_37589# a_3392_37949# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X546 a_37354_61190# a_16362_61190# a_37446_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5460 VDD a_26495_36341# a_26319_36341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5461 a_22319_39913# a_21387_39679# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5462 a_38037_41831# a_38345_42044# a_38011_42035# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5463 a_5091_69685# a_5208_70063# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5464 vcm_commonmode VSS a_29414_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5465 VSS a_6978_58487# a_6782_58951# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5466 a_29205_42693# a_29513_42333# a_28717_42917# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5467 vcm_commonmode a_16362_22544# a_44474_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5468 a_2568_29245# a_2317_28892# a_2347_28918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X5469 a_4333_29423# a_1915_35015# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X547 VSS a_23847_47919# a_23540_48981# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X5470 a_43378_57174# a_16362_57174# a_43470_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5471 VDD a_21021_46805# a_21051_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5472 a_26310_67214# a_16362_67214# a_26402_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5473 a_5604_39215# a_4941_35727# a_5414_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X5474 VDD a_12981_59343# a_25306_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5475 a_4792_41167# a_4314_40821# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X5476 VSS a_22521_37692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5477 a_9583_10703# a_9484_11989# a_9414_10383# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5478 VDD config_2_in[12] a_1591_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5479 VDD a_7436_46983# a_7387_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X548 a_19596_34215# a_18627_34239# a_19559_34473# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X5480 VDD a_3049_14343# a_2926_15253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X5481 a_25953_32143# a_25605_32259# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5482 a_6671_51183# a_5909_51433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5483 a_21382_22544# a_16746_22542# a_21290_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5484 a_3394_68413# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5485 VDD a_12907_56399# a_16362_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X5486 a_30818_24520# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5487 a_3805_30083# a_3854_29977# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5488 a_28708_52105# a_27627_51733# a_28361_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5489 a_12970_34191# a_12793_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X549 a_5785_25321# a_5085_24759# a_6143_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X5490 a_20378_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5491 a_2882_54813# a_2124_54715# a_2319_54684# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X5492 a_36746_17890# a_12899_11471# a_36350_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5493 VDD a_3987_19623# a_9955_21807# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5494 a_34342_16886# a_12899_11471# a_34834_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5495 VSS a_13357_32143# a_26065_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5496 a_46482_72234# VDD a_46390_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5497 a_19678_69222# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5498 VSS a_12983_63151# a_23694_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5499 a_20682_64202# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X55 VDD a_20359_29199# a_30104_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3e+11p ps=5.26e+06u w=1e+06u l=150000u M=2
X550 VSS a_39503_43957# a_12907_56399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5500 a_47394_15882# a_12727_13353# a_47886_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5501 VSS a_11067_21583# a_47790_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5502 a_2007_65002# a_2099_64757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5503 VDD a_34759_31029# a_34698_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X5504 a_31330_20902# a_12985_7663# a_31822_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5505 a_4960_40847# a_4259_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5506 a_10109_73487# a_9353_72399# a_10037_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5507 a_31330_16886# a_16362_16520# a_31422_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5508 a_36548_49871# a_36464_49783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5509 VDD a_12901_58799# a_41370_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X551 vcm_commonmode a_16362_63198# a_49494_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5510 VDD a_8531_70543# a_34895_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5511 VSS a_12907_56399# a_16362_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X5512 VDD a_6417_62215# a_7393_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5513 VSS a_12727_15529# a_37750_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5514 a_6825_66665# a_2952_66139# a_6515_67477# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5515 a_7931_10357# a_7736_10499# a_8241_10749# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X5516 VSS a_10239_16911# a_10423_17455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X5517 a_41766_11866# a_12985_16367# a_41370_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5518 VDD a_2840_53511# a_5515_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5519 VSS a_4351_26159# a_4528_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X552 VDD a_8933_22583# a_10665_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.145e+12p ps=1.829e+07u w=1e+06u l=150000u M=4
X5520 VSS a_2656_45895# a_3983_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X5521 a_35647_35877# a_33963_35507# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5522 a_10562_69135# a_9485_69141# a_10400_69513# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5523 VDD a_10492_60809# a_10667_60735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5524 a_30722_56170# a_12257_56623# a_30326_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5525 VDD a_12899_10927# a_27314_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5526 a_24794_15484# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5527 a_21290_12870# a_12877_16911# a_21782_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5528 a_24698_21906# a_12985_7663# a_24302_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5529 a_32928_31171# a_4811_34855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X553 a_6457_64489# a_1823_76181# a_6375_64489# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X5530 a_24515_43493# a_20899_44211# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5531 a_42374_66210# a_10975_66407# a_42866_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5532 a_28410_12504# a_16746_12502# a_28318_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5533 VSS a_1586_21959# a_1591_29973# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5534 vcm_commonmode a_16362_60186# a_37446_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5535 vcm_commonmode a_16362_19532# a_37446_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5536 a_4809_18785# a_4591_18543# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5537 a_17927_31573# a_4443_46607# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5538 a_11525_57953# a_11307_57711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5539 a_9963_50959# a_4298_58951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X554 a_26706_16886# a_12727_13353# a_26310_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5540 a_9485_69141# a_9319_69141# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5541 VDD a_17682_50095# a_23631_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5542 a_4897_27247# a_4627_27613# a_4807_27613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5543 vcm_commonmode VSS a_21382_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5544 VSS a_15775_40229# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5545 a_39758_63198# a_15439_49525# a_39362_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5546 a_15223_41807# a_15193_41781# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5547 VSS a_7841_12167# a_8041_15279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X5548 a_25306_11866# a_10055_58791# a_25798_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5549 VSS a_38628_47349# a_29927_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X555 a_5065_66959# a_4307_67477# a_3668_56311# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X5550 a_46786_8854# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5551 VDD a_12516_7093# a_22294_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5552 VSS a_8167_11561# a_7803_11703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X5553 VDD a_21712_43781# a_21616_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5554 VDD a_12727_58255# a_18278_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5555 a_13975_44527# a_13798_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5556 a_16707_40183# a_15775_40229# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X5557 a_32795_39679# a_31280_40517# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5558 VDD a_11400_26133# a_11430_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5559 a_20505_29967# a_14625_30761# a_20433_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X556 a_12883_31421# a_3339_30503# a_12787_31421# VSS sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5560 a_12371_53903# a_12120_54019# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X5561 a_27406_18528# a_16746_18526# a_27314_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5562 a_26447_36367# a_12641_36596# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=0p ps=0u w=420000u l=150000u
X5563 VDD a_6559_22671# a_9135_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5564 a_19282_67214# a_12983_63151# a_19774_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5565 a_49402_56170# a_12947_56817# a_49894_56492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5566 a_23790_65528# a_18611_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5567 a_20286_62194# a_12355_15055# a_20778_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5568 VSS a_10515_22671# a_30722_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5569 a_2107_51183# a_1591_51183# a_2012_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X557 a_39127_48463# a_20635_29415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X5570 VSS a_12901_66665# a_44778_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5571 a_24556_49551# a_6835_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X5572 a_2764_52271# a_1683_52271# a_2417_52513# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X5573 a_40458_66210# a_16746_66212# a_40366_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5574 a_33668_41831# a_32795_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5575 a_5913_74273# a_5695_74031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X5576 a_33338_61190# a_12981_59343# a_33830_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5577 a_42466_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5578 a_7931_10357# a_7775_10625# a_8076_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X5579 vcm_commonmode a_16362_14512# a_28410_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X558 a_15775_34239# a_14076_35077# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X5580 a_10660_16367# a_10543_16580# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5581 a_33734_8854# a_12947_8725# a_33338_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5582 a_19678_22910# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5583 a_11999_67477# a_11711_67325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5584 a_14655_47919# a_5039_42167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X5585 a_11794_58575# a_11710_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X5586 VSS a_12985_7663# a_23694_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5587 a_1846_64491# a_2163_64381# a_2121_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X5588 a_5541_53359# a_1952_60431# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5589 a_45478_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X559 VSS a_1643_57685# a_1591_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5590 a_26802_56492# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5591 a_11902_27497# a_8935_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5592 a_24331_44581# a_22632_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X5593 a_10295_47919# a_9779_47919# a_10200_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X5594 a_18158_46831# a_5831_39189# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5595 a_21686_71230# a_12947_71576# a_21290_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5596 VSS a_12516_7093# a_48794_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5597 a_44474_65206# a_16746_65208# a_44382_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5598 VSS a_28959_49783# a_28789_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.72e+11p ps=4.36e+06u w=650000u l=150000u
X5599 VSS a_4043_44343# a_2656_45895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X56 a_44382_15882# a_16362_15516# a_44474_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X560 VDD a_14747_31599# a_14926_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X5600 VSS a_22989_48437# a_23577_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X5601 a_43378_20902# a_16362_20536# a_43470_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5602 a_46482_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5603 a_27016_29587# a_27169_30083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X5604 VDD a_2847_45503# a_2834_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5605 VSS a_12985_19087# a_31726_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5606 VSS a_26815_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5607 VSS a_2847_51157# a_2781_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X5608 VSS a_12355_15055# a_38754_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5609 a_34434_57174# a_16746_57176# a_34342_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X561 a_12663_40871# a_32555_43777# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X5610 a_35742_18894# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5611 a_42770_60186# a_12981_59343# a_42374_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5612 vcm_commonmode a_16362_8488# a_48490_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5613 a_42770_19898# a_12895_13967# a_42374_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5614 a_13353_30511# a_12786_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5615 a_17366_67214# a_16746_67216# a_17274_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5616 a_7168_55107# a_6467_55527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5617 a_25702_70226# a_12901_66665# a_25306_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5618 a_47486_56170# a_16746_56172# a_47394_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5619 a_48794_17890# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X562 VSS a_12404_34191# a_12510_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5620 a_41261_28335# a_28817_29111# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=0p ps=0u w=650000u l=150000u M=2
X5621 VDD a_11067_23759# a_16362_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X5622 a_28152_44869# a_27183_44581# a_28115_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5623 VSS a_4674_40277# a_4615_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X5624 a_12672_18115# a_10055_58791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5625 a_7037_19385# a_3247_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5626 a_20378_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5627 a_35438_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5628 a_7217_53047# a_7803_55509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5629 VDD a_15439_49525# a_39362_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X563 a_38450_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5630 VDD a_1761_4399# a_1933_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5631 a_40366_59182# a_12901_58799# a_40858_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5632 a_7142_61225# a_5024_67885# a_7060_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5633 a_11340_25321# a_11069_23983# a_11245_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X5634 VDD a_8453_51727# a_10426_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X5635 a_12662_15939# a_10055_58791# a_12580_15939# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5636 a_22753_29967# a_5915_35943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5637 a_10860_47919# a_9779_47919# a_10513_48161# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5638 a_2369_66415# a_2325_66657# a_2203_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5639 a_28714_61190# a_12355_15055# a_28318_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X564 a_6835_23983# a_6451_22895# a_6989_24233# VSS sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5640 VSS a_12899_10927# a_25702_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5641 VDD a_5024_67885# a_9654_65577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X5642 a_7295_60751# a_7311_60975# a_7449_60431# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5643 a_35438_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5644 VDD config_1_in[7] a_1591_4399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5645 VDD VDD a_16270_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5646 a_33338_8854# a_16362_8488# a_33430_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5647 a_1761_11471# a_1591_11471# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5648 VDD VDD a_47394_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5649 a_5629_31849# a_3607_34639# a_5547_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X565 a_5594_36727# a_5963_36585# a_5897_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5650 VSS a_25939_51157# a_26397_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X5651 a_41462_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5652 a_2847_9813# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5653 a_7460_31055# a_6835_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=150000u
X5654 a_36392_43677# a_35647_42405# a_36579_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X5655 a_30818_58500# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5656 VSS a_12899_11471# a_29718_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5657 a_26706_13874# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5658 VSS a_10055_58791# a_30722_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5659 VSS a_3215_68351# a_3149_68425# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X566 a_25263_41001# a_24331_40767# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X5660 a_11759_63927# a_11803_64239# a_12157_64015# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X5661 a_27406_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5662 a_17766_71552# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5663 VDD a_11067_67279# a_17274_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5664 VDD a_5963_36585# a_7215_36201# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5665 a_32730_68218# a_12901_66959# a_32334_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5666 a_2787_32679# a_6655_46261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5667 VDD a_6515_67477# a_7107_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5668 a_8113_24527# a_6162_28487# a_8031_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X5669 a_37699_27221# a_38210_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X567 a_38754_69222# a_12516_7093# a_38358_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5670 a_2216_42997# a_2040_43401# a_2360_43389# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5671 a_17274_61190# a_16362_61190# a_17366_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5672 a_38754_66210# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5673 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5674 a_22015_28111# a_35959_30485# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5675 VSS a_33591_32375# a_28547_51175# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X5676 a_45782_67214# a_12727_67753# a_45386_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5677 VSS a_11067_13095# a_42770_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5678 vcm_commonmode a_16362_63198# a_29414_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5679 a_36350_23914# a_12947_23413# a_36842_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X568 VSS a_10975_66407# a_35742_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5680 a_50198_39208# ctopn a_49876_41198# VSS sky130_fd_pr__nfet_01v8_lvt ad=4.025e+12p pd=3.144e+07u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u M=4
X5681 VSS a_37885_42333# a_37577_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X5682 a_36350_19898# a_16362_19532# a_36442_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5683 a_7553_48469# a_7387_48469# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X5684 a_40858_21508# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5685 a_40458_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5686 a_22749_50613# a_22531_51017# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X5687 a_43378_65206# a_16362_65206# a_43470_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5688 a_3911_16065# a_1586_9991# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5689 a_35742_59182# a_12727_58255# a_35346_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X569 a_31822_69544# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5690 a_32121_40741# a_32795_39679# a_33668_39655# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5691 a_13983_40719# a_13835_41001# a_13620_40871# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X5692 a_18370_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5693 VDD a_12727_13353# a_33338_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5694 a_7640_45577# a_6725_45205# a_7293_45173# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5695 a_32823_29397# a_40323_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X5696 a_20964_31029# a_20905_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5697 a_17939_36129# a_18127_35797# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5698 a_18674_69222# a_12516_7093# a_18278_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5699 VSS a_2216_16885# a_2150_17289# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X57 a_10897_9839# a_10862_10091# a_10659_9813# VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X570 a_15193_44005# a_15775_44581# a_16648_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X5700 VDD a_10472_52423# a_9271_52789# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5701 VSS a_5749_60039# a_5707_59887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X5702 a_8117_12559# a_3327_9308# a_8117_12879# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5703 a_34434_10496# a_16746_10494# a_34342_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5704 VDD a_12877_14441# a_46390_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5705 a_18045_39105# a_17799_38591# a_18672_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5706 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5707 a_41370_13874# a_16362_13508# a_41462_13508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5708 VDD a_19946_51157# a_19502_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X5709 a_17366_20536# a_16746_20534# a_17274_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X571 a_26402_63198# a_16746_63200# a_26310_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5710 a_20378_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5711 a_15261_51433# a_14859_51183# a_15097_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X5712 a_34342_67214# a_16362_67214# a_34434_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5713 VSS VSS a_36746_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5714 a_20682_72234# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5715 VSS a_12355_65103# a_19678_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5716 VSS a_28305_28879# a_35263_28879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8025e+11p ps=3.77e+06u w=650000u l=150000u
X5717 a_47394_66210# a_16362_66210# a_47486_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5718 VDD a_12899_11471# a_19282_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5719 a_2702_45743# a_2656_45895# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X572 vcm_commonmode a_16362_60186# a_23390_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5720 a_1643_64213# a_1846_64491# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5721 a_25104_51183# a_8123_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X5722 VSS a_8459_71285# a_7707_70741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5723 a_17366_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5724 a_33734_71230# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5725 a_32426_69222# a_16746_69224# a_32334_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5726 VDD a_11619_63151# a_11711_67325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.646e+11p ps=2.94e+06u w=420000u l=150000u
X5727 a_47886_11468# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5728 a_7939_30503# a_8123_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5729 a_2847_44629# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X573 vcm_commonmode a_16362_19532# a_23390_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5730 a_37846_68540# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5731 VDD a_1952_60431# a_4533_55799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X5732 a_31330_24918# VSS a_31422_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5733 VDD a_12983_63151# a_41370_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5734 VDD a_5135_50069# a_6646_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5735 a_20635_29415# a_35539_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5736 VSS a_41427_52263# a_41967_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5737 a_2520_43023# a_2040_43401# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X5738 a_34834_9460# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5739 a_6521_58773# a_6361_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X574 VSS a_24800_44129# a_23901_44220# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X5740 a_41462_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5741 VDD a_4571_26677# a_8189_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5742 VSS a_13620_40871# a_12641_42036# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5743 a_24394_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5744 VDD a_12985_19087# a_44382_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5745 a_15775_36965# a_13557_37999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X5746 a_6825_23555# a_4427_30511# a_6743_23555# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5747 a_41261_28335# a_20635_29415# a_41441_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X5748 VSS a_13005_35823# a_12641_37684# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5749 a_5326_51005# a_2595_47653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X575 a_27806_59504# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5750 VDD a_12985_16367# a_24302_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5751 vcm_commonmode a_16362_65206# a_33430_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5752 a_7195_65564# a_7039_65469# a_7340_65693# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X5753 VSS a_2411_26133# a_3013_42301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5754 result_out[3] a_1644_58229# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X5755 a_38358_64202# a_11067_13095# a_38850_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5756 a_4025_10749# a_3981_10357# a_3859_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5757 VDD a_10975_66407# a_45386_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5758 a_42866_62516# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5759 a_11281_30511# a_11155_30663# a_11183_30761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X576 a_26433_39631# a_26267_39631# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X5760 a_32334_9858# a_12546_22351# a_32826_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5761 a_22063_47594# a_20853_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X5762 a_27710_62194# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5763 a_20927_35877# a_19780_37253# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X5764 a_10321_74575# a_10109_73487# a_10239_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5765 vcm_commonmode a_16362_57174# a_23390_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5766 VSS a_12727_58255# a_31726_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5767 a_32730_21906# a_12985_7663# a_32334_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5768 VSS a_11067_67279# a_31726_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5769 VSS a_2411_19605# a_2369_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X577 VDD a_34711_47375# a_34987_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5770 VDD a_10515_22671# a_35346_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5771 a_22127_37737# a_22521_37692# a_20827_37737# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X5772 a_6473_62313# a_6417_62215# a_5497_63303# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X5773 a_45782_20902# a_11067_67279# a_45386_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5774 VDD a_12727_67753# a_18278_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5775 VDD a_12257_56623# a_48398_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5776 a_28810_24520# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5777 a_40762_69222# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5778 a_2203_66415# a_1757_66415# a_2107_66415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5779 a_18370_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X578 a_15097_51183# a_13925_51727# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X5780 a_14049_42869# a_13716_43047# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5781 a_37888_43983# a_37711_43983# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5782 VDD a_7162_60039# a_5749_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X5783 VSS a_1642_18231# a_1591_17999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5784 VSS a_19807_28111# a_32232_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X5785 a_35742_12870# a_10055_58791# a_35346_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5786 VDD a_18045_41281# a_18856_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5787 a_8497_54697# a_7479_54439# a_8082_54599# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X5788 a_50198_39208# a_49984_39288# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u M=8
X5789 VSS a_14983_51157# a_18034_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u M=4
X579 a_36520_42693# a_36392_43677# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X5790 a_7299_59887# a_7210_55081# a_7162_60039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5791 a_18674_22910# a_11067_21583# a_18278_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5792 vcm_commonmode a_16362_23548# a_42466_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5793 a_20286_70226# a_12516_7093# a_20778_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5794 a_41370_58178# a_16362_58178# a_41462_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5795 VDD a_12727_15529# a_22294_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5796 a_34359_50639# a_34411_50613# a_33360_51701# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X5797 VDD a_12707_26159# a_13059_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5798 a_18278_9858# a_16362_9492# a_18370_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5799 a_37939_43455# a_2021_22325# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X58 VDD a_12257_56623# a_49402_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X580 a_37446_20536# a_16746_20534# a_37354_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5800 a_6721_64239# a_6095_44807# a_6375_64489# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X5801 a_5803_74397# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X5802 a_29322_20902# a_12985_7663# a_29814_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5803 a_2509_47349# a_2291_47753# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X5804 a_44778_68218# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5805 a_29322_16886# a_16362_16520# a_29414_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5806 a_41370_17890# a_12899_10927# a_41862_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5807 VSS a_1645_42453# a_1593_42479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5808 a_30326_11866# a_16362_11500# a_30418_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5809 a_13975_34191# a_13798_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X581 a_26748_7638# a_30788_28487# a_30746_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X5810 a_11709_65569# a_11491_65327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X5811 a_48490_17524# a_16746_17522# a_48398_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5812 a_19282_12870# a_12877_16911# a_19774_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5813 VSS a_10791_15529# a_11714_14557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X5814 a_23790_10464# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5815 a_34738_18894# a_12899_10927# a_34342_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5816 VDD a_12725_44527# a_27891_41495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5817 VDD a_5411_59317# a_5333_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X5818 a_32426_22544# a_16746_22542# a_32334_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5819 a_8307_32687# a_6243_30662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X582 a_40458_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5820 vcm_commonmode a_16362_70226# a_41462_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5821 a_5411_12791# a_4429_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5822 VSS a_12727_67753# a_21686_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5823 a_47790_59182# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5824 VDD a_2292_43291# a_2592_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X5825 VSS a_22132_40865# a_21233_40956# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X5826 a_5136_34551# a_4495_35925# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5827 a_8361_15529# a_7987_15431# a_8289_15529# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5828 VSS a_10275_21495# a_10151_21379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X5829 a_45386_16886# a_12899_11471# a_45878_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X583 VDD a_12901_66665# a_18278_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5830 VDD a_40921_41245# a_40527_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5831 VDD a_27429_35301# a_28056_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5832 vcm_commonmode VSS a_19374_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5833 a_31726_64202# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5834 a_5447_56860# a_5291_56765# a_5592_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X5835 VSS a_30991_29397# a_27752_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5836 VDD a_4812_13879# a_6607_13879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5837 vcm_commonmode a_16362_13508# a_49494_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5838 VDD a_28441_36389# a_29068_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5839 a_5645_10383# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X584 VSS a_28757_27247# a_31127_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X5840 VDD a_19596_40743# a_19500_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X5841 VDD a_3295_54421# a_10975_55535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5842 a_44273_30287# a_41597_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5843 a_10697_72399# a_10509_73193# a_10615_72399# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5844 a_36442_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5845 a_7387_69929# a_6921_72943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X5846 VSS a_12877_14441# a_35742_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5847 a_23447_28853# a_18053_28879# a_23845_29245# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5848 a_33802_47375# a_33868_47349# a_33635_47695# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.8675e+11p ps=3.79e+06u w=650000u l=150000u
X5849 a_39854_7452# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X585 a_5483_74244# a_5779_75093# a_5737_75369# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5850 a_35742_7850# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5851 VSS a_12901_58799# a_24698_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5852 a_21686_56170# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5853 a_23593_35303# a_23901_35516# a_23567_35507# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5854 VSS a_6008_69679# a_6676_69455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5855 a_6263_15645# a_2292_17179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X5856 a_18278_18894# a_12895_13967# a_18770_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5857 VSS a_5447_56860# a_5378_56989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5858 a_22786_16488# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5859 VDD a_2223_28617# a_4065_24233# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X586 VDD a_11780_69679# a_11955_69653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5860 VDD a_12947_71576# a_39362_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5861 VDD VDD a_49402_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5862 VSS VDD a_45782_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5863 a_40366_67214# a_12983_63151# a_40858_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5864 a_26402_13508# a_16746_13506# a_26310_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5865 vcm_commonmode a_16362_10496# a_23390_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5866 a_22671_43439# a_1761_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X5867 a_39454_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5868 VSS a_28688_50247# a_28648_50101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5869 a_3112_19319# a_3143_22364# a_3254_19453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X587 a_40762_72234# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5870 a_11335_10076# a_11179_9981# a_11480_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X5871 vcm_commonmode a_16362_60186# a_48490_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5872 vcm_commonmode a_16362_19532# a_48490_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5873 VSS a_10515_22671# a_28714_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5874 a_25702_55166# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5875 a_38450_66210# a_16746_66212# a_38358_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5876 a_37577_42693# a_37885_42333# a_37551_42333# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X5877 a_26706_9858# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5878 a_9989_46831# a_9821_46831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X5879 a_40762_22910# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 a_2107_69513# a_1591_69141# a_2012_69501# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X5880 a_37354_21906# a_16362_21540# a_37446_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5881 VSS a_20881_28111# a_23303_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5882 VSS a_38436_29941# a_38969_29217# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5883 a_30875_36919# a_29943_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5884 a_11801_52047# a_11759_51959# a_9240_53877# VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X5885 a_5749_18297# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5886 VSS a_24800_35425# a_23901_35516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X5887 VDD a_15443_29941# a_14354_32117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5888 a_26310_68218# a_12727_67753# a_26802_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5889 a_43470_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X589 a_18370_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5890 a_30818_66532# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5891 VSS a_12899_10927# a_33734_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5892 a_25398_60186# a_16746_60188# a_25306_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5893 VDD a_12727_58255# a_29322_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5894 a_25398_19532# a_16746_19530# a_25306_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5895 a_14372_29429# a_13390_29575# a_14289_29687# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5896 a_30326_56170# a_16362_56170# a_30418_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5897 VSS config_1_in[12] a_1626_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5898 a_22448_37253# a_21479_36965# a_22352_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5899 a_44778_21906# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X59 a_20286_64202# a_16362_64202# a_20378_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X590 VSS a_12355_65103# a_39758_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5900 a_25300_38567# a_24331_38591# a_25263_38825# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X5901 VDD a_75162_40202# a_75111_40050# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5902 a_47394_57174# a_12257_56623# a_47886_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5903 a_11661_71855# a_11617_72097# a_11495_71855# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X5904 VSS a_28103_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5905 a_6909_41935# a_6269_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5906 VSS VDD a_42770_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5907 a_31330_62194# a_12355_15055# a_31822_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5908 a_13097_36367# a_12671_36694# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5909 a_34738_13874# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X591 a_4818_47414# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X5910 a_11022_48285# a_9945_47919# a_10860_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5911 a_16746_67216# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X5912 a_7199_62839# a_7077_62313# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X5913 a_7125_31375# a_2235_30503# a_6835_31055# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=2.34e+06u as=0p ps=0u w=650000u l=150000u
X5914 a_4647_63937# a_1586_66567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5915 vcm_commonmode VSS a_37446_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5916 a_17670_23914# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5917 a_47790_12870# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5918 VSS a_11067_21583# a_21686_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5919 a_30722_7850# VDD a_30326_7850# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X592 a_20612_37607# a_20827_37737# a_20754_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5920 a_18370_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5921 a_11082_14557# a_10956_14459# a_10678_14443# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X5922 a_33203_34191# a_33026_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X5923 a_24794_57496# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5924 VDD a_2939_33535# a_2926_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5925 VSS a_35431_31751# a_25787_28327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X5926 VDD a_28691_49783# a_28639_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X5927 vcm_commonmode a_16362_68218# a_38450_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5928 a_47486_7484# VDD a_47394_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5929 a_12621_59343# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X593 a_32334_65206# a_12355_65103# a_32826_65528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5930 a_30843_52521# a_2959_47113# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X5931 VSS a_77285_39738# a_77098_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5932 VSS a_5147_50943# a_5081_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X5933 a_26465_48463# a_26187_48801# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5934 VDD a_2787_32679# a_6069_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5935 a_38454_34191# a_38277_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5936 a_7289_62607# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5937 a_27710_15882# a_12877_14441# a_27314_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5938 VSS a_12877_16911# a_24698_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5939 VSS a_12981_62313# a_36746_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 VDD a_12899_11471# a_39362_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5940 a_20904_30761# a_5363_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X5941 a_16744_41605# a_15775_41317# a_16648_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X5942 vcm_commonmode a_16362_9492# a_28410_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5943 VSS a_4351_26703# a_8369_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5944 a_7917_12265# a_7841_12167# a_7799_12265# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5945 VSS a_1761_31055# a_32327_35839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X5946 VSS a_12355_15055# a_49798_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5947 VDD a_12687_34191# a_12793_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5948 a_45478_57174# a_16746_57176# a_45386_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5949 a_22294_7850# VSS a_22386_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X595 a_6921_72943# a_5599_74549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X5950 a_46786_18894# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5951 a_4417_22671# a_4083_22351# a_4333_22351# VDD sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X5952 VDD a_6059_14165# a_5943_15492# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X5953 a_19492_52245# a_4758_45369# a_19715_52271# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X5954 VSS a_28747_37503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X5955 a_2629_54447# a_2250_54813# a_2557_54447# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5956 VSS a_2595_47653# a_4669_51005# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5957 VDD a_11659_66567# a_9513_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5958 vcm_commonmode a_16362_18528# a_24394_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5959 a_34834_22512# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X596 a_6444_16367# a_5363_16367# a_6097_16609# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X5960 a_28810_58500# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5961 a_32426_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5962 a_2746_16885# a_2596_16911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.184e+11p pd=2.2e+06u as=0p ps=0u w=840000u l=150000u
X5963 VSS a_10055_58791# a_28714_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5964 a_41462_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5965 VSS a_4417_22671# a_8377_24847# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X5966 a_12381_35836# a_32003_35307# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5967 VDD a_14831_50095# a_29829_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X5968 a_21290_71230# a_16362_71230# a_21382_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5969 a_26706_62194# a_12981_62313# a_26310_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X597 a_37446_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5970 VDD a_2511_42479# a_2292_43291# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X5971 VDD a_3357_67257# a_3387_66998# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5972 a_11763_62581# a_11943_63125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5973 VDD a_1923_54591# a_1643_57685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5974 a_4149_48469# a_3983_48469# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5975 a_1846_63403# a_2163_63293# a_2121_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X5976 a_38358_72234# VDD a_38850_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5977 a_38850_21508# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5978 a_38450_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5979 a_42866_70548# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X598 VDD a_33694_30761# a_33797_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5980 a_35346_14878# a_16362_14512# a_35438_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5981 a_6095_54697# a_5531_53903# a_5877_54421# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5982 a_42374_60186# a_16362_60186# a_42466_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5983 a_17830_49373# a_16753_49007# a_17668_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X5984 VDD a_28361_51701# a_28251_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X5985 VDD a_10244_26159# a_10472_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X5986 a_25306_70226# a_16362_70226# a_25398_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5987 VDD a_12047_57685# a_12034_58077# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X5988 VDD a_12985_16367# a_32334_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5989 a_18840_47375# a_18626_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X599 a_22181_50645# a_22015_50645# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X5990 a_17670_64202# a_12355_65103# a_17274_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5991 VSS a_5594_36727# a_5547_36495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5992 VDD a_12875_31751# a_12215_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X5993 a_30716_51701# a_2775_46025# a_30845_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X5994 a_10589_10383# a_9484_11989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5995 VDD config_1_in[14] a_1591_22895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X5996 a_39459_44527# a_39282_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X5997 a_39362_13874# a_16362_13508# a_39454_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5998 VDD a_12546_22351# a_45386_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X5999 a_27155_40871# a_27263_40871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_42466_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.957e+14p ps=2.64812e+09u w=800000u l=150000u
X60 a_29814_24520# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X600 a_4060_70223# a_3372_70197# a_3452_70537# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6000 a_42283_42359# a_41351_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6001 a_6435_10901# a_6260_10927# a_6614_10927# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6002 VDD a_28717_42917# a_29205_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6003 a_18370_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6004 VSS a_1950_59887# a_10189_60797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6005 a_36746_67214# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6006 a_17797_40517# a_18105_40157# a_13576_40413# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X6007 VDD a_11067_67279# a_28318_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6008 a_31117_28879# a_20635_29415# a_31117_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6009 a_20661_49917# a_20282_49551# a_20589_49917# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X601 VSS a_5239_20693# a_3987_19623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X6010 a_43774_68218# a_12901_66959# a_43378_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6011 VSS a_12355_65103# a_40762_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6012 VDD a_2411_18517# a_11480_10205# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6013 a_28318_61190# a_16362_61190# a_28410_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6014 VSS a_11763_57399# a_11080_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6015 vcm_commonmode a_16362_56170# a_44474_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6016 a_2012_39037# a_1895_38842# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6017 vcm_commonmode a_16362_21540# a_38450_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6018 a_5211_24759# a_8625_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=6
X6019 a_1761_52815# a_1591_52815# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X602 VDD a_77568_40202# a_77381_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6020 VDD a_10055_58791# a_18278_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6021 VSS a_38210_30199# a_38239_32375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6022 vcm_commonmode a_16362_66210# a_27406_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6023 VDD a_14831_50095# a_32310_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X6024 a_16362_13508# a_11067_23759# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X6025 a_14809_47919# a_5039_42167# a_14737_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6026 a_31422_64202# a_16746_64204# a_31330_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6027 a_3254_9661# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6028 a_29322_24918# VSS a_29414_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6029 a_1683_5059# a_1681_5175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X603 a_22294_57174# a_12257_56623# a_22786_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6030 VDD a_19459_29423# a_19626_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6031 a_36842_63520# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6032 a_40394_28585# a_32823_29397# a_40086_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.25e+11p pd=2.65e+06u as=0p ps=0u w=1e+06u l=150000u
X6033 a_46786_59182# a_12727_58255# a_46390_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6034 VDD a_12355_15055# a_40366_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6035 a_29414_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6036 VDD a_12815_19319# a_12815_19087# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X6037 VDD a_12727_13353# a_44382_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6038 a_21879_30663# a_14646_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6039 a_29718_69222# a_12516_7093# a_29322_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X604 VDD a_16928_35303# a_16832_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X6040 a_21382_56170# a_16746_56172# a_21290_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6041 a_22690_17890# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6042 a_8543_36469# a_8902_36469# a_8679_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X6043 a_45478_10496# a_16746_10494# a_45386_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6044 a_22062_31287# a_2787_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6045 a_4972_51017# a_3891_50645# a_4625_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6046 a_43678_31029# a_43680_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X6047 a_35932_41953# a_35647_41317# a_36579_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X6048 VSS a_11069_23983# a_11163_25321# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6049 a_1849_31599# a_1683_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X605 a_33734_55166# a_12869_2741# a_33338_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6050 a_45386_67214# a_16362_67214# a_45478_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6051 VSS VSS a_47790_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6052 a_26273_48801# a_6835_46823# a_26187_48801# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6053 a_15925_30287# a_3339_30503# a_15829_30287# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X6054 a_31726_72234# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6055 VSS a_12139_71829# a_5877_70197# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6056 a_35838_69544# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6057 a_24302_10862# a_16362_10496# a_24394_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6058 a_35346_59182# a_16362_59182# a_35438_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6059 VSS a_2847_9813# a_1929_10651# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X606 a_8375_40847# a_8384_40303# a_8017_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X6060 a_33727_38825# a_33764_38567# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6061 a_13762_41046# a_13067_38517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X6062 a_11710_58487# a_12407_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6063 a_20161_48463# a_19991_48463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6064 a_18278_69222# a_16362_69222# a_18370_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6065 VDD a_1689_10396# a_1633_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6066 VDD a_12981_62313# a_17274_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6067 a_7802_45199# a_6725_45205# a_7640_45577# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6068 VDD a_8273_42479# a_9445_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6069 a_22386_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X607 VSS a_13143_29575# a_14444_29429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X6070 a_24698_55166# VSS a_24302_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6071 a_2012_15101# a_1895_14906# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6072 VDD a_4032_53047# a_3231_53047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6073 VDD a_3355_25071# a_4351_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6074 a_36350_65206# a_12355_65103# a_36842_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6075 VSS a_26631_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X6076 a_37830_28111# a_37527_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X6077 a_39362_58178# a_16362_58178# a_39454_58178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6078 a_25702_63198# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6079 a_5173_61225# a_4985_61021# a_5091_60981# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X608 a_32730_20902# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6080 vcm_commonmode a_16362_58178# a_21382_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6081 vcm_commonmode a_16362_71230# a_35438_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6082 a_21616_43781# a_20743_43493# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6083 a_1846_63403# a_2124_63419# a_2080_63517# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6084 a_33760_40743# a_32887_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6085 a_39362_17890# a_12899_10927# a_39854_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6086 VSS a_12947_23413# a_39758_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6087 a_7001_36495# a_6653_36611# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6088 a_36746_20902# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6089 a_25313_31599# a_24746_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X609 a_2012_33927# a_4503_21523# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X6090 a_32867_28879# a_33008_28853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6091 a_4437_34639# a_2011_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6092 a_15315_52271# a_7050_53333# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=0p ps=0u w=650000u l=150000u M=2
X6093 a_43870_15484# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6094 a_43774_21906# a_12985_7663# a_43378_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6095 a_9869_67745# a_9651_67503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6096 a_40366_12870# a_12877_16911# a_40858_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6097 a_9945_73807# a_8003_72917# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X6098 a_4918_58255# a_4792_58371# a_4514_58387# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6099 a_14049_36341# a_13123_38231# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X61 a_41766_69222# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X610 a_44474_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6100 a_24029_39355# a_35647_40229# a_36520_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6101 VDD a_10515_22671# a_46390_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6102 a_23298_22910# a_10515_23975# a_23790_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6103 VSS a_12546_22351# a_36746_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6104 a_16362_58178# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X6105 VDD a_10515_23975# a_30326_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6106 a_2835_23222# a_1689_10396# a_2376_23047# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X6107 VDD a_12727_67753# a_29322_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6108 a_2805_22869# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6109 VDD a_32029_41829# a_33484_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X611 VSS a_12901_66665# a_30722_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6110 a_11893_65871# a_11521_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X6111 vcm_commonmode a_16362_70226# a_39454_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6112 a_30326_64202# a_16362_64202# a_30418_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6113 a_33734_13874# a_12877_16911# a_33338_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6114 VDD a_4443_46607# a_8367_44343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6115 a_9263_24501# a_7377_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6116 a_29414_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6117 VDD a_13957_36121# a_13987_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6118 a_29620_37479# a_28747_37503# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6119 vcm_commonmode VSS a_40458_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X612 a_4220_57685# a_4482_57863# a_4440_57711# VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6120 a_2150_17289# a_1757_16917# a_2040_17289# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X6121 a_46786_9858# a_12985_19087# a_46390_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6122 VDD a_23467_41237# a_23415_41263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6123 VDD a_12877_14441# a_20286_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6124 a_46786_12870# a_10055_58791# a_46390_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6125 a_44382_11866# a_10055_58791# a_44874_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6126 a_2100_24759# a_2223_28617# a_2242_24893# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6127 a_29718_64202# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6128 a_34342_68218# a_12727_67753# a_34834_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6129 a_29718_22910# a_11067_21583# a_29322_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X613 VDD a_12985_16367# a_44382_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6130 a_27314_21906# a_11067_21583# a_27806_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6131 a_15207_30511# a_14361_29967# a_15986_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u M=2
X6132 a_27314_17890# a_16362_17524# a_27406_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6133 a_2369_15101# a_2325_14709# a_2203_15113# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6134 a_31330_70226# a_12516_7093# a_31822_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6135 a_33430_60186# a_16746_60188# a_33338_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6136 VDD a_12727_58255# a_37354_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6137 a_33430_19532# a_16746_19530# a_33338_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6138 a_31422_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6139 a_16362_70226# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X614 a_28817_29111# a_38883_29217# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6140 a_23911_35823# a_23734_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6141 a_19678_56170# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6142 a_46482_18528# a_16746_18526# a_46390_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6143 a_8753_66103# a_8958_65961# a_8916_65987# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6144 vcm_commonmode a_16362_15516# a_43470_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6145 a_17274_13874# a_12727_15529# a_17766_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6146 a_28056_40517# a_28152_40517# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6147 a_5169_29673# a_4497_29673# a_5087_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6148 VDD a_10513_48161# a_10403_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6149 a_2012_49917# a_1895_49722# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X615 VSS a_1915_35015# a_3803_35523# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X6150 a_21782_11468# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6151 VDD a_1959_26703# a_2099_59861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X6152 a_30091_35253# a_30267_35253# a_30219_35279# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X6153 a_30418_23548# a_16746_23546# a_30326_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6154 VDD a_2292_17179# a_2596_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X6155 a_12231_65301# a_12056_65327# a_12410_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6156 a_11865_24527# a_9955_20969# a_11793_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X6157 a_1644_63669# a_1823_63677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6158 a_18497_47741# a_17787_47349# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6159 a_4987_52508# a_4792_52539# a_5297_52271# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X616 a_6361_57711# a_5823_57961# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6160 a_19374_61190# a_16746_61192# a_19282_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6161 a_12123_46831# a_11067_47695# a_11760_46983# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6162 VSS a_11067_23759# a_16362_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X6163 VDD a_30912_39429# a_30816_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X6164 VSS a_12727_67753# a_32730_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6165 a_20378_15516# a_16746_15514# a_20286_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6166 a_1945_43023# a_1593_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=0p ps=0u w=840000u l=150000u
X6167 vcm_commonmode a_16362_14512# a_47486_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6168 a_52778_39936# a_52590_39936# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.66e+06u as=0p ps=0u w=500000u l=150000u M=2
X6169 VSS a_1689_10396# a_1633_12342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X617 a_5169_13353# a_5399_13255# a_5023_13255# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X6170 VSS a_7939_30503# a_25605_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6171 a_7125_46653# a_7090_46419# a_6655_46261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6172 a_27167_32509# a_5363_30503# a_27417_32509# VSS sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X6173 a_43378_19898# a_11067_67279# a_43870_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6174 a_19026_31375# a_13353_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6175 a_19774_8456# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6176 a_2283_32362# a_2235_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6177 a_39372_37479# a_38499_37503# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6178 VSS a_28959_49783# a_28909_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X6179 a_47486_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X618 a_33668_38341# a_32795_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6180 a_40762_71230# a_12947_71576# a_40366_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6181 a_38450_9492# a_16746_9490# a_38358_9858# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6182 VDD a_4571_26677# a_7267_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6183 a_28810_66532# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6184 a_25306_63198# a_12981_62313# a_25798_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6185 VSS a_36392_43677# a_35493_43421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X6186 a_5616_43567# a_4701_43567# a_5269_43809# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6187 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X6188 VDD a_12947_8725# a_29322_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6189 VSS a_12985_19087# a_25702_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X619 a_29718_64202# a_12355_65103# a_29322_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6190 a_24394_14512# a_16746_14510# a_24302_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6191 vcm_commonmode a_16362_11500# a_21382_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6192 a_5043_19306# a_5135_19061# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X6193 VSS a_7479_57175# a_6515_62037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6194 a_14287_51175# a_30440_31573# a_30021_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X6195 a_37446_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6196 a_30520_50345# a_27869_50095# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6197 a_20778_19500# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6198 VSS a_77285_40202# a_77098_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6199 VDD a_12257_56623# a_22294_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X62 VDD a_1586_21959# a_10883_18007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X620 a_32779_27497# a_20359_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X6200 a_36442_67214# a_16746_67216# a_36350_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6201 a_12689_55311# a_12659_54965# a_12605_55311# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X6202 a_18977_27791# a_18126_28023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6203 a_14049_36341# a_13123_38231# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6204 VSS a_7162_59575# a_6382_61127# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6205 a_29322_62194# a_12355_15055# a_29814_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6206 VSS a_4528_26159# a_5087_24643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6207 a_35346_22910# a_16362_22544# a_35438_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6208 a_1586_40455# a_4535_43031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6209 a_4343_60405# a_4148_60547# a_4653_60797# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X621 VDD a_12901_66959# a_34342_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6210 a_49494_66210# a_16746_66212# a_49402_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6211 VSS a_21479_42405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X6212 VDD a_17222_27247# a_22808_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X6213 a_48398_21906# a_16362_21540# a_48490_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6214 a_19071_28111# a_17222_27247# a_18977_28111# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X6215 a_10299_20969# a_6816_19355# a_9872_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X6216 a_17670_72234# VDD a_17274_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6217 a_12981_59343# a_12712_59343# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6218 a_47790_61190# a_12355_15055# a_47394_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6219 VSS a_12899_10927# a_44778_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X622 VSS a_11067_46823# a_40783_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6220 VDD a_5135_50069# a_5909_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6221 a_8206_28879# a_5087_29423# a_8206_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X6222 a_5595_12167# a_1929_10651# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6223 a_23271_50943# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6224 a_25398_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6225 vcm_commonmode a_16362_8488# a_41462_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6226 a_2775_46025# a_2847_45503# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X6227 a_19446_51183# a_19946_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X6228 VDD a_26523_29199# a_43680_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6229 VSS a_4215_51157# a_27167_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X623 a_28855_48801# a_26514_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6230 a_9557_64757# a_9280_65327# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X6231 vcm_commonmode a_16362_8488# a_17366_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6232 a_38959_29967# a_35815_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6233 a_6769_40125# a_4314_40821# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6234 a_38209_30761# a_33694_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X6235 a_31000_38341# a_30127_38053# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6236 a_21686_17890# a_12899_11471# a_21290_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6237 a_2107_69513# a_1757_69141# a_2012_69501# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X6238 VSS a_12899_11471# a_48794_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6239 a_45782_13874# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_22690_12870# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6240 a_40402_28111# a_40457_27765# a_40233_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X6241 a_31422_72234# VDD a_31330_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6242 a_46482_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6243 a_36842_71552# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6244 a_28714_23914# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6245 a_11449_62313# a_11395_62037# a_9643_63125# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6246 a_27406_8488# a_16746_8486# a_27314_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6247 a_32334_15882# a_12727_13353# a_32826_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6248 VSS a_11067_21583# a_32730_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6249 a_29414_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X625 a_75475_38962# a_75199_38962# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6250 a_21948_34973# a_21479_34239# a_22352_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6251 a_3026_18543# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X6252 a_16746_13506# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X6253 VDD a_2686_70223# a_4181_73193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6254 a_19282_71230# a_16362_71230# a_19374_71230# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6255 a_49402_59182# a_12901_58799# a_49894_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6256 a_36629_27791# a_36459_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6257 a_18674_15882# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6258 a_5803_11293# a_5179_10927# a_5695_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6259 VDD a_4312_19061# a_1586_9991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X626 a_34738_63198# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6260 a_25702_16886# a_12727_13353# a_25306_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6261 VSS a_12727_15529# a_22690_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6262 VSS a_43321_29941# a_43269_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6263 VSS a_37551_42333# a_37491_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6264 a_2928_67191# a_1770_14441# a_3070_67325# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6265 VSS a_12981_62313# a_47790_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6266 VSS a_4427_30511# a_6099_23983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6267 a_15681_27247# a_12349_25847# a_15871_27247# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X6268 a_5239_45717# a_5064_45743# a_5418_45743# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6269 VSS a_52778_39198# a_19967_41781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X627 a_33041_51157# a_33313_51157# a_33712_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u M=2
X6270 a_37750_69222# a_12516_7093# a_37354_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6271 VSS a_11659_66567# a_11764_65845# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X6272 VSS a_3339_43023# a_7757_21379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6273 a_8475_44343# a_8143_44982# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6274 VSS a_10975_66407# a_34738_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6275 a_2317_28892# a_2847_21781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6276 vcm_commonmode a_16362_60186# a_22386_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6277 a_26802_59504# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6278 vcm_commonmode a_16362_19532# a_22386_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6279 a_26671_50095# a_26321_50095# a_26576_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X628 VDD a_9669_26703# a_11251_26159# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6280 a_5906_28585# a_5073_27247# a_5823_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X6281 a_36442_20536# a_16746_20534# a_36350_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6282 a_45878_22512# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6283 a_12713_36483# a_24515_34789# a_25447_34743# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X6284 a_3595_73487# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6285 VDD a_12901_66665# a_17274_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6286 a_35438_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6287 a_24698_63198# a_15439_49525# a_24302_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6288 VDD a_23051_28023# a_22762_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6289 a_10423_30761# a_6459_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X629 VSS a_28691_49783# a_28639_49551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6290 VSS a_12355_65103# a_38754_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6291 VSS a_19096_44129# a_19559_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X6292 VDD a_11710_58487# a_11893_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6293 VDD a_12899_11471# a_38358_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6294 VDD a_8857_14709# a_8747_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6295 a_35838_14480# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6296 a_30561_48829# a_14831_50095# a_30479_48576# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6297 a_3509_58487# a_3618_58487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6298 a_2150_28662# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X6299 a_36442_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X63 a_19374_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X630 a_47790_62194# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6300 VSS a_21049_41245# a_20741_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6301 a_17044_28335# a_12985_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6302 a_49894_21508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6303 a_49494_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6304 a_46390_14878# a_16362_14512# a_46482_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6305 VSS a_2747_72007# a_2571_72040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6306 a_32730_55166# a_11067_47695# a_32334_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6307 a_13381_38365# a_13111_37999# a_13291_37999# VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6308 VSS a_6619_16341# a_5535_18012# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X6309 VSS a_19807_28111# a_35079_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X631 vcm_commonmode a_16362_57174# a_43470_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6310 a_17869_28585# a_15799_29941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6311 a_30762_49641# a_30520_50345# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6312 VSS a_38327_44759# a_38140_44501# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6313 a_43470_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6314 a_30219_35279# a_13097_36367# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6315 VDD a_10472_54135# a_9547_54421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6316 a_39854_13476# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6317 a_36350_10862# a_12985_16367# a_36842_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6318 VSS a_35815_31751# a_21187_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6319 a_27422_29789# a_5363_30503# a_26221_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 VSS a_2292_17179# a_2369_15101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6320 VDD a_29926_30511# a_30939_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6321 a_32772_7638# a_30788_28487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6322 VDD a_12985_16367# a_43378_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6323 a_15146_27907# a_14471_28585# a_15064_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6324 a_4406_73853# a_1923_73087# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6325 a_28714_64202# a_12355_65103# a_28318_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6326 VSS a_15074_50871# a_14681_50247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6327 VSS a_11763_21237# a_11480_23957# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6328 VDD a_12901_66959# a_33338_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6329 a_4263_32259# a_2216_28309# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X633 VSS a_3143_22364# a_3985_22901# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6330 VDD a_12985_7663# a_26310_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6331 a_26310_9858# a_12546_22351# a_26802_9460# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6332 VSS a_23789_39100# a_23733_39126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6333 VSS a_9624_65301# a_9543_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.355e+11p ps=3.94e+06u w=650000u l=150000u
X6334 VDD a_31084_30485# a_21371_52263# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6335 VSS a_17039_51157# a_18257_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6336 a_29414_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6337 a_26310_62194# a_16362_62194# a_26402_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6338 a_41141_28879# a_34759_31029# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6339 a_2163_57853# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X634 VSS a_3325_18543# a_5265_28157# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X6340 a_30418_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6341 vcm_commonmode a_16362_57174# a_42466_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6342 a_18674_56170# a_12257_56623# a_18278_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6343 a_29718_72234# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6344 vcm_commonmode a_16362_67214# a_25398_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6345 a_2163_56765# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6346 VSS a_34759_31029# a_40961_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X6347 VDD a_6619_73719# a_6098_73095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X6348 a_5081_51017# a_3891_50645# a_4972_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6349 VDD a_12727_67753# a_37354_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X635 a_19678_56170# a_12257_56623# a_19282_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6350 a_34834_64524# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6351 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X6352 VDD a_10055_58791# a_29322_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6353 a_31422_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6354 a_27406_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6355 VSS a_26020_30199# a_25971_29967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6356 a_47886_63520# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6357 VSS a_12355_15055# a_23694_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6358 a_22995_30663# a_3339_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6359 a_20682_18894# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X636 vcm_commonmode a_16362_67214# a_26402_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6360 a_8491_41383# a_14298_32143# a_15162_32463# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X6361 VSS a_6459_30511# a_14013_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6362 a_2773_4943# a_2603_4943# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X6363 a_37750_22910# a_11067_21583# a_37354_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6364 VDD a_7571_29199# a_20993_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X6365 a_28056_35077# a_27183_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6366 a_32426_56170# a_16746_56172# a_32334_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6367 a_33734_17890# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6368 a_9927_60809# a_9577_60437# a_9832_60797# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X6369 a_9123_57399# a_9135_56623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X637 a_1757_26159# a_1591_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6370 a_35346_60186# a_12727_58255# a_35838_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6371 a_3805_30083# a_3325_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6372 a_29068_35303# a_28195_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6373 VDD a_7189_35015# a_5963_36585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X6374 a_48794_8854# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6375 a_13620_40871# a_13835_41001# a_13762_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X6376 a_43378_68218# a_16362_68218# a_43470_68218# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6377 VDD a_15439_49525# a_24302_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6378 vcm_commonmode a_16362_58178# a_19374_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6379 VSS a_16087_31751# a_15911_31784# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X638 a_30418_65206# a_16746_65208# a_30326_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6380 a_1761_39215# a_1591_39215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X6381 VDD a_23567_35507# a_23593_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6382 VSS a_12381_35836# a_26495_35253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6383 a_1757_16917# a_1591_16917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6384 a_42801_27497# a_41842_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6385 a_24561_41583# a_14293_41807# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X6386 VDD a_38171_34191# a_38277_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6387 a_2150_28335# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6388 a_25306_71230# a_12901_66665# a_25798_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6389 a_46390_59182# a_16362_59182# a_46482_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X639 VDD a_3541_19385# a_3571_19126# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6390 a_9872_20175# a_4792_20443# a_10131_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X6391 a_20378_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6392 VDD a_30788_28487# a_33591_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.25e+11p ps=2.85e+06u w=1e+06u l=150000u
X6393 VDD a_11067_67279# a_12727_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X6394 a_2107_18543# a_1591_18543# a_2012_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X6395 VDD a_12981_62313# a_28318_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6396 a_49798_69222# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6397 a_8935_27791# a_8662_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6398 a_12473_36341# a_31819_35073# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6399 VDD a_37551_42333# a_37577_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X64 a_28361_51701# a_28143_52105# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X640 a_11074_22895# a_11130_22869# a_11067_47695# VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X6400 a_9301_49557# a_9135_49557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6401 a_1846_56875# a_2124_56891# a_2080_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6402 a_35742_8854# a_12947_8725# a_35346_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6403 VSS a_13909_39747# a_39055_39913# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6404 a_9223_22895# a_4798_23759# a_9223_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=4.1e+11p ps=2.82e+06u w=1e+06u l=150000u
X6405 VDD a_8273_42479# a_9367_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6406 a_10145_60405# a_9927_60809# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X6407 a_29322_70226# a_12516_7093# a_29814_70548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6408 a_22531_51017# a_22015_50645# a_22436_51005# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X6409 VSS a_12901_58799# a_43774_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X641 a_2215_29967# a_1591_29973# a_2107_30345# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X6410 a_40762_56170# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6411 a_37354_18894# a_12895_13967# a_37846_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6412 VSS VSS a_37750_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6413 VDD a_3247_20495# a_4842_45467# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6414 a_2012_49917# a_1895_49722# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6415 vcm_commonmode a_16362_71230# a_46482_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6416 a_41862_16488# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6417 VSS a_12901_66959# a_26706_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6418 a_23694_66210# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6419 VSS a_37520_49783# a_36464_49783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X642 VSS a_35647_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X6420 a_30722_67214# a_12727_67753# a_30326_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6421 VDD a_4792_20443# a_12821_20175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6422 a_21290_23914# a_12947_23413# a_21782_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6423 a_21290_19898# a_16362_19532# a_21382_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6424 vcm_commonmode a_16362_10496# a_42466_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6425 VDD a_1803_20719# a_1945_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6426 VDD a_35403_50069# a_34579_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6427 VSS a_2847_18517# a_2781_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6428 a_28410_23548# a_16746_23546# a_28318_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6429 vcm_commonmode a_16362_20536# a_25398_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X643 VDD a_12727_67753# a_38358_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6430 a_34251_52263# a_35263_28879# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=150000u
X6431 VDD a_27337_38565# a_27320_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6432 a_8082_54599# a_8199_58229# a_8219_54447# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X6433 a_9653_69831# a_9314_69367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6434 a_40458_61190# a_16746_61192# a_40366_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6435 a_27406_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6436 a_20682_59182# a_12727_58255# a_20286_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6437 a_44778_55166# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6438 a_44778_13874# a_12877_16911# a_44382_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6439 a_7107_40847# a_6927_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X644 a_35838_64524# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6440 a_30679_43493# a_29913_43457# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X6441 a_27710_65206# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6442 a_5091_60981# a_3295_62083# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6443 a_18370_15516# a_16746_15514# a_18278_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6444 a_27806_17492# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6445 a_42985_46831# a_20267_30503# a_42997_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X6446 VDD a_12877_14441# a_31330_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6447 a_25306_18894# a_16362_18528# a_25398_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6448 a_37446_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6449 VDD a_25939_51157# a_25926_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X645 a_30021_31599# a_28757_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.085e+11p pd=7.38e+06u as=0p ps=0u w=650000u l=150000u M=2
X6450 a_5795_27497# a_4248_29967# a_5639_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.8525e+11p pd=1.87e+06u as=5.6875e+11p ps=5.65e+06u w=650000u l=150000u
X6451 a_9789_73807# a_9353_72399# a_9707_73807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6452 a_4717_65569# a_4499_65327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X6453 a_45386_68218# a_12727_67753# a_45878_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6454 a_44474_60186# a_16746_60188# a_44382_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6455 a_17670_57174# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6456 a_44474_19532# a_16746_19530# a_44382_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6457 VDD a_12727_58255# a_48398_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6458 vcm_commonmode a_16362_16520# a_41462_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6459 a_12703_38517# a_12879_38517# a_12831_38543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.008e+11p ps=1.32e+06u w=420000u l=150000u
X646 a_32426_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6460 VSS VSS a_21686_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6461 VDD a_1586_45431# a_4535_43031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6462 a_27406_70226# a_16746_70228# a_27314_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6463 a_33430_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6464 a_7622_61839# a_7580_61751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6465 a_32334_66210# a_16362_66210# a_32426_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6466 vcm_commonmode a_16362_11500# a_19374_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6467 VSS a_26523_29199# a_43495_28487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6468 a_28318_13874# a_12727_15529# a_28810_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6469 a_32826_11468# a_32772_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X647 a_2629_63151# a_2250_63517# a_2557_63151# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6470 a_18770_19500# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6471 VDD VDD a_18278_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6472 VDD a_2511_23983# a_2411_19605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6473 a_22786_68540# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6474 a_30326_7850# VDD a_30818_7452# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6475 a_38784_42589# a_38499_42943# a_39372_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6476 a_49402_67214# a_12983_63151# a_49894_67536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6477 a_17366_62194# a_16746_62196# a_17274_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6478 a_11902_27497# a_7369_24233# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6479 a_13005_43983# a_12579_44310# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X648 a_19885_50095# a_19715_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6480 a_22762_27791# a_4811_34855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6481 VSS a_3799_31063# a_2473_34293# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6482 a_6641_37903# a_5993_37039# a_6559_37583# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6483 a_24698_7850# VDD a_24302_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6484 a_18379_46831# a_3339_32463# a_18016_46983# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6485 VDD a_1803_20719# a_32327_40191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6486 a_18445_46805# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6487 a_18626_47375# a_18539_47617# a_18222_47507# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6488 a_43870_57496# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6489 a_49798_22910# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X649 a_38450_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6490 a_4681_13621# a_4057_13647# a_4968_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6491 a_26802_67536# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6492 a_23298_64202# a_11067_13095# a_23790_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6493 VDD a_10975_66407# a_30326_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6494 a_25450_28995# a_9529_28335# a_25368_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6495 VDD a_23731_28023# a_23051_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X6496 VSS a_4227_73791# a_4161_73865# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6497 a_35438_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6498 VSS a_12877_16911# a_43774_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6499 VDD a_10515_22671# a_20286_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X65 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u M=777
X650 a_20282_49551# a_20156_49667# a_19878_49683# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6500 VSS a_7295_44647# a_40233_31605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6501 a_16270_7850# VSS a_16362_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6502 VSS a_10515_23975# a_26706_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6503 a_35742_70226# a_34251_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6504 a_19780_39429# a_18811_39141# a_19743_39095# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X6505 a_34434_68218# a_16746_68220# a_34342_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6506 a_30722_20902# a_11067_67279# a_30326_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6507 VSS config_1_in[2] a_1591_11471# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6508 VDD a_13390_29575# a_14289_29687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5795e+11p ps=2.99e+06u w=420000u l=150000u
X6509 a_33697_50359# a_33826_50075# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X651 a_7009_72105# a_6271_72943# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.05e+11p pd=2.61e+06u as=0p ps=0u w=1e+06u l=150000u
X6510 a_49876_37608# ctopp a_50198_39208# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=9.32e+06u as=0p ps=0u w=2e+06u l=150000u M=4
X6511 a_47486_67214# a_16746_67216# a_47394_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6512 a_2250_58077# a_2124_57979# a_1846_57963# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6513 a_12579_44310# a_12621_44099# a_12579_43983# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X6514 a_46390_22910# a_16362_22544# a_46482_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6515 a_12196_21583# a_5535_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.6875e+11p pd=4.35e+06u as=0p ps=0u w=650000u l=150000u
X6516 a_20682_12870# a_10055_58791# a_20286_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6517 a_10680_52245# a_32582_51701# VSS VSS sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u M=4
X6518 a_32730_63198# a_15439_49525# a_32334_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6519 VDD a_12663_39783# a_12651_39997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X652 VSS a_12907_56399# a_16362_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X6520 a_17274_55166# VSS a_17766_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6521 a_40458_7484# VDD a_40366_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6522 a_11902_27247# a_7369_24233# a_12092_27247# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u M=2
X6523 VSS a_18016_46983# a_17311_46833# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6524 a_38754_61190# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6525 a_37446_59182# a_16746_59184# a_37354_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6526 a_40366_71230# a_16362_71230# a_40458_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6527 a_45782_62194# a_12981_62313# a_45386_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6528 a_1757_69141# a_1591_69141# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6529 VSS a_12895_13967# a_42770_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X653 VSS a_12355_15055# a_24698_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6530 a_39685_27791# a_37699_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X6531 a_16362_7484# VDD a_16270_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6532 a_12757_8207# a_12479_8545# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X6533 a_28714_72234# VDD a_28318_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6534 VDD a_5535_18012# a_10394_19605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X6535 a_22631_29199# a_22577_29111# a_22441_28879# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X6536 a_17670_10862# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6537 vcm_commonmode a_16362_9492# a_21382_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6538 a_6921_20969# a_2339_38129# a_6825_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6539 a_5447_56860# a_5252_56891# a_5757_56623# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X654 a_7162_60039# a_6559_59879# a_7299_59887# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X6540 a_4807_27613# a_4627_27613# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6541 a_2104_33597# a_1987_33402# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6542 VSS a_28152_44869# a_28115_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6543 a_15661_29199# a_10506_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=2
X6544 a_8453_51727# a_8051_52047# a_8289_52047# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X6545 vcm_commonmode VSS a_38450_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6546 a_44382_70226# a_16362_70226# a_44474_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6547 a_43774_14878# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6548 a_36842_9460# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6549 VSS a_77002_39738# a_76744_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X655 a_20378_57174# a_16746_57176# a_20286_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6550 a_32730_59182# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6551 a_34834_72556# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6552 a_26706_24918# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6553 a_30326_16886# a_12899_11471# a_30818_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6554 VDD a_1689_10396# a_1863_42729# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X6555 VDD a_12985_19087# a_46390_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6556 a_34342_62194# a_16362_62194# a_34434_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6557 VDD a_12981_59343# a_34342_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6558 a_2104_31599# a_1987_31812# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X6559 a_4726_20541# a_3247_20495# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X656 VSS a_4083_22351# a_4417_22671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.005e+11p ps=2.84e+06u w=650000u l=150000u
X6560 a_49750_39288# a_42165_36367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6561 a_47886_71552# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6562 a_2847_12863# a_2672_12937# a_3026_12925# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6563 VDD a_11067_67279# a_47394_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6564 a_17274_72234# VSS a_17366_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6565 VSS a_12727_58255# a_19678_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6566 VSS a_11067_67279# a_19678_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6567 a_21382_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6568 a_47394_61190# a_16362_61190# a_47486_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6569 VSS a_12877_14441# a_20682_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X657 a_21686_18894# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6570 a_21479_34239# a_19596_34215# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X6571 VDD a_5024_67885# a_6825_66665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6572 a_2203_39049# a_1757_38677# a_2107_39049# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X6573 VSS config_2_in[11] a_1591_46287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6574 VDD a_10055_58791# a_37354_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6575 a_2215_36495# a_1591_36501# a_2107_36873# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X6576 a_4001_56377# a_3668_56311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6577 VDD a_12947_71576# a_24302_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6578 a_5805_15279# a_5639_15279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6579 VSS a_15189_39889# a_15221_39631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X658 a_1823_72381# a_2847_66389# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6580 a_48490_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6581 a_3523_13967# a_2283_15797# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6582 a_17711_40183# a_13576_40413# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6583 a_24394_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6584 a_48794_69222# a_12516_7093# a_48398_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6585 VSS a_10975_66407# a_45782_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6586 vcm_commonmode a_16362_60186# a_33430_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6587 a_34434_21540# a_16746_21538# a_34342_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6588 a_2008_28487# a_2223_28617# a_2150_28662# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X6589 vcm_commonmode a_16362_19532# a_33430_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 VDD a_26753_37981# a_26359_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X6590 a_4227_37887# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6591 VDD a_10055_58791# a_12727_58255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u M=3
X6592 a_2923_45743# a_2775_46025# a_2560_45895# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X6593 a_23390_66210# a_16746_66212# a_23298_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6594 a_7523_62581# a_9544_61635# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X6595 a_5803_74397# a_5179_74031# a_5695_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6596 a_4065_70767# a_2686_70223# a_3983_70767# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6597 a_47486_20536# a_16746_20534# a_47394_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6598 a_6377_38133# a_5631_38127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6599 a_22294_21906# a_16362_21540# a_22386_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X66 a_36746_12870# a_10055_58791# a_36350_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X660 VSS a_2223_28617# a_3707_28995# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X6600 result_out[2] a_1644_56053# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6601 VDD a_15439_49525# a_32334_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6602 a_32187_40513# a_12357_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6603 VDD a_12901_66665# a_28318_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6604 a_18278_11866# a_16362_11500# a_18370_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6605 VSS a_2689_65103# a_6905_63151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X6606 VDD a_15253_37692# a_14859_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X6607 VDD a_12899_10927# a_36350_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6608 VSS a_33764_41831# a_33727_42089# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X6609 a_28410_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X661 a_32920_34191# a_32743_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6610 VSS a_12355_65103# a_49798_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6611 a_37446_12504# a_16746_12502# a_37354_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6612 VDD a_12899_11471# a_49402_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6613 VDD a_21856_36513# a_22536_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X6614 a_47486_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6615 a_13848_44135# a_13944_43957# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6616 a_11341_62063# a_11299_62215# a_9643_63125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X6617 a_37354_69222# a_16362_69222# a_37446_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6618 VSS a_12257_56623# a_39758_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6619 a_32334_57174# a_12257_56623# a_32826_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X662 VSS a_6614_21237# a_5085_24759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X6620 a_5437_11791# a_4429_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X6621 a_41462_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6622 a_12901_67279# a_11619_56615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X6623 a_43774_55166# VSS a_43378_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6624 a_23643_29245# a_23051_28023# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6625 a_26706_65206# a_10975_66407# a_26310_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6626 a_6559_27907# a_6773_27805# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X6627 a_7433_65327# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6628 a_9135_22895# a_7187_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=6.565e+11p pd=5.92e+06u as=0p ps=0u w=650000u l=150000u
X6629 VDD a_12901_66959# a_44382_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X663 VDD a_1799_29556# a_4719_33239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6630 a_27236_50095# a_26155_50095# a_26889_50337# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6631 a_32730_12870# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6632 a_7755_68591# a_7707_70741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6633 a_44778_63198# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6634 VSS a_9314_69367# a_10055_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6635 vcm_commonmode a_16362_58178# a_40458_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6636 a_12092_27247# a_11711_27247# a_11902_27497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6637 VSS a_2560_45895# a_2007_45717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6638 VDD a_38115_52263# a_39219_52271# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X6639 vcm_commonmode a_16362_68218# a_23390_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X664 VSS a_35033_38780# a_34725_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u
X6640 a_34639_38825# a_35033_38780# a_34699_38771# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X6641 a_37750_7850# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6642 a_11574_22869# a_12349_25847# a_12355_23983# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6643 a_29718_56170# a_12257_56623# a_29322_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6644 a_2743_36278# a_2473_34293# a_2284_36103# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X6645 a_14008_51727# a_13735_51727# a_13925_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X6646 a_7901_13077# a_8071_13255# a_8029_13353# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6647 a_25321_29673# a_9529_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6648 a_42374_22910# a_10515_23975# a_42866_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6649 a_12565_8545# a_11067_67279# a_12479_8545# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X665 a_38754_22910# a_11067_21583# a_38358_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6650 VSS VDD a_47790_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6651 VDD a_12727_67753# a_48398_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6652 a_45878_64524# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6653 VSS a_12981_62313# a_21686_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6654 a_3417_33231# a_2939_33535# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6655 a_5345_47919# a_5179_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6656 a_18370_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6657 VSS a_12631_28585# a_15661_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X6658 vcm_commonmode a_16362_59182# a_26402_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6659 a_48490_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X666 a_36579_39095# a_35647_39141# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X6660 VDD a_15828_38695# a_15193_41781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6661 a_26218_48981# a_26662_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X6662 a_35742_23914# a_10515_23975# a_35346_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6663 a_30418_57174# a_16746_57176# a_30326_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6664 a_31726_18894# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6665 a_4259_40847# a_4314_40821# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6666 a_35838_56492# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6667 a_28714_9858# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6668 a_48794_22910# a_11067_21583# a_48398_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6669 a_15541_46831# a_5039_42167# a_15457_46831# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X667 a_40366_70226# a_12516_7093# a_40858_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6670 a_8994_63927# a_9643_63125# a_9589_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6671 a_39389_52271# a_39219_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6672 VDD a_5023_13255# a_4995_13103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6673 a_46390_60186# a_12727_58255# a_46882_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6674 a_18278_56170# a_16362_56170# a_18370_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6675 VDD a_11067_66191# a_12662_15939# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6676 VSS a_18627_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X6677 VDD a_10964_25615# a_13335_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X6678 VDD a_5259_39367# a_3759_39991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X6679 a_39854_55488# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X668 VDD a_12727_15529# a_42374_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6680 a_19282_23914# a_12947_23413# a_19774_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6681 a_23298_72234# VDD a_23790_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6682 a_19282_19898# a_16362_19532# a_19374_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6683 a_34738_70226# a_12901_66665# a_34342_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6684 a_49402_12870# a_12877_16911# a_49894_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6685 a_23790_21508# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6686 a_23390_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6687 a_20286_14878# a_16362_14512# a_20378_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6688 a_38450_61190# a_16746_61192# a_38358_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6689 vcm_commonmode a_16362_17524# a_35438_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X669 VDD a_12985_19087# a_23298_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6690 a_11981_20495# a_5535_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6691 VDD a_11887_19087# a_11763_21237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6692 VSS a_12985_16367# a_39758_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6693 vcm_commonmode VSS a_49494_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6694 a_8569_25071# a_8215_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6695 VDD VSS a_16270_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6696 vcm_commonmode VSS a_39454_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6697 a_3210_47741# a_2595_47653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6698 a_11296_14557# a_11082_14557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6699 a_26802_12472# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X67 VDD a_33264_37601# a_33668_38341# VSS sky130_fd_pr__nfet_01v8 ad=8.3123e+14p pd=8.36296e+09u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X670 a_8016_68047# a_7707_70741# a_7761_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X6700 VDD a_27535_30503# a_31551_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6701 a_24302_13874# a_16362_13508# a_24394_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6702 VDD a_12546_22351# a_30326_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6703 a_11759_59575# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X6704 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X6705 a_21686_67214# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6706 a_49494_7484# VDD a_49402_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6707 a_1757_49557# a_1591_49557# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X6708 a_44382_63198# a_12981_62313# a_44874_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6709 VSS a_35079_46831# a_18979_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X671 a_36350_60186# a_12727_58255# a_36842_60508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6710 VSS a_1952_60431# a_1985_53387# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6711 vcm_commonmode a_16362_16520# a_39454_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6712 VSS a_3541_19385# a_3475_19453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6713 a_48398_18894# a_12895_13967# a_48890_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6714 VDD a_25484_37253# a_25388_37253# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X6715 a_22094_51433# a_22164_51157# a_19946_51157# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.3e+11p pd=5.26e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6716 a_43470_14512# a_16746_14510# a_43378_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6717 vcm_commonmode a_16362_11500# a_40458_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6718 VSS a_8367_44343# a_8308_44111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6719 a_23928_28585# a_23303_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X672 VSS a_12516_7093# a_11067_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X6720 a_26402_24552# VDD a_26310_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6721 vcm_commonmode a_16362_21540# a_23390_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6722 a_26815_42405# a_23567_42035# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X6723 a_39454_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6724 VSS config_1_in[14] a_1591_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6725 a_20351_49525# a_20156_49667# a_20661_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X6726 a_12318_71855# a_8575_74853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6727 a_8453_64757# a_6515_62037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=0p ps=0u w=1e+06u l=150000u
X6728 a_16746_62196# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X6729 a_5533_17455# a_5363_17455# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X673 VDD VSS a_25306_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6730 VDD a_38454_43983# a_38999_44527# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6731 a_21782_63520# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6732 VSS a_36607_34191# a_36713_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6733 a_43537_27497# a_41597_29967# a_9503_26151# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X6734 a_31726_59182# a_12727_58255# a_31330_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6735 a_16362_16520# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X6736 a_24302_7850# VSS a_24394_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6737 a_25798_18496# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6738 a_43378_69222# a_12901_66959# a_43870_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6739 a_5879_16367# a_5529_16367# a_5784_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X674 a_49402_20902# a_12985_7663# a_49894_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6740 a_29414_15516# a_16746_15514# a_29322_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6741 vcm_commonmode a_16362_12504# a_26402_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6742 vcm_commonmode a_16362_63198# a_38450_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6743 VDD a_4215_51157# a_26155_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6744 a_30418_10496# a_16746_10494# a_30326_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6745 VDD a_6579_42255# a_6473_40277# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6746 a_2283_32362# a_2235_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X6747 a_4308_45431# a_4458_45565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6748 VDD a_1923_54591# a_2464_54813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6749 a_28714_57174# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X675 a_49402_16886# a_16362_16520# a_49494_16520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6750 a_5905_44905# a_5715_44343# a_5823_44905# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X6751 a_30326_67214# a_16362_67214# a_30418_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6752 VSS a_5085_24759# a_6649_25615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6753 VSS a_11067_47695# a_32730_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6754 VSS a_6559_59663# a_7622_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6755 a_8396_29199# a_8273_42479# a_8206_28879# VSS sky130_fd_pr__nfet_01v8 ad=2.925e+11p pd=2.2e+06u as=0p ps=0u w=650000u l=150000u
X6756 a_20778_69544# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6757 a_44474_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6758 VSS a_15193_42917# a_16707_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X6759 a_20286_59182# a_16362_59182# a_20378_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X676 a_12539_59663# a_11251_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X6760 a_29814_19500# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6761 a_4503_21523# a_4839_21495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X6762 VSS a_3983_12879# a_5457_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X6763 a_1987_33402# a_1867_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6764 a_2592_43023# a_1591_43029# a_2520_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6765 a_8489_74549# a_8271_74953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X6766 a_34391_48682# a_34221_47695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6767 VDD a_3305_38671# a_5631_38127# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6768 VSS a_3295_54421# a_10975_55535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6769 a_40762_17890# a_12899_11471# a_40366_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X677 a_2775_46025# a_2847_45503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X6770 VDD a_5915_30287# a_7561_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6771 a_23734_29941# a_15548_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6772 a_5963_20149# a_8256_20969# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X6773 VDD a_9670_24527# a_12702_25615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X6774 VDD a_11719_28023# a_11968_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6775 a_47790_23914# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6776 VSS a_77002_40202# a_76744_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6777 a_48490_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6778 a_21290_65206# a_12355_65103# a_21782_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6779 a_4458_45565# a_4500_45289# a_4458_45315# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X678 VDD a_26514_47375# a_28108_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.5e+11p ps=5.1e+06u w=1e+06u l=150000u
X6780 a_25204_38567# a_24331_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6781 VDD a_21233_44220# a_20839_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6782 VSS a_9955_20969# a_12082_25077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6783 a_24302_58178# a_16362_58178# a_24394_58178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6784 a_37750_15882# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6785 VDD a_2451_72373# a_10321_74575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6786 vcm_commonmode a_16362_71230# a_20378_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6787 a_20655_34743# a_21049_34717# a_20715_34717# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X6788 VSS a_12727_15529# a_41766_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6789 VSS a_2451_72373# a_2882_73309# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X679 a_41351_38053# a_39468_37479# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X6790 a_19374_64202# a_16746_64204# a_19282_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6791 a_8111_18825# a_8539_18231# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6792 VDD a_11521_58951# a_11759_59575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6793 a_24302_17890# a_12899_10927# a_24794_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6794 VSS a_27891_41495# a_23789_39100# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6795 VDD a_12947_71576# a_32334_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6796 a_21686_20902# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6797 VSS a_12947_23413# a_24698_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6798 VDD a_6515_62037# a_6473_62313# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6799 VSS a_7862_34025# a_26157_31605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X68 a_34342_11866# a_10055_58791# a_34834_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X680 a_6921_72943# a_6453_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X6800 a_9914_68279# a_10379_66389# a_10325_66415# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6801 VDD a_10515_22671# a_31330_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6802 a_2847_42313# a_2401_41941# a_2751_42313# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X6803 a_11345_53359# a_11303_53511# a_10680_54171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6804 a_46786_70226# a_43267_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6805 a_45478_68218# a_16746_68220# a_45386_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6806 VDD a_4571_26677# a_4517_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6807 a_17670_18894# a_12899_10927# a_17274_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6808 a_2789_71855# a_2747_72007# a_2322_72631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6809 VDD a_10973_16609# a_10863_16733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X681 a_27891_41495# a_27999_41495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X6810 vcm_commonmode a_16362_70226# a_24394_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6811 a_10678_14443# a_10995_14333# a_10953_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6812 a_6646_50639# a_3325_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X6813 VDD a_6515_62037# a_8497_54697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6814 a_20378_8488# a_16746_8486# a_20286_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6815 a_33449_30305# a_19626_31751# a_33363_30305# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X6816 a_10717_17209# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6817 VSS a_9307_30663# a_10515_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6818 a_36746_62194# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6819 a_26701_29739# a_27016_29587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X682 a_33819_42359# a_32887_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X6820 a_31726_12870# a_10055_58791# a_31330_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6821 a_43774_63198# a_15439_49525# a_43378_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6822 VSS a_12727_58255# a_40762_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6823 VDD a_35932_38689# a_35033_38780# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X6824 VSS a_11067_67279# a_40762_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6825 a_28318_55166# VSS a_28810_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6826 a_11573_9839# a_2411_18517# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6827 a_19500_42919# a_18627_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6828 VDD a_12727_58255# a_22294_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6829 VSS a_12877_14441# a_18674_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X683 VDD a_7293_42721# a_7183_42845# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X6830 vcm_commonmode a_16362_61190# a_27406_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6831 a_37846_24520# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6832 VSS a_4528_26159# a_6743_23555# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6833 a_31422_18528# a_16746_18526# a_31330_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6834 VDD a_11067_21583# a_41370_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6835 a_10311_20175# a_9955_21807# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+12p pd=1.031e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X6836 a_5455_37039# a_5701_37013# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.646e+11p pd=2.94e+06u as=0p ps=0u w=420000u l=150000u
X6837 a_4060_70223# a_3280_70501# a_3452_70537# VSS sky130_fd_pr__nfet_01v8 ad=1.87e+11p pd=1.93e+06u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X6838 VDD a_2944_63400# a_2882_63517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X6839 a_28714_10862# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X684 a_39362_12870# a_12877_16911# a_39854_12472# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6840 VSS a_32227_48169# a_33957_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X6841 a_2847_19605# a_2672_19631# a_3026_19631# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6842 a_12056_60975# a_10975_60975# a_11709_61217# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X6843 a_3663_39991# a_3305_38671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6844 a_1915_20394# a_2007_20149# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X6845 a_5254_67503# a_4906_67509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6846 a_47790_64202# a_12355_65103# a_47394_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6847 a_22627_51017# a_22181_50645# a_22531_51017# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X6848 a_38358_20902# a_12985_7663# a_38850_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6849 a_5414_39215# a_5490_41365# a_5604_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X685 a_4680_32687# a_4563_32900# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6850 a_45878_72556# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6851 a_38358_16886# a_16362_16520# a_38450_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6852 VDD a_12985_7663# a_45386_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6853 vcm_commonmode a_16362_14512# a_32426_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6854 a_42466_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6855 a_48490_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6856 a_45386_62194# a_16362_62194# a_45478_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6857 a_37750_56170# a_12257_56623# a_37354_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6858 a_28318_72234# VSS a_28410_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6859 a_2012_26159# a_1853_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X686 VSS a_7000_43541# a_11067_67279# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X6860 a_32426_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6861 VDD a_12877_16911# a_35346_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6862 VDD a_8295_47388# a_12899_3311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X6863 vcm_commonmode a_16362_67214# a_44474_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6864 VSS a_3031_47679# a_2965_47753# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6865 VDD a_10515_23975# a_18278_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6866 VSS a_8531_70543# a_33856_50101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6867 VDD a_27236_50095# a_27411_50069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6868 a_4161_73865# a_2971_73493# a_4052_73865# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X6869 VDD a_10055_58791# a_48398_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X687 a_43870_10464# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6870 a_9219_71285# a_9063_71553# a_9364_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X6871 a_18278_64202# a_16362_64202# a_18370_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6872 a_46482_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6873 VSS a_13692_44527# a_13798_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6874 a_22386_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6875 a_7565_31751# a_7295_32259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6876 vcm_commonmode a_16362_59182# a_34434_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6877 VSS a_12546_22351# a_38754_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6878 a_77086_40693# a_75794_40594# vcm_commonmode VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=500000u M=2
X6879 a_12671_37782# a_12641_37684# a_12599_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X688 VSS a_2216_28309# a_5136_34551# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6880 VDD a_12621_44099# a_22352_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6881 vcm_commonmode a_16362_69222# a_17366_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6882 a_7847_39872# a_7373_40847# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X6883 a_6817_37289# a_5631_38127# a_6745_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6884 VDD a_4891_47388# a_27201_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6885 VSS a_19333_48463# a_19991_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X6886 a_33597_50141# a_30928_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6887 a_21382_67214# a_16746_67216# a_21290_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6888 a_48794_9858# a_12985_19087# a_48398_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6889 a_29943_36965# a_27600_36165# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X689 a_26310_71230# a_12901_66665# a_26802_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6890 a_45478_21540# a_16746_21538# a_45386_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6891 a_20286_22910# a_16362_22544# a_20378_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6892 a_36001_31055# a_32823_29397# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6893 VSS a_6775_53877# a_10503_52828# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X6894 a_19374_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6895 VDD a_11067_23759# a_16362_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X6896 a_3137_16367# a_3023_16341# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X6897 VSS a_12139_71829# a_12073_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X6898 a_10667_60735# a_1950_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6899 a_33338_21906# a_16362_21540# a_33430_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X69 a_33484_41605# a_32611_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X690 a_26802_20504# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6900 VDD a_15439_49525# a_43378_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6901 a_35438_13508# a_16746_13506# a_35346_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6902 a_35431_31751# a_29927_29199# a_35665_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X6903 a_14444_29429# a_13239_29575# a_14372_29429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6904 a_23631_50069# a_14831_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6905 a_6725_49557# a_6559_49557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6906 VSS a_10515_22671# a_37750_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6907 a_44382_71230# a_12901_66665# a_44874_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6908 VSS a_4351_67279# a_11883_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6909 a_13051_46831# a_5039_42167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X691 VSS a_12727_67753# a_41766_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X6910 a_35683_50613# a_30928_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=5.72e+06u as=0p ps=0u w=1e+06u l=150000u
X6911 VSS a_8575_74853# a_11661_71855# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6912 a_23507_43177# a_23901_43132# a_23567_43123# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X6913 a_48398_69222# a_16362_69222# a_48490_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6914 VDD a_8827_17215# a_8814_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6915 a_35346_8854# a_12985_19087# a_35838_8456# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6916 VDD a_12981_62313# a_47394_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6917 VSS a_11303_53511# a_11127_53544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6918 a_2952_66139# a_4075_69143# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X6919 VSS a_32971_35281# a_32917_35307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X692 a_26402_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6920 VSS a_29513_42333# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X6921 a_28410_57174# a_16746_57176# a_28318_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6922 a_29718_18894# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6923 a_2702_46070# a_2656_45895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X6924 a_45878_8456# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6925 a_41766_8854# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6926 VSS a_38837_46983# a_38805_47081# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6927 a_30722_13874# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6928 a_1770_14441# a_1591_14191# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X6929 a_31422_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X693 a_1761_49007# a_1591_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X6930 a_76648_40202# a_76744_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6931 VDD a_1586_9991# a_5363_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X6932 a_4404_20719# a_3969_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X6933 a_21782_71552# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6934 a_42466_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6935 VSS a_27560_34337# a_29119_34473# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X6936 a_17766_61512# a_13183_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6937 a_15745_30287# a_13390_29575# a_15443_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6725e+11p ps=2.43e+06u w=650000u l=150000u
X6938 a_17670_8854# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X6939 a_25398_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X694 a_1643_29397# a_1799_29556# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X6940 a_35647_42405# a_34699_42035# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X6941 a_3491_42239# a_3316_42313# a_3670_42301# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6942 a_2203_49929# a_1757_49557# a_2107_49929# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X6943 a_42770_66210# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6944 a_2012_30333# a_1895_30138# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6945 a_30565_30199# a_40691_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6946 a_40366_23914# a_12947_23413# a_40858_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X6947 a_40366_19898# a_16362_19532# a_40458_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6948 VSS a_12985_19087# a_27710_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6949 a_13059_27791# a_11602_25071# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X695 VSS a_38867_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X6950 a_8592_58255# a_7963_58255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X6951 vcm_commonmode a_16362_20536# a_44474_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6952 VSS a_2529_24825# a_2463_24893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6953 VDD a_1761_52815# a_26267_39631# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X6954 a_46482_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6955 a_43378_55166# VSS a_43470_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6956 a_9349_30761# a_9307_30663# a_9161_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6957 VDD a_14831_50095# a_23669_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X6958 a_33830_18496# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6959 a_33734_24918# a_12899_2767# a_33338_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X696 a_29322_64202# a_16362_64202# a_29414_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6960 VSS a_12981_62313# a_32730_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6961 a_8753_31055# a_8215_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6962 VSS a_15660_49257# a_12355_15055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u M=2
X6963 a_29269_44545# a_29391_44031# a_30264_44007# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X6964 a_42466_71230# a_16746_71232# a_42374_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6965 a_3141_59887# a_2785_60151# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6966 a_29414_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6967 a_22690_69222# a_12516_7093# a_22294_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6968 VDD a_9529_28335# a_25462_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.8668e+12p ps=1.774e+07u w=1e+06u l=150000u M=4
X6969 vcm_commonmode a_16362_12504# a_34434_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X697 VDD a_12981_62313# a_29322_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X6970 a_46882_17492# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6971 a_43378_14878# a_12877_14441# a_43870_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6972 a_46786_23914# a_10515_23975# a_46390_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6973 a_3040_68425# a_2125_68053# a_2693_68021# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X6974 a_44382_18894# a_16362_18528# a_44474_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6975 a_12671_37455# a_12417_37782# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X6976 VSS a_2843_71829# a_7289_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=2
X6977 a_8539_18231# a_5535_18012# a_8937_18319# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X6978 vcm_commonmode a_16362_22544# a_17366_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6979 VDD a_17475_51157# a_17462_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X698 VDD a_9624_65301# a_10147_65984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X6980 a_26310_24918# VSS a_26802_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X6981 a_7337_45565# a_7293_45173# a_7171_45577# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6982 a_33802_47375# a_22015_28111# a_33730_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X6983 a_21382_20536# a_16746_20534# a_21290_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6984 VDD a_12907_56399# a_16362_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X6985 a_30818_22512# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6986 VDD a_31280_40517# a_31184_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X6987 a_8491_27023# a_12815_4399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X6988 a_22727_29199# a_18053_28879# a_22631_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.08e+11p pd=1.94e+06u as=0p ps=0u w=650000u l=150000u
X6989 a_20378_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X699 vcm_commonmode VSS a_39454_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6990 a_36746_15882# a_12877_14441# a_36350_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6991 VDD a_20635_29415# a_43537_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6992 a_19678_67214# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6993 a_4514_58387# a_4831_58497# a_4789_58621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X6994 a_46482_70226# a_16746_70228# a_46390_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6995 a_7407_18038# a_7377_18012# a_7335_18038# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6996 a_9963_29967# a_8739_28879# a_10045_30287# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u
X6997 a_11477_69679# a_11433_69921# a_11311_69679# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X6998 a_2840_53511# a_6743_54447# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X6999 VSS a_12355_65103# a_23694_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_8364_47919# a_6863_42692# a_8143_48246# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X70 a_19678_64202# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X700 VDD a_2325_45173# a_2215_45199# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7000 a_49798_56170# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7001 a_16928_44007# a_15959_44031# a_16891_44265# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X7002 VDD a_12899_11471# a_23298_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7003 a_20778_14480# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7004 a_47394_13874# a_12727_15529# a_47886_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7005 VDD a_12947_8725# a_30326_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7006 a_21382_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7007 a_10003_55862# a_9821_55862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7008 VDD a_6516_53511# a_6467_53359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7009 VDD a_22989_48437# a_23850_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 VDD a_19439_32143# a_4443_46607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X7010 VSS a_4891_47388# a_22951_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7011 a_41862_68540# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7012 a_36442_62194# a_16746_62196# a_36350_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7013 vcm_commonmode a_16362_8488# a_43470_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7014 a_7896_18695# a_8111_18825# a_8038_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X7015 a_7634_57961# a_6515_62037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7016 a_37846_58500# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7017 a_31330_14878# a_16362_14512# a_31422_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7018 a_8361_15529# a_7959_15279# a_8197_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X7019 VSS a_16228_28335# a_17459_31145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X702 VDD a_38171_43983# a_38277_43983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7020 a_5345_47919# a_5179_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7021 a_19374_72234# VDD a_19282_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7022 VSS a_10055_58791# a_37750_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7023 a_49494_61190# a_16746_61192# a_49402_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7024 vcm_commonmode a_16362_17524# a_46482_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7025 VSS a_12947_56817# a_26706_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7026 vcm_commonmode a_16362_8488# a_19374_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7027 VDD a_12727_13353# a_27314_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7028 a_24794_13476# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7029 a_21290_10862# a_12985_16367# a_21782_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X703 VDD a_5039_42167# a_11619_56615# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u M=4
X7030 a_53260_40156# a_7841_12167# a_53906_40254# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=0p ps=0u w=800000u l=150000u
X7031 VDD a_14524_48437# a_10975_66407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X7032 a_42374_64202# a_11067_13095# a_42866_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7033 a_29414_8488# a_16746_8486# a_29322_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7034 a_2589_62839# a_2605_60975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7035 a_28410_10496# a_16746_10494# a_28318_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7036 a_20649_36391# a_20623_36595# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7037 a_2325_10081# a_2107_9839# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7038 a_12875_31751# a_7695_31573# a_13049_31627# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7039 VSS a_14049_42869# a_13983_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X704 a_21290_9858# a_16362_9492# a_21382_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7040 a_3870_60563# a_4148_60547# a_4104_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7041 VSS a_10984_58487# a_6417_62215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7042 a_25104_51183# a_8123_56399# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7043 VDD a_22843_29415# a_36613_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7044 a_18770_69544# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7045 a_8296_56873# a_7773_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.35e+11p pd=2.47e+06u as=0p ps=0u w=1e+06u l=150000u
X7046 VDD a_12727_67753# a_22294_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7047 a_28670_30663# a_28513_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X7048 a_32826_63520# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7049 VSS a_3572_56311# a_2419_55687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X705 VDD a_12546_22351# a_20286_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7050 a_27406_16520# a_16746_16518# a_27314_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7051 a_1644_56053# a_1591_54447# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7052 a_5037_32687# a_4993_32929# a_4871_32687# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X7053 VDD a_1586_45431# a_7387_48469# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7054 a_4241_18543# a_4075_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7055 a_22690_22910# a_11067_21583# a_22294_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7056 a_19282_65206# a_12355_65103# a_19774_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7057 a_24413_39087# a_23987_39126# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7058 a_26706_58178# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7059 a_39454_69222# a_16746_69224# a_39362_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X706 a_45782_8854# a_12947_8725# a_45386_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7060 a_20286_60186# a_12727_58255# a_20778_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7061 vcm_commonmode a_16362_66210# a_36442_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7062 a_47790_72234# VDD a_47394_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7063 a_40458_64202# a_16746_64204# a_40366_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7064 VSS a_18126_28023# a_18084_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7065 a_16746_59184# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X7066 a_38358_24918# VSS a_38450_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7067 a_42466_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7068 VDD a_11659_66567# a_11711_67325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7069 a_7749_49929# a_6559_49557# a_7640_49929# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X707 a_10101_51183# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7070 a_8117_12879# a_1929_12131# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7071 a_19678_20902# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7072 a_2596_16911# a_1591_16917# a_2520_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.66e+10p ps=1.3e+06u w=420000u l=150000u
X7073 VSS a_5085_24759# a_5087_23145# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7074 VSS a_12981_59343# a_34738_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7075 a_8079_43732# a_8171_43541# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7076 VSS a_20359_27791# a_20881_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u M=2
X7077 a_11281_30511# a_9367_29397# a_11372_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7078 VSS a_12901_66665# a_17670_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7079 a_13146_51005# a_2419_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X708 a_13983_42895# a_13835_43177# a_13620_43047# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7080 VDD a_1586_51335# a_11711_50645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7081 a_31330_59182# a_16362_59182# a_31422_59182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7082 a_11424_23983# a_7841_22895# a_11121_23957# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X7083 a_45782_24918# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7084 a_2011_34837# a_4903_29975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7085 a_6155_15279# a_5805_15279# a_6060_15279# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X7086 VSS a_6372_38279# a_8656_34639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7087 VSS a_12727_58255# a_38754_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7088 a_28318_9858# a_12546_22351# a_28810_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7089 a_34434_55166# VDD a_34342_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X709 VDD a_8485_71855# a_9782_71311# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X7090 a_35742_16886# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7091 VSS a_11067_67279# a_38754_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7092 a_4852_23413# a_3972_25615# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X7093 VSS a_3357_67257# a_3291_67325# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7094 a_5245_61225# a_3295_62083# a_5173_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7095 a_28980_41831# a_28011_41855# a_28943_42089# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7096 a_35185_43781# a_35493_43421# a_30412_42589# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7097 a_17366_65206# a_16746_65208# a_17274_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7098 a_12484_25935# a_12349_25847# a_12394_25615# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X7099 a_18811_42405# a_16928_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X71 a_2319_54684# a_2163_54589# a_2464_54813# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X710 VSS a_2375_76372# a_1823_77821# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7100 a_49402_71230# a_16362_71230# a_49494_71230# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7101 a_48794_15882# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7102 a_22294_18894# a_12895_13967# a_22786_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7103 VSS VSS a_22690_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7104 a_4699_18909# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7105 a_19374_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7106 VDD a_11067_23759# a_16362_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X7107 vcm_commonmode a_16362_71230# a_31422_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7108 a_22536_35303# a_21663_35327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7109 VDD a_5749_60039# a_5515_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X711 a_34342_63198# a_12981_62313# a_34834_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7110 VDD a_19531_49007# a_19715_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7111 VDD a_12947_71576# a_43378_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7112 a_28115_40183# a_27183_40229# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X7113 VDD a_12355_15055# a_39362_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7114 VDD a_1586_69367# a_7755_74581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7115 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7116 a_43470_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7117 a_11311_69679# a_10865_69679# a_11215_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7118 VSS a_26319_38517# a_24892_38237# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7119 VDD config_1_in[3] a_1591_13103# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X712 a_22260_39655# a_20713_40193# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X7120 VSS a_16744_41605# a_16707_41271# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X7121 a_28239_52105# a_27793_51733# a_28143_52105# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X7122 a_26402_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7123 a_28714_18894# a_12899_10927# a_28318_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7124 VSS a_12727_13353# a_25702_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7125 a_28618_32143# a_14646_29423# a_27890_32459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X7126 a_9028_63695# a_8994_63927# a_8773_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X7127 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7128 a_16707_34473# a_15775_34239# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7129 VSS a_24800_43041# a_34823_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X713 VSS a_37557_32463# a_38013_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X7130 VDD a_12901_66665# a_47394_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7131 a_37354_11866# a_16362_11500# a_37446_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7132 a_6269_43567# a_5791_43541# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7133 a_34943_51335# a_35495_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7134 a_5426_39465# a_3949_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7135 a_4227_37887# a_4052_37961# a_4406_37949# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7136 a_30326_68218# a_12727_67753# a_30818_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7137 a_9649_58255# a_7210_55081# a_9215_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7138 a_41766_66210# a_12983_63151# a_41370_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7139 VDD a_2589_55535# a_2882_56989# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X714 VSS a_12901_58799# a_44778_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7140 vcm_commonmode a_16362_62194# a_25398_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7141 a_26310_58178# a_10515_22671# a_26802_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7142 VSS a_9370_69831# a_9319_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7143 VDD a_2244_22583# a_2021_22325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7144 VSS a_12877_14441# a_29718_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7145 a_26706_11866# a_26748_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7146 VSS a_33798_31145# a_33593_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7147 VDD a_1586_40455# a_6559_49557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7148 a_39454_22544# a_16746_22542# a_39362_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7149 a_22808_27497# a_19889_27497# a_12869_2741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X715 a_41766_56170# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7150 a_28789_50613# a_29055_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7151 a_30557_49783# a_26397_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7152 VSS config_2_in[13] a_1591_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7153 VSS a_3327_9308# a_7803_11703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7154 a_38754_64202# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7155 a_33261_51433# a_33313_51157# a_10687_52553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u M=2
X7156 a_45782_65206# a_10975_66407# a_45386_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7157 a_8497_72105# a_2451_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7158 a_36350_21906# a_11067_21583# a_36842_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7159 a_36350_17890# a_16362_17524# a_36442_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X716 VDD a_19889_27497# a_22026_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u M=4
X7160 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7161 a_40458_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7162 a_26631_35877# a_25484_37253# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X7163 a_43378_63198# a_16362_63198# a_43470_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7164 a_2012_19631# a_1867_20175# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X7165 a_11413_12015# a_10935_11989# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7166 VDD a_18979_30287# a_43539_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X7167 a_33430_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7168 a_35742_57174# a_10515_22671# a_35346_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7169 VDD a_2847_66389# a_2834_66781# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X717 a_38358_18894# a_12895_13967# a_38850_18496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7170 a_37750_8854# a_12947_8725# a_37354_8854# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7171 VDD a_3325_69135# a_4075_69143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7172 a_11082_14557# a_10995_14333# a_10678_14443# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=420000u l=150000u
X7173 vcm_commonmode a_16362_68218# a_42466_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7174 a_18674_67214# a_12727_67753# a_18278_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7175 VSS a_10659_9813# a_9484_11989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7176 a_31873_37253# a_32181_36893# a_31847_36893# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7177 a_48794_56170# a_12257_56623# a_48398_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7178 VDD a_35932_37601# a_35033_37692# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X7179 VDD a_12877_16911# a_46390_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X718 a_27314_12870# a_16362_12504# a_27406_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7180 VDD a_5064_45743# a_5239_45717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7181 VDD a_13390_29575# a_15851_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.025e+12p ps=6.05e+06u w=1e+06u l=150000u
X7182 VDD a_12907_56399# a_16362_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X7183 VSS a_14983_51157# a_14941_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X7184 VDD a_11667_63303# a_11619_63151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7185 a_20378_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7186 VDD a_10515_23975# a_29322_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7187 a_4357_69929# a_2952_66139# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7188 VDD a_15607_46805# a_35228_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7189 a_4621_36611# a_4495_35925# a_4525_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X719 a_6835_23983# a_5531_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7190 a_20682_70226# a_16955_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7191 vcm_commonmode a_16362_59182# a_45478_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7192 a_41141_32463# a_35815_31751# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X7193 VDD a_7289_70767# a_7387_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X7194 VDD a_12877_14441# a_19282_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7195 VSS a_37527_29397# a_16863_29415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=2
X7196 vcm_commonmode a_16362_69222# a_28410_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7197 a_34342_24918# a_12899_3311# a_34834_24520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7198 VSS a_3983_16617# a_4630_15823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X7199 a_32426_67214# a_16746_67216# a_32334_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X72 VSS a_14926_31849# a_17554_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.46e+11p ps=5.58e+06u w=650000u l=150000u M=2
X720 a_33430_14512# a_16746_14510# a_33338_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7200 a_40581_31599# a_40233_31605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X7201 VSS a_16510_8760# a_16746_8486# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X7202 VDD a_4427_30511# a_6099_23983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7203 a_37846_66532# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7204 a_31330_22910# a_16362_22544# a_31422_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7205 VDD a_12355_65103# a_41370_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7206 a_39454_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7207 a_8493_27791# a_3607_34639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7208 a_37354_56170# a_16362_56170# a_37446_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7209 a_34834_7452# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X721 a_42866_16488# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7210 a_2371_28335# a_2223_28617# a_2008_28487# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7211 a_23694_61190# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7212 a_22386_59182# a_16746_59184# a_22294_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7213 a_8076_10383# a_7862_10383# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7214 vcm_commonmode a_16362_58178# a_49494_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7215 a_30722_62194# a_12981_62313# a_30326_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7216 a_25388_37253# a_24515_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7217 a_2560_45895# a_2775_46025# a_2702_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X7218 VDD VDD a_44382_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7219 VSS VDD a_40762_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X722 a_16746_70228# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7220 a_42374_72234# VDD a_42866_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7221 VDD a_2163_63293# a_2124_63419# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7222 a_38358_62194# a_12355_15055# a_38850_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7223 a_5885_39759# a_3305_38671# a_5731_40079# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X7224 a_6369_10927# a_5179_10927# a_6260_10927# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X7225 a_42866_60508# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7226 VSS VDD a_16666_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u M=2
X7227 a_32334_7850# VDD a_32826_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7228 VSS a_4215_51157# a_24683_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7229 a_27710_60186# a_23395_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X723 VDD config_2_in[9] a_1591_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7230 a_26402_58178# a_16746_58180# a_26310_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7231 vcm_commonmode VSS a_23390_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7232 a_27710_19898# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7233 a_43445_28335# a_18703_29199# a_43227_28309# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7234 a_21686_9858# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7235 a_26706_7850# VDD a_26310_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7236 VDD VSS a_35346_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7237 a_4513_55357# a_4035_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7238 a_23850_48463# a_23631_50069# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7239 a_10035_60431# a_1950_59887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X724 a_11067_66191# a_5039_42167# a_13413_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X7240 a_2847_71615# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7241 VDD a_10975_66407# a_18278_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7242 a_39758_71230# a_12947_71576# a_39362_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7243 a_28810_22512# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7244 a_32826_71552# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7245 a_40762_67214# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7246 a_18370_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7247 a_2055_61225# a_1770_14441# a_1959_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7248 a_2107_9839# a_1757_9839# a_2012_9839# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X7249 a_32334_61190# a_16362_61190# a_32426_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X725 VSS a_12901_66959# a_27710_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7250 a_35742_10862# a_12546_22351# a_35346_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7251 VSS a_2008_28487# a_1683_27399# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7252 vcm_commonmode a_16362_21540# a_42466_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7253 a_18770_14480# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7254 a_18674_20902# a_11067_67279# a_18278_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7255 a_26311_31849# a_25263_29981# a_26239_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7256 a_19684_41605# a_18811_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X7257 VDD a_3987_19623# a_4043_44343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7258 VDD a_10055_58791# a_22294_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7259 a_6185_23145# a_4427_25071# a_6089_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X726 VDD a_38837_46983# a_38805_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X7260 a_40458_72234# VDD a_40366_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7261 a_18278_7850# VSS a_18370_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7262 a_1761_9295# a_1591_9295# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7263 a_29322_14878# a_16362_14512# a_29414_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7264 a_2926_33231# a_1849_33237# a_2764_33609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7265 a_41370_15882# a_12727_13353# a_41862_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7266 a_44874_18496# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7267 a_44778_24918# VSS a_44382_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7268 VSS a_10975_66407# a_30722_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7269 VDD a_25269_27791# a_27250_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u M=2
X727 VDD a_10607_58799# a_7773_63927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7270 a_48490_15516# a_16746_15514# a_48398_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7271 vcm_commonmode a_16362_12504# a_45478_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7272 VDD a_28757_27247# a_30663_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X7273 a_19282_10862# a_12985_16367# a_19774_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7274 a_21479_42405# a_19596_42919# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X7275 a_34738_58178# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7276 a_42466_7484# VDD a_42374_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7277 vcm_commonmode a_16362_22544# a_28410_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7278 a_34738_16886# a_12727_13353# a_34342_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7279 a_32426_20536# a_16746_20534# a_32334_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X728 a_16362_24552# VDD a_16270_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7280 a_17670_68218# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7281 a_1761_30511# a_1591_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X7282 a_47790_57174# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7283 VSS a_27411_50069# a_27869_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X7284 a_11763_62581# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7285 VDD a_12899_10927# a_21290_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7286 a_30633_48829# a_17682_50095# a_30561_48829# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7287 a_18370_7484# VDD a_18278_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7288 a_29175_28335# a_28902_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7289 VSS a_39176_44527# a_39282_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X729 a_31726_67214# a_12727_67753# a_31330_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7290 a_30127_38053# a_29361_38017# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X7291 a_22386_12504# a_16746_12502# a_22294_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7292 a_34434_63198# a_16746_63200# a_34342_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7293 vcm_commonmode a_16362_11500# a_49494_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7294 a_35647_41317# a_33764_41831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X7295 vcm_commonmode a_16362_9492# a_23390_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7296 a_35838_59504# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7297 a_33593_31287# a_33798_31145# a_33756_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7298 a_32426_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7299 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X73 a_31184_36165# a_31280_36165# VDD VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u M=2
X730 a_23258_50639# a_22181_50645# a_23096_51017# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7300 a_48890_19500# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7301 a_2672_30345# a_1591_29973# a_2325_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7302 a_47486_62194# a_16746_62196# a_47394_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7303 a_22294_69222# a_16362_69222# a_22386_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7304 VSS a_12257_56623# a_24698_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7305 a_18278_16886# a_12899_11471# a_18770_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7306 a_38850_9460# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7307 a_17712_7638# a_18979_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X7308 a_1643_57685# a_1846_57963# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7309 a_2107_44655# a_1757_44655# a_2012_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X731 a_6155_15279# a_5639_15279# a_6060_15279# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X7310 a_3202_68047# a_2125_68053# a_3040_68425# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7311 a_40366_65206# a_12355_65103# a_40858_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7312 a_26402_11500# a_16746_11498# a_26310_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7313 VDD a_12985_19087# a_48398_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7314 a_33015_40513# a_12357_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7315 a_2479_50899# a_2419_48783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X7316 VDD a_12895_13967# a_25306_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7317 a_7801_46653# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7318 a_2319_73180# a_2163_73085# a_2464_73309# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X7319 a_38450_64202# a_16746_64204# a_38358_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X732 a_46482_13508# a_16746_13506# a_46390_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7320 VDD a_5208_70063# a_5295_69135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X7321 VDD a_1954_61677# a_3983_59887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7322 VSS a_28639_49551# a_28648_50101# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7323 a_40762_20902# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7324 VSS a_12947_23413# a_43774_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7325 VSS a_2411_18517# a_11173_12015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7326 a_2752_62723# a_2605_60975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7327 VSS a_12381_43957# a_12800_43983# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7328 a_12727_15529# a_12355_15055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X7329 a_43378_56170# a_12947_56817# a_43870_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X733 vcm_commonmode a_16362_10496# a_43470_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7330 a_29814_69544# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7331 a_26310_66210# a_10975_66407# a_26802_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7332 a_30818_64524# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7333 a_2672_9839# a_1757_9839# a_2325_10081# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X7334 VSS a_4571_26677# a_7755_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7335 VSS a_12727_13353# a_33734_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7336 VDD a_39331_34191# a_11067_23759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X7337 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7338 VDD a_1586_51335# a_1591_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7339 a_29322_59182# a_16362_59182# a_29414_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X734 a_10391_49855# a_10216_49929# a_10570_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7340 a_31117_29199# a_30788_28487# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7341 a_26020_30199# a_7939_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7342 a_4775_32687# a_4259_32687# a_4680_32687# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X7343 a_20682_23914# a_10515_23975# a_20286_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7344 VSS a_9011_74879# a_6224_73095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X7345 a_2347_28918# a_2011_34837# a_2347_29245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7346 a_20778_56492# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7347 a_46390_9858# a_16362_9492# a_46482_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7348 a_38754_72234# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7349 a_47394_55166# VSS a_47886_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X735 result_out[1] a_1644_54965# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X7350 VSS a_12516_7093# a_42770_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7351 a_15959_42943# a_15193_42917# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X7352 a_34342_58178# a_10515_22671# a_34834_58500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7353 a_36324_34191# a_36147_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7354 a_12165_65327# a_10975_65327# a_12056_65327# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X7355 a_21737_49249# a_21519_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X7356 a_31330_60186# a_12727_58255# a_31822_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7357 a_34738_11866# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7358 VSS a_5601_11471# a_5483_11140# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7359 a_40458_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X736 vcm_commonmode a_16362_20536# a_26402_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7360 a_36357_47375# a_12907_27023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7361 a_7901_57961# a_7580_61751# a_7467_57863# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X7362 a_37307_29423# a_37527_29397# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7363 a_19780_39429# a_18811_39141# a_19684_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7364 VDD a_23901_43132# a_23507_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7365 a_17670_21906# a_17712_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7366 a_35487_49871# a_35676_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7367 vcm_commonmode a_16362_71230# a_29414_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7368 VSS a_15548_30761# a_21879_30663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7369 a_47790_10862# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X737 a_29414_23548# a_16746_23546# a_29322_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7370 VDD a_36116_44765# a_35217_44509# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X7371 a_31004_44869# a_30035_44581# a_30967_44535# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7372 a_8679_36495# a_5363_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7373 a_38628_47349# a_38805_47081# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7374 a_24794_55488# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7375 a_10531_31055# a_10280_31171# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7376 VSS a_12981_59343# a_45782_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7377 a_1846_57963# a_2163_57853# a_2121_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X7378 a_1915_35015# a_3983_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X7379 VDD a_4429_14191# a_5731_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X738 VDD a_36600_49159# a_36551_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X7380 a_4499_20719# a_3983_20719# a_4404_20719# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X7381 a_23390_61190# a_16746_61192# a_23298_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7382 vcm_commonmode a_16362_17524# a_20378_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7383 VDD a_12899_2767# a_33338_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7384 a_6683_37815# a_6377_38133# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7385 VDD a_42188_43677# a_42224_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7386 a_27710_13874# a_12877_16911# a_27314_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7387 VSS a_12985_16367# a_24698_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7388 VDD a_2847_38975# a_2834_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7389 a_8583_33551# a_3339_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X739 VDD a_8566_39215# a_9821_46831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X7390 VSS a_22989_48437# a_23019_48463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X7391 a_47394_72234# VSS a_47486_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7392 VSS a_12727_58255# a_49798_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7393 a_45478_55166# VDD a_45386_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7394 VSS a_11067_67279# a_49798_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7395 a_46786_16886# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7396 a_39758_7850# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7397 a_3417_31599# a_2939_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7398 VSS a_1923_54591# a_4273_55357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7399 vcm_commonmode a_16362_16520# a_24394_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X74 vcm_commonmode a_16362_23548# a_43470_23548# VSS sky130_fd_pr__nfet_01v8 ad=1.55518e+14p pd=1.74372e+09u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X740 VSS a_19096_36513# a_18197_36604# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X7400 a_34834_20504# a_33864_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7401 VDD a_10515_23975# a_37354_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7402 VDD VDD a_41370_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7403 a_34434_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7404 a_33338_18894# a_12895_13967# a_33830_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7405 a_8489_74549# a_8271_74953# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7406 a_37354_64202# a_16362_64202# a_37446_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7407 VDD a_17867_32117# a_17798_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7408 a_31422_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7409 a_41462_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X741 a_21686_59182# a_12727_58255# a_21290_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7410 a_37520_49783# a_35676_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7411 VSS a_6835_46823# a_26259_47491# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7412 VDD a_11763_62581# a_11395_62037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7413 a_11893_65871# a_11619_63151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7414 a_5913_74273# a_5695_74031# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X7415 a_17199_49007# a_16753_49007# a_17103_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X7416 a_24394_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7417 a_26706_60186# a_12981_59343# a_26310_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7418 a_31648_43781# a_30679_43493# a_31611_43447# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7419 a_26706_19898# a_12895_13967# a_26310_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X742 a_7000_43541# a_7847_40847# a_8375_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7420 a_1959_61225# a_1768_16367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7421 a_1644_66933# a_1823_66941# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X7422 a_38358_70226# a_12516_7093# a_38850_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7423 a_6841_14013# a_4812_13879# a_6769_14013# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7424 VDD a_20635_29415# a_39305_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X7425 a_38450_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7426 a_35346_12870# a_16362_12504# a_35438_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7427 VSS a_1915_35015# a_4437_34639# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7428 VSS a_15557_52245# a_15315_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7429 VSS a_12901_66959# a_35742_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X743 VSS a_10515_22671# a_48794_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7430 vcm_commonmode a_16362_63198# a_23390_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7431 VSS a_10055_58791# a_12257_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7432 a_48398_11866# a_16362_11500# a_48490_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7433 a_9765_32143# a_9318_32509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7434 VSS config_1_in[3] a_1591_13103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7435 a_40613_41605# a_40921_41245# a_13909_41923# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7436 a_5592_56989# a_5378_56989# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7437 a_37446_23548# a_16746_23546# a_37354_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7438 a_6883_37019# a_3607_34639# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7439 a_12621_36091# a_35647_35877# a_36579_35831# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X744 a_45782_55166# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7440 a_7969_58799# a_3668_56311# a_7871_59049# VSS sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X7441 VSS a_24331_39679# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7442 a_18811_41317# a_18045_41281# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X7443 a_18370_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7444 a_28251_51727# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7445 VSS a_12727_67753# a_39758_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7446 a_36746_65206# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7447 VDD a_5269_43809# a_5159_43933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7448 a_25263_29981# a_25368_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X7449 a_25398_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X745 a_23303_31171# a_15548_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X7450 a_41766_9858# a_12985_19087# a_41370_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7451 a_14287_27247# a_11866_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.8025e+11p pd=3.77e+06u as=0p ps=0u w=650000u l=150000u
X7452 VDD a_12889_40977# a_12831_41085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7453 a_6743_29673# a_5449_25071# a_6825_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X7454 VSS a_7707_70741# a_7289_70767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X7455 VDD a_12546_22351# a_18278_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7456 vcm_commonmode a_16362_64202# a_27406_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7457 a_6792_43719# a_6269_43567# a_6934_43894# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X7458 a_33734_58178# a_12901_58799# a_33338_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7459 a_10717_17209# a_2143_15271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X746 a_37354_8854# a_16362_8488# a_37446_8488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7460 a_11480_10205# a_11266_10205# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7461 a_17670_9858# a_12985_19087# a_17274_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7462 a_9955_20969# a_7187_23439# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7463 a_32730_23914# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7464 a_29322_22910# a_16362_22544# a_29414_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7465 a_11377_30761# a_10595_30511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7466 a_32227_48169# a_31753_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.1125e+11p pd=1.95e+06u as=0p ps=0u w=650000u l=150000u
X7467 a_36842_61512# a_36717_47375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7468 a_44474_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7469 a_46786_57174# a_10515_22671# a_46390_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X747 a_10338_19631# a_10394_19605# a_8933_22583# VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X7470 VDD a_12907_27023# a_30745_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7471 a_41370_66210# a_16362_66210# a_41462_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7472 VSS a_2315_24540# a_2981_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X7473 a_30835_38695# a_30943_38695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7474 a_12727_67753# a_11067_67279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X7475 a_5607_44343# a_5715_44343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7476 vcm_commonmode a_16362_56170# a_17366_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7477 a_2203_30345# a_1757_29973# a_2107_30345# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X7478 a_29718_67214# a_12727_67753# a_29322_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7479 a_5805_15279# a_5639_15279# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X748 a_28714_65206# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7480 a_5735_37699# a_5631_38127# a_5639_37699# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7481 a_22690_15882# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7482 VDD a_2417_33205# a_2307_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7483 VDD a_35036_34191# a_35142_34191# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7484 a_11323_70045# a_8575_74853# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7485 a_19678_59182# a_12727_58255# a_19282_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7486 a_25517_37455# a_25091_37782# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7487 a_48490_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7488 a_31726_70226# a_31768_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7489 a_30418_68218# a_16746_68220# a_30326_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X749 a_11866_27791# a_9179_22351# a_11794_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.025e+12p pd=6.05e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7490 VSS a_27239_36341# a_13576_37149# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7491 VSS a_23628_35823# a_23734_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7492 a_6641_27907# a_4427_25071# a_6559_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7493 a_6559_27907# a_4427_25071# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7494 a_35838_67536# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7495 a_2199_33609# a_1683_33237# a_2104_33597# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X7496 VSS a_10949_72719# a_10969_71631# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7497 a_45386_24918# VSS a_45878_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7498 a_35346_57174# a_16362_57174# a_35438_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7499 a_7761_37583# a_3305_38671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X75 a_19678_22910# a_11067_21583# a_19282_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X750 a_26353_34215# a_26661_34428# a_13484_39325# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X7500 a_12703_38517# a_12801_38517# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7501 a_21686_62194# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7502 VSS a_7619_62581# a_7553_62927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X7503 a_24800_35425# a_24331_34239# a_25204_34215# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7504 a_18278_67214# a_16362_67214# a_18370_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7505 VDD a_12981_59343# a_17274_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7506 a_7828_31849# a_7281_29423# a_7571_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X7507 a_33430_9492# a_16746_9490# a_33338_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7508 a_39673_28111# a_39727_27765# a_39685_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7509 a_48398_56170# a_16362_56170# a_48490_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X751 a_19374_15516# a_16746_15514# a_19282_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7510 a_11964_18543# a_11049_18543# a_11617_18785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7511 VDD a_12947_8725# a_24302_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7512 VSS a_10515_23975# a_35742_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7513 VSS a_12985_19087# a_20682_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7514 VDD a_12899_11471# a_42374_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7515 VSS a_15775_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7516 a_6993_20969# a_4792_20443# a_6921_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7517 a_5087_24643# a_4333_22895# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7518 VDD a_35932_38689# a_36520_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7519 a_22786_24520# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X752 VSS a_11067_23759# a_16362_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X7520 a_29269_40741# a_29943_41317# a_30875_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7521 a_49402_23914# a_12947_23413# a_49894_23516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7522 a_49402_19898# a_16362_19532# a_49494_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7523 VSS a_28446_31375# a_30008_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7524 a_7695_31573# a_7390_32693# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X7525 a_12815_16519# a_12580_15939# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7526 a_38450_72234# VDD a_38358_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7527 a_2307_52637# a_1923_54591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7528 a_25398_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7529 VDD a_9219_11471# a_10103_11079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X753 a_28785_47919# a_6831_63303# a_28524_47919# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X7530 a_23192_27791# a_22567_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=150000u
X7531 a_39362_15882# a_12727_13353# a_39854_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7532 VSS a_11067_21583# a_39758_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7533 a_43870_13476# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7534 a_6459_30511# a_5915_30511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X7535 a_40366_10862# a_12985_16367# a_40858_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7536 VSS a_10975_66407# a_28714_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7537 a_1644_58229# a_1591_56623# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7538 a_9379_15039# a_9204_15113# a_9558_15101# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X7539 a_5909_51433# a_3325_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X754 a_6841_40125# a_3305_38671# a_6769_40125# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7540 VDD VSS a_46390_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7541 VDD a_12879_38517# a_12703_38517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7542 a_23298_20902# a_12985_7663# a_23790_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7543 a_26802_23516# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7544 a_26402_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7545 VSS a_17863_44211# a_17803_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X7546 a_30967_44535# a_30035_44581# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7547 a_30818_72556# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7548 a_23298_16886# a_16362_16520# a_23390_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7549 VDD a_12985_7663# a_30326_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X755 a_3173_66169# a_2840_66103# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7550 a_19878_49683# a_20156_49667# a_20112_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7551 VDD a_12901_58799# a_33338_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7552 VDD a_10975_66407# a_29322_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7553 a_33734_11866# a_12985_16367# a_33338_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7554 a_30326_62194# a_16362_62194# a_30418_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7555 a_18848_27765# a_18307_27791# a_18977_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X7556 VDD a_24683_48463# a_23830_49525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7557 VDD a_4037_58773# a_3618_58487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7558 a_29414_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7559 a_42466_17524# a_16746_17522# a_42374_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X756 a_10501_65871# a_10147_65984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7560 VDD a_6097_16609# a_5987_16733# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7561 a_22690_56170# a_12257_56623# a_22294_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7562 VSS a_3307_18259# a_2411_18517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X7563 VDD a_12877_16911# a_20286_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7564 a_46786_10862# a_12546_22351# a_46390_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7565 VDD a_9869_67745# a_9759_67869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7566 VDD a_10515_22671# a_19282_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7567 a_34342_66210# a_10975_66407# a_34834_66532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7568 a_29814_14480# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7569 a_29718_20902# a_11067_67279# a_29322_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X757 a_20378_10496# a_16746_10494# a_20286_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7570 VDD a_8935_27791# a_11866_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7571 a_41766_59182# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7572 a_27314_15882# a_16362_15516# a_27406_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7573 a_6927_65871# a_3143_66972# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7574 a_31422_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7575 a_3229_27791# a_2315_24540# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7576 a_9865_14441# a_7841_12167# a_9865_14191# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7577 a_46482_16520# a_16746_16518# a_46390_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7578 vcm_commonmode a_16362_13508# a_43470_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7579 a_19678_12870# a_10055_58791# a_19282_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X758 a_26310_18894# a_16362_18528# a_26402_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7580 VSS a_34391_48682# a_31768_55394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7581 a_17274_11866# a_10055_58791# a_17766_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7582 a_2325_45173# a_2107_45577# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7583 VDD a_5331_18517# a_5318_18909# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7584 vcm_commonmode a_16362_23548# a_26402_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7585 a_22386_8488# a_16746_8486# a_22294_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7586 a_30599_28023# a_28757_27247# a_30745_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7587 a_30418_21540# a_16746_21538# a_30326_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7588 VDD a_6649_25615# a_7841_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7589 a_7073_51433# a_6671_51183# a_6909_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X759 a_47486_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7590 a_28251_51727# a_27627_51733# a_28143_52105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7591 a_45782_58178# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7592 VDD a_12901_66959# a_27314_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7593 a_28714_68218# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7594 a_11074_22895# a_11574_22869# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7595 a_15212_31375# a_14361_29967# a_14939_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=3.4735e+11p ps=3.68e+06u w=650000u l=150000u
X7596 VDD a_30412_42589# a_35185_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7597 VSS a_11067_23759# a_16362_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X7598 a_19374_18528# a_16746_18526# a_19282_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7599 a_5291_56765# a_3295_54421# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X76 VDD a_16824_28309# a_15799_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X760 a_46390_68218# a_12727_67753# a_46882_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7600 a_1761_50639# a_1591_50639# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X7601 a_20378_13508# a_16746_13506# a_20286_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7602 a_27588_52271# a_8491_57487# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7603 VSS a_16824_28309# a_15799_29941# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X7604 a_11943_63125# a_12231_60949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7605 a_36395_43177# a_35463_42943# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7606 a_18944_31055# a_3339_32463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X7607 a_45478_63198# a_16746_63200# a_45386_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7608 VSS a_20623_36595# a_20563_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X7609 VSS a_10515_22671# a_22690_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X761 a_42866_7452# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7610 VSS a_12901_66665# a_36746_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7611 a_41820_41501# a_41443_41855# a_42316_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7612 a_33856_42693# a_32887_42405# a_33760_42693# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7613 a_7901_74281# a_6098_73095# a_7829_74281# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7614 a_22991_28111# a_4811_34855# a_22857_28111# VSS sky130_fd_pr__nfet_01v8 ad=2.5025e+11p pd=2.07e+06u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X7615 VSS a_11067_66191# a_12580_15939# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7616 a_28810_64524# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7617 a_25306_61190# a_12981_59343# a_25798_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7618 a_34434_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7619 a_33338_69222# a_16362_69222# a_33430_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X762 a_3137_37589# a_2971_37589# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7620 VDD a_13669_39605# a_16699_37999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7621 a_30485_49257# a_30005_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7622 a_12725_44527# a_12559_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7623 a_7987_40821# a_7847_39872# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7624 a_37446_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7625 a_27974_32459# a_26505_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X7626 a_3013_42301# a_2969_41909# a_2847_42313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7627 a_1757_71317# a_1591_71317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7628 VSS a_7925_72399# a_9161_72737# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7629 a_18770_56492# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X763 a_18674_57174# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7630 a_36442_65206# a_16746_65208# a_36350_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7631 VSS VSS a_41766_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7632 a_29322_60186# a_12727_58255# a_29814_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7633 a_35346_20902# a_16362_20536# a_35438_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7634 a_38450_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7635 a_39742_44527# a_39565_44527# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7636 a_49494_64202# a_16746_64204# a_49402_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7637 a_41370_57174# a_12257_56623# a_41862_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7638 a_30849_50959# a_30663_51727# a_30415_50871# VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X7639 a_4253_67753# a_4211_67655# a_4169_67753# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X764 a_45478_60186# a_16746_60188# a_45386_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7640 VSS a_1952_60431# a_2721_55329# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7641 a_33041_51157# a_4482_57863# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7642 a_17670_70226# a_12901_66665# a_17274_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7643 a_39454_56170# a_16746_56172# a_39362_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7644 a_31422_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7645 VSS a_12727_13353# a_44778_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7646 a_47790_18894# a_12899_10927# a_47394_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7647 a_41766_12870# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7648 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7649 a_6713_72765# a_6327_72917# a_6641_72765# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X765 VDD a_12727_58255# a_49402_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7650 VDD a_4681_13621# a_4629_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7651 a_13047_29575# a_13390_29575# a_13287_29423# VSS sky130_fd_pr__nfet_01v8 ad=3.8025e+11p pd=3.77e+06u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X7652 a_21290_9858# a_12546_22351# a_21782_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7653 a_31822_17492# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7654 a_31726_23914# a_10515_23975# a_31330_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7655 a_4818_47741# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7656 VSS a_32365_37692# a_32057_37479# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7657 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7658 vcm_commonmode a_16362_62194# a_44474_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7659 a_45386_58178# a_10515_22671# a_45878_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X766 a_45478_19532# a_16746_19530# a_45386_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7660 VSS a_12899_10927# a_17670_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7661 a_4443_46607# a_19439_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X7662 a_10509_73193# a_8003_72917# a_10509_72943# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7663 vcm_commonmode VSS a_27406_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7664 a_21686_15882# a_12877_14441# a_21290_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7665 VSS a_12877_14441# a_48794_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7666 a_45782_11866# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7667 a_31422_70226# a_16746_70228# a_31330_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7668 VDD a_6720_15279# a_6895_15253# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7669 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X767 a_20286_67214# a_16362_67214# a_20378_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7670 a_28714_21906# a_28756_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7671 a_17600_50345# a_17493_50639# a_17682_50095# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X7672 a_32334_13874# a_12727_15529# a_32826_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7673 a_13835_41001# a_13107_41317# a_14039_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7674 a_33430_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7675 a_5639_27247# a_4427_25071# a_5795_27497# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7676 a_16746_11498# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X7677 a_21382_62194# a_16746_62196# a_21290_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7678 a_22786_58500# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7679 a_37354_8854# a_12985_19087# a_37846_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X768 a_25702_58178# a_12901_58799# a_25306_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7680 a_18674_13874# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7681 a_25702_14878# a_12727_15529# a_25306_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7682 VSS a_2292_17179# a_5957_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7683 VSS a_10055_58791# a_22690_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7684 a_19374_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7685 a_15911_31784# a_2235_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7686 VDD VSS a_44382_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7687 vcm_commonmode a_16362_17524# a_31422_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7688 a_7281_29423# a_6743_29673# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7689 a_47886_8456# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X769 VSS VSS a_22690_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7690 a_43774_8854# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7691 a_37750_67214# a_12727_67753# a_37354_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7692 VSS a_11067_13095# a_34738_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7693 a_30967_41001# a_31004_40743# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X7694 a_19678_8854# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7695 a_8381_51727# a_4298_58951# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X7696 VDD a_4399_48084# a_4287_48634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7697 a_10471_65002# a_10501_65871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X7698 a_35346_65206# a_16362_65206# a_35438_65206# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7699 a_15483_49007# a_10515_63143# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=0p ps=0u w=650000u l=150000u
X77 a_17274_21906# a_11067_21583# a_17766_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X770 VSS a_13620_43047# a_12889_40977# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7700 a_45878_20504# a_43270_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7701 VDD a_10515_23975# a_48398_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7702 a_45478_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7703 VSS a_12985_19087# a_29718_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7704 VSS a_21712_43781# a_21049_41245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X7705 a_48398_64202# a_16362_64202# a_48490_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7706 VDD a_14049_40693# a_14079_41046# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7707 VSS a_1586_45431# a_9135_49557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7708 a_19780_38341# a_18811_38053# a_19684_38341# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7709 vcm_commonmode a_16362_69222# a_47486_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X771 a_29915_41959# a_30023_41959# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7710 VDD a_12877_14441# a_38358_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7711 a_35838_12472# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7712 VDD a_24800_41953# a_23901_42044# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X7713 VDD a_10531_31055# a_15548_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.65e+12p ps=1.53e+07u w=1e+06u l=150000u M=4
X7714 VDD a_10789_74273# a_10679_74397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7715 VDD a_4339_64521# a_9177_60214# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X7716 VSS a_8177_37013# a_7244_39189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7717 a_49494_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7718 a_46390_12870# a_16362_12504# a_46482_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7719 a_12507_35862# a_12325_35862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X772 a_18770_7452# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7720 a_25398_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7721 a_28902_27791# a_28817_29111# a_28599_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7722 a_35049_30511# a_34759_31029# a_34977_30511# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7723 a_42770_61190# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7724 a_34579_50613# a_35224_49871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7725 a_41462_59182# a_16746_59184# a_41370_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7726 a_8129_38377# a_5631_38127# a_7948_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.45e+11p pd=2.69e+06u as=7.55e+11p ps=3.51e+06u w=1e+06u l=150000u
X7727 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X7728 a_35438_24552# VDD a_35346_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7729 a_39362_66210# a_16362_66210# a_39454_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X773 VSS a_8625_20175# a_5211_24759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X7730 a_30715_41835# a_12357_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7731 a_4052_73865# a_3137_73493# a_3705_73461# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X7732 a_25702_71230# a_21371_50959# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7733 a_24394_69222# a_16746_69224# a_24302_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7734 a_2325_26401# a_2107_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7735 a_21187_29415# a_34482_29941# a_36199_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X7736 vcm_commonmode a_16362_66210# a_21382_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7737 a_39854_11468# a_39223_32463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7738 a_23298_24918# VSS a_23390_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7739 VDD a_12983_63151# a_33338_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X774 a_30008_30511# a_29942_30663# a_29926_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7740 VSS a_7862_34025# a_22922_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X7741 a_26310_7850# VDD a_26802_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7742 VDD a_30557_49783# a_30525_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.4e+11p ps=2.68e+06u w=1e+06u l=150000u
X7743 a_8397_35407# a_5915_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7744 VDD a_4968_60405# a_4906_60431# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X7745 a_33430_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7746 a_29414_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7747 a_26310_60186# a_16362_60186# a_26402_60186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7748 a_4681_13621# a_5227_13621# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7749 vcm_commonmode a_16362_8488# a_45478_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X775 a_18627_34239# a_16928_35303# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X7750 a_19525_28585# a_17278_28309# a_19442_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7751 a_25926_51549# a_24849_51183# a_25764_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7752 vcm_commonmode VSS a_42466_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7753 a_16362_66210# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7754 a_16948_27253# a_11430_26159# a_16865_27511# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7755 VDD a_2325_29941# a_2215_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7756 a_29718_70226# a_29760_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7757 a_28410_68218# a_16746_68220# a_28318_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7758 vcm_commonmode a_16362_65206# a_25398_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7759 VDD a_20027_27221# a_20359_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X776 a_28810_61512# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7760 VDD a_30788_28487# a_35069_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X7761 a_30722_24918# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7762 a_6649_25615# a_4528_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7763 a_27314_23914# a_16362_23548# a_27406_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7764 VDD a_10975_66407# a_37354_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7765 a_34834_62516# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7766 VDD a_12546_22351# a_29322_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7767 a_44778_58178# a_12901_58799# a_44382_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7768 a_8173_70543# a_6921_72943# a_7755_70543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X7769 a_43495_28487# a_41842_27221# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X777 a_8273_42479# a_7815_42453# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X7770 a_27267_39605# a_12641_37684# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7771 a_16961_28585# a_11902_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X7772 a_19678_62194# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7773 a_47886_61512# a_43362_28879# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7774 VSS a_12727_58255# a_23694_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7775 a_20682_16886# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7776 VSS a_11067_67279# a_23694_19898# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7777 a_8941_59663# a_5024_67885# a_7107_58487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7778 VDD a_15607_46805# a_40086_28335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7779 a_13528_36055# a_12889_35537# a_13670_36189# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X778 a_26514_47375# a_26259_47491# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X7780 vcm_commonmode a_16362_56170# a_28410_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7781 a_37750_20902# a_11067_67279# a_37354_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7782 a_33734_15882# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7783 a_30326_8854# a_16362_8488# a_30418_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7784 VDD a_20635_29415# a_33049_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X7785 a_12892_37455# a_12641_37684# a_12671_37782# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7786 a_11308_22057# a_10073_23439# a_8295_47388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X7787 a_4441_62327# a_1591_64239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7788 VDD a_12355_15055# a_24302_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7789 VSS a_2589_55535# a_2882_56989# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X779 a_34434_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7790 VDD a_9491_12297# a_10351_12879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7791 vcm_commonmode a_16362_23548# a_34434_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7792 a_2325_36469# a_2107_36873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X7793 a_1861_5059# a_1761_6031# a_1765_5059# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7794 a_2108_12015# a_1761_11471# a_1887_12342# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7795 a_4706_40847# a_4314_40821# a_4960_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X7796 VDD a_3491_42239# a_3949_41935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X7797 vcm_commonmode a_16362_22544# a_47486_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7798 a_34823_44535# a_35217_44509# a_24800_43041# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X7799 a_22063_47594# a_20853_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X78 a_23774_49551# a_23830_49525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X780 VSS a_4399_48084# a_4287_48634# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7800 VDD a_12907_56399# a_16362_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X7801 VSS a_41289_43421# a_40981_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7802 a_28810_72556# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7803 a_46390_57174# a_16362_57174# a_46482_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7804 a_4630_15823# a_3911_16065# a_4067_15797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X7805 a_8205_26409# a_4528_26159# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X7806 VSS a_10717_53113# a_10651_53181# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7807 a_22294_11866# a_16362_11500# a_22386_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7808 VDD a_12899_10927# a_40366_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7809 VDD a_12981_59343# a_28318_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X781 a_19894_51433# a_19946_51157# a_6559_59879# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X7810 a_49798_67214# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7811 VDD a_1915_11092# a_1867_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7812 a_11710_28335# a_11747_28639# a_11527_28701# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7813 a_9556_67503# a_8772_63927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7814 VDD a_33597_50141# a_33697_50359# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7815 a_41462_12504# a_16746_12502# a_41370_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7816 a_3607_34639# a_3063_34319# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X7817 VSS a_1950_59887# a_11753_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7818 a_24394_22544# a_16746_22542# a_24302_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7819 VSS a_12263_20969# a_12196_21583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X782 a_33338_66210# a_16362_66210# a_33430_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7820 a_39758_59182# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7821 VSS a_12257_56623# a_43774_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7822 a_39758_17890# a_12899_11471# a_39362_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7823 a_37354_16886# a_12899_11471# a_37846_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7824 a_49494_72234# VDD a_49402_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7825 VSS a_1586_9991# a_5363_16367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7826 a_21859_35831# a_20927_35877# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7827 VSS a_12983_63151# a_26706_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7828 a_23694_64202# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7829 a_9497_10383# a_9642_10357# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X783 a_9872_20969# a_7187_23439# a_9955_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+12p pd=1.273e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X7830 a_30722_65206# a_10975_66407# a_30326_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7831 a_4067_23145# a_2317_28892# a_3985_22901# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7832 a_21290_21906# a_11067_21583# a_21782_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7833 VSS a_21049_34717# a_20741_35077# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7834 a_21290_17890# a_16362_17524# a_21382_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7835 vcm_commonmode a_16362_61190# a_36442_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7836 a_28410_21540# a_16746_21538# a_28318_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7837 a_11067_63143# a_14634_47349# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X7838 a_5695_47919# a_5345_47919# a_5600_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X7839 a_7812_61839# a_7829_60431# a_7622_61839# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X784 a_5269_43809# a_5051_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7840 a_40458_18528# a_16746_18526# a_40366_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7841 VDD a_12901_58799# a_44382_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7842 a_12283_40183# a_12677_40157# a_12249_43457# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X7843 a_20682_57174# a_10515_22671# a_20286_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7844 a_8289_52047# a_7933_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7845 a_41427_52263# a_41059_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7846 a_15566_49257# a_5039_42167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7847 a_44778_11866# a_12985_16367# a_44382_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7848 a_21663_35327# a_17863_36595# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X7849 a_7895_47158# a_7644_46805# a_7436_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X785 VSS a_33839_28309# a_32167_29611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7850 a_18045_38017# a_18351_37503# a_19224_37479# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7851 a_12539_62063# a_11067_63143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7852 VDD a_18328_31573# a_17927_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7853 a_18370_13508# a_16746_13506# a_18278_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7854 a_27806_15484# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7855 a_13909_35395# a_18627_35327# a_19559_35561# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7856 VDD a_12877_16911# a_31330_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7857 a_8222_47741# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7858 a_12921_35279# a_12651_35645# a_12831_35645# VSS sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7859 a_48890_69544# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X786 a_19774_19500# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7860 a_45386_66210# a_10975_66407# a_45878_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X7861 a_8747_14735# a_8123_14741# a_8639_15113# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7862 a_75162_40202# a_75258_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7863 VSS a_8556_10357# a_8494_10383# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X7864 a_2325_38645# a_2107_39049# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7865 a_17670_55166# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7866 VDD a_17709_48761# a_17739_48502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7867 vcm_commonmode a_16362_14512# a_41462_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7868 VDD a_35932_37601# a_36520_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7869 vcm_commonmode a_16362_59182# a_30418_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X787 VDD VDD a_28318_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7870 a_30079_47375# a_26417_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X7871 VDD a_12985_19087# a_41370_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7872 a_41232_28879# a_28841_29575# a_41059_29199# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X7873 VDD a_1915_45908# a_1867_45743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X7874 a_28318_11866# a_10055_58791# a_28810_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7875 VDD a_4717_20961# a_4607_21085# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7876 a_37534_51701# a_37459_51183# a_38704_52047# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u M=4
X7877 a_18278_68218# a_12727_67753# a_18770_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7878 VDD a_12516_7093# a_25306_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7879 a_22786_66532# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X788 VSS VDD a_24698_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7880 a_49402_65206# a_12355_65103# a_49894_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7881 a_17366_60186# a_16746_60188# a_17274_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7882 a_9828_56311# a_8123_56399# a_9970_56445# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7883 a_17366_19532# a_16746_19530# a_17274_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7884 VSS a_8933_22583# a_10528_20495# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7885 VDD a_12985_19087# a_17274_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7886 VSS a_23631_50069# a_23577_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7887 VDD a_7637_53877# a_3228_54171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X7888 a_4941_35727# a_5079_35639# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X7889 a_22294_56170# a_16362_56170# a_22386_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X789 VDD a_4119_70741# a_7100_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X7890 a_26343_30761# a_25321_29673# a_26247_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7891 a_8891_22351# a_8015_21807# a_8671_22671# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X7892 a_39362_57174# a_12257_56623# a_39854_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7893 VDD a_7695_31573# a_12591_31029# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.646e+11p ps=2.94e+06u w=420000u l=150000u
X7894 VSS VDD a_34738_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7895 a_43870_55488# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7896 a_49798_20902# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7897 a_5258_54223# a_4889_55535# a_5089_53903# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7898 VDD a_1929_12131# a_5867_11995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7899 VSS a_10995_14333# a_10956_14459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X79 a_17274_17890# a_16362_17524# a_17366_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X790 a_2426_35951# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7900 VSS a_27983_40871# a_12663_39783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7901 a_2215_40669# a_1591_40303# a_2107_40303# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X7902 a_26802_65528# a_21371_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7903 a_23298_62194# a_12355_15055# a_23790_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7904 VSS a_6372_38279# a_6377_38133# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7905 a_24223_31171# a_23626_31573# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X7906 a_16746_19530# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X7907 a_26867_29739# a_26191_29397# a_26694_29473# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7908 a_12161_31849# a_3339_30503# a_12245_31599# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7909 VSS a_12901_66665# a_47790_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X791 VSS a_4647_63937# a_4608_63811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7910 a_39758_12870# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7911 a_45478_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7912 a_10771_25731# a_9751_25071# a_10699_25731# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X7913 VSS a_32327_40191# a_32273_40513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7914 VSS a_12985_16367# a_43774_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7915 a_32121_42369# a_32795_42943# a_33668_42919# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X7916 VDD VSS a_20286_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7917 VSS a_12985_7663# a_26706_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7918 a_41766_61190# a_12355_15055# a_41370_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7919 a_11266_10205# a_11179_9981# a_10862_10091# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X792 a_4607_21085# a_3983_20719# a_4499_20719# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X7920 a_29814_56492# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7921 a_27009_47919# a_22989_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7922 a_24698_71230# a_12947_71576# a_24302_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7923 VDD a_30440_31573# a_14287_51175# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X7924 a_47486_65206# a_16746_65208# a_47394_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7925 VDD a_13909_41923# a_40613_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X7926 VDD a_7295_44647# a_39035_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7927 a_5258_54223# a_3325_49551# a_5172_54223# VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X7928 a_36980_37253# a_36107_36965# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X7929 VSS a_17449_46831# a_18243_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X793 a_29269_44545# a_29391_44031# a_30323_44265# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X7930 a_25398_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7931 a_49494_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7932 a_46390_20902# a_16362_20536# a_46482_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7933 a_20682_10862# a_12546_22351# a_20286_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7934 a_38197_32143# a_12907_27023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7935 a_6927_56873# a_4119_70741# a_7009_56623# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X7936 a_24743_48437# a_24209_48463# a_25129_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7937 a_37446_57174# a_16746_57176# a_37354_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7938 a_38754_18894# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7939 a_6099_73193# a_6224_73095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X794 VSS a_12473_41781# a_12892_41807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X7940 a_43470_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7941 a_45782_60186# a_12981_59343# a_45386_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7942 a_45782_19898# a_12895_13967# a_45386_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7943 VSS a_12899_11471# a_42770_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7944 a_27901_52513# a_27683_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X7945 a_8332_38377# a_5363_30503# a_8228_38377# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.7e+11p ps=2.74e+06u w=1e+06u l=150000u
X7946 a_28714_70226# a_12901_66665# a_28318_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7947 a_40458_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7948 VDD a_5755_14709# a_6914_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X7949 a_13987_35862# a_12889_35537# a_13528_36055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X795 a_10528_20495# a_9955_21807# a_9263_24501# VSS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=2.4e+06u as=9.3275e+11p ps=9.37e+06u w=650000u l=150000u
X7950 a_40675_27791# a_40402_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7951 a_32555_43777# a_12357_37999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7952 a_30375_51335# a_2775_46025# a_30542_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7953 a_33430_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7954 vcm_commonmode a_16362_17524# a_29414_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7955 VSS a_5791_43541# a_5725_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7956 a_14365_46805# a_5039_42167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X7957 a_13097_40719# a_12831_41085# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7958 vcm_commonmode a_16362_12504# a_30418_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7959 vcm_commonmode a_16362_63198# a_42466_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X796 a_37750_23914# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X7960 a_18674_62194# a_12981_62313# a_18278_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7961 a_24208_39453# a_19629_39631# a_23987_39126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7962 a_43378_59182# a_12901_58799# a_43870_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7963 a_36842_7452# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7964 VSS a_8575_74853# a_11477_69679# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7965 a_32730_57174# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7966 VSS a_22151_29941# a_22097_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7967 VDD a_25417_51425# a_25307_51549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7968 a_34834_70548# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7969 a_36725_27497# a_20359_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X797 VDD a_18105_40157# a_17711_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X7970 a_35615_30199# a_33641_29967# a_35849_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7971 VDD VDD a_46390_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7972 VSS a_33080_37149# a_33727_36649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X7973 a_6607_13879# a_4429_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7974 VSS VDD a_42770_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7975 a_7773_63927# a_10607_58799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u M=2
X7976 a_1925_22583# a_2021_22325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7977 a_34342_60186# a_16362_60186# a_34434_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7978 VSS a_17475_51157# a_17409_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7979 a_4333_22671# a_3143_22364# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X798 a_28943_42089# a_28011_41855# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X7980 a_41351_39141# a_40403_37683# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X7981 a_20778_59504# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7982 a_44474_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7983 a_5343_72221# a_1923_73087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X7984 a_17274_70226# a_16362_70226# a_17366_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X7985 a_23498_28585# a_17869_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.55e+11p pd=5.31e+06u as=0p ps=0u w=1e+06u l=150000u
X7986 a_2663_43541# a_2872_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X7987 VSS a_8491_57487# a_9370_58575# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7988 a_2111_38279# a_2339_38129# a_2285_38155# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7989 a_15457_46831# a_10515_63143# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X799 VSS a_11067_21583# a_41766_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7990 a_9589_63401# a_3024_67191# a_9505_63401# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7991 VSS VDD a_18674_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X7992 a_10476_74031# a_10239_74575# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X7993 a_32426_62194# a_16746_62196# a_32334_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X7994 VSS a_12621_44099# a_22411_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X7995 a_2557_64239# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7996 a_6008_69679# a_3143_66972# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.46e+11p pd=5.58e+06u as=0p ps=0u w=650000u l=150000u M=2
X7997 VDD a_12546_22351# a_37354_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7998 a_23694_9858# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7999 a_28714_7850# VDD a_28318_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_7803_55509# a_8307_66415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X80 a_21290_70226# a_12516_7093# a_21782_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X800 a_38450_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8000 a_35742_68218# a_12901_66959# a_35346_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8001 VSS a_23395_32463# a_43439_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8002 a_8105_21263# a_7757_21379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X8003 a_48794_67214# a_12727_67753# a_48398_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8004 VSS a_11067_13095# a_45782_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8005 vcm_commonmode a_16362_66210# a_19374_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8006 VSS a_1586_36727# a_1683_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8007 a_23390_64202# a_16746_64204# a_23298_64202# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8008 a_46390_65206# a_16362_65206# a_46482_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8009 VSS a_6521_58773# a_5612_58229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X801 VDD a_18848_27765# a_17358_31069# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8010 a_38754_59182# a_12727_58255# a_38358_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8011 VSS a_12947_56817# a_35742_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8012 VDD a_12355_15055# a_32334_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8013 a_9782_71311# a_9063_71553# a_9219_71285# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X8014 a_12541_63401# a_10515_63143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8015 VDD a_12727_13353# a_36350_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8016 a_6457_64239# a_1823_76181# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X8017 a_7030_31055# a_6243_30662# a_6917_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X8018 VDD a_12877_14441# a_49402_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8019 a_37446_10496# a_16746_10494# a_37354_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X802 VSS a_1586_40455# a_1775_47381# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8020 VDD a_8643_48767# a_8630_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8021 vcm_commonmode VSS a_34434_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8022 VDD a_18979_30287# a_33603_47081# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X8023 a_4797_62063# a_4441_62327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8024 VSS a_16101_31029# a_18637_29451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8025 a_40762_62194# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8026 VDD a_15607_46805# a_38295_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X8027 a_37354_67214# a_16362_67214# a_37446_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8028 VSS VSS a_39758_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8029 a_44474_7484# VDD a_44382_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X803 a_44874_57496# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8030 a_23385_31171# a_22399_32143# a_23303_31171# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8031 a_23694_72234# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8032 a_32334_55166# a_11067_47695# a_32826_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8033 a_26433_39631# a_26267_39631# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X8034 a_5073_27247# a_4807_27613# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8035 a_41862_24520# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8036 a_25447_36919# a_25484_37253# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X8037 VSS a_5779_75093# a_5483_74244# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8038 VDD a_12983_63151# a_44382_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8039 VSS a_12815_19319# a_12815_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X804 a_27183_44581# a_23567_44211# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X8040 VSS a_1586_40455# a_1591_40303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8041 a_32730_10862# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8042 vcm_commonmode a_16362_9492# a_25398_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8043 VDD a_29545_35841# a_30080_36391# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8044 a_16666_55166# VSS a_16270_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8045 a_18627_35327# a_15011_34717# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X8046 a_44474_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8047 a_5441_27791# a_5175_27791# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8048 VSS a_12981_59343# a_30722_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8049 a_33689_29423# a_33694_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X805 a_27806_67536# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8050 a_27406_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8051 VSS a_4578_40455# a_4941_35727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8052 a_29147_50069# a_29561_49667# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X8053 a_28056_44869# a_28152_44869# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8054 VDD a_11035_47893# a_11022_48285# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8055 a_12226_57711# a_2419_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8056 a_42374_20902# a_12985_7663# a_42866_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8057 a_42374_16886# a_16362_16520# a_42466_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8058 a_17670_63198# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8059 VDD a_10975_66407# a_48398_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X806 a_20027_27221# a_7571_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8060 a_45878_62516# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8061 a_13015_43493# a_12249_43457# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X8062 VSS a_19594_35823# a_23451_35823# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8063 a_8056_13967# a_8026_13885# a_7953_13967# VSS sky130_fd_pr__nfet_01v8 ad=5.6875e+11p pd=4.35e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X8064 vcm_commonmode a_16362_57174# a_26402_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8065 a_4214_73487# a_3137_73493# a_4052_73865# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8066 a_32334_72234# VSS a_32426_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8067 a_35742_21906# a_12985_7663# a_35346_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8068 a_2713_35925# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8069 a_7155_43567# a_6269_43567# a_6792_43719# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X807 VDD a_10975_66407# a_31330_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8070 VDD a_4351_67279# a_23753_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8071 a_30418_55166# VDD a_30326_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8072 a_31726_16886# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8073 a_32951_27247# a_20359_29199# a_32862_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X8074 VDD a_10515_22671# a_38358_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8075 a_48890_14480# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8076 a_48794_20902# a_11067_67279# a_48398_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8077 VDD a_10515_23975# a_22294_23914# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8078 VDD clk_vcm a_77664_40024# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8079 VDD config_2_in[2] a_1591_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X808 VSS a_3020_54135# a_2327_54135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8080 a_22294_64202# a_16362_64202# a_22386_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8081 a_43774_69222# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8082 VSS a_8117_30287# a_8561_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X8083 a_7640_42479# a_6725_42479# a_7293_42721# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X8084 VDD a_1586_18695# a_1591_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8085 a_22132_40865# a_21479_40229# a_22352_40517# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8086 a_38754_12870# a_10055_58791# a_38358_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8087 VDD a_26397_51183# a_31186_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8088 vcm_commonmode a_16362_23548# a_45478_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8089 a_19282_21906# a_11067_21583# a_19774_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X809 VDD a_39836_38567# a_39740_38567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X8090 VSS a_41289_36893# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X8091 a_3449_54201# a_2840_53511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8092 a_23298_70226# a_12516_7093# a_23790_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8093 a_19282_17890# a_16362_17524# a_19374_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8094 VDD a_12727_15529# a_25306_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8095 a_49402_10862# a_12985_16367# a_49894_10464# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8096 a_23390_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8097 a_20286_12870# a_16362_12504# a_20378_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8098 a_48398_9858# a_16362_9492# a_48490_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8099 VSS a_12901_66959# a_20682_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X81 VDD a_12727_15529# a_23298_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X810 VDD a_6515_62037# a_7289_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.6e+11p ps=7.72e+06u w=1e+06u l=150000u
X8100 a_5259_39367# a_4314_40821# a_5426_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X8101 a_47790_68218# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8102 a_38450_18528# a_16746_18526# a_38358_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8103 vcm_commonmode a_16362_15516# a_35438_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8104 a_33338_11866# a_16362_11500# a_33430_11500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8105 VDD a_38076_31573# a_30788_28487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8106 a_11521_58951# a_11943_63125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8107 a_4517_26703# a_3301_27791# a_4433_26703# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8108 a_5453_72097# a_5235_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X8109 a_11429_16367# a_10239_16367# a_11320_16367# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X811 a_27314_57174# a_16362_57174# a_27406_57174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8110 a_22386_23548# a_16746_23546# a_22294_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8111 VDD a_2672_45577# a_2847_45503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8112 a_11396_55535# a_8199_58229# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X8113 a_36615_29199# a_11067_46823# a_36425_28879# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X8114 a_2215_12559# a_1591_12565# a_2107_12937# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X8115 a_35438_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8116 a_26802_10464# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8117 VSS a_10515_32143# a_12244_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8118 VSS a_10515_22671# a_41766_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8119 a_10515_32143# a_4903_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X812 VDD config_2_in[1] a_1591_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X8120 VSS a_12727_67753# a_24698_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8121 a_8577_48841# a_7387_48469# a_8468_48841# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X8122 a_21686_65206# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8123 a_44382_61190# a_12981_59343# a_44874_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8124 vcm_commonmode a_16362_14512# a_39454_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8125 VSS a_13835_36649# a_16707_36919# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8126 a_8485_71855# a_8539_71829# a_8497_72105# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8127 a_48398_16886# a_12899_11471# a_48890_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8128 VSS a_10286_26311# a_10521_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8129 VDD a_2191_68565# a_4719_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X813 VDD a_2971_48463# a_2595_47653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8130 a_2369_51183# a_2325_51425# a_2203_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X8131 a_35346_19898# a_11067_67279# a_35838_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8132 VDD a_22989_48437# a_25961_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X8133 VSS a_21856_36513# a_20957_36604# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=3.83e+06u
X8134 a_10317_67191# a_10379_66389# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8135 a_19675_49525# a_19878_49683# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8136 a_39454_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8137 VDD a_2787_30503# a_26191_29397# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X8138 a_32730_71230# a_12947_71576# a_32334_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8139 a_1643_29397# a_1799_29556# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X814 a_31422_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8140 a_4989_42255# a_4446_40553# a_4771_42167# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8141 a_17274_63198# a_12981_62313# a_17766_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8142 a_14625_30761# a_10531_31055# a_14471_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8143 a_16746_60188# a_11803_55311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8144 a_22749_50613# a_22531_51017# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8145 VSS a_12901_58799# a_27710_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8146 VDD a_11067_46823# a_41211_28023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8147 a_11902_46831# a_4674_40277# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8148 a_21782_61512# a_17507_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8149 a_16362_14512# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X815 a_47790_15882# a_12877_14441# a_47394_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8150 a_3583_37961# a_3137_37589# a_3487_37961# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=360000u l=150000u
X8151 a_31726_57174# a_10515_22671# a_31330_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8152 a_10557_47919# a_10513_48161# a_10391_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X8153 a_25798_16488# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8154 a_18851_51017# a_18501_50645# a_18756_51005# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X8155 a_35529_27497# a_20359_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8156 a_20713_40193# a_21387_39679# a_22319_39913# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8157 VSS a_38345_42044# a_38037_41831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8158 a_43378_67214# a_12983_63151# a_43870_67536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8159 a_29414_13508# a_16746_13506# a_29322_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X816 VSS a_12877_16911# a_44778_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8160 vcm_commonmode a_16362_10496# a_26402_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8161 a_6980_45565# a_6361_44655# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8162 a_29679_37737# a_29361_38017# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X8163 VSS a_15253_43421# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X8164 VSS a_2012_33927# a_2568_29245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8165 VDD a_5915_35943# a_8395_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X8166 a_4693_36611# a_3305_38671# a_4621_36611# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8167 a_5731_37039# a_5701_37013# a_5625_37039# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8168 a_29887_32375# a_30052_32117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8169 a_40895_43447# a_39244_41953# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X817 a_17365_49007# a_17321_49249# a_17199_49007# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X8170 a_28714_55166# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8171 a_2847_23743# a_2672_23817# a_3026_23805# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8172 a_43774_22910# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8173 VSS a_16928_42919# a_16891_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8174 a_21169_49007# a_21003_49007# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8175 a_20993_28879# a_10873_27497# a_20747_27765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8176 a_20778_67536# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8177 VSS a_36600_49159# a_36551_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8178 a_10328_21379# a_10275_21495# a_10233_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X8179 a_30326_24918# VSS a_30818_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X818 VDD a_10515_22671# a_21290_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8180 a_2125_34863# a_2011_34837# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8181 a_29829_29673# a_4811_34855# a_28963_28853# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8182 a_20286_57174# a_16362_57174# a_20378_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8183 VSS a_12899_10927# a_36746_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8184 a_40762_15882# a_12877_14441# a_40366_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8185 a_4031_50247# a_4127_50069# a_4429_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X8186 a_33338_56170# a_16362_56170# a_33430_56170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8187 VSS a_10515_23975# a_20682_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8188 VDD a_4685_37583# a_7847_39872# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8189 a_17366_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X819 a_26310_7850# VSS a_26402_7484# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8190 a_47790_21906# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8191 VSS a_12546_22351# a_33734_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8192 VSS VDD a_45782_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8193 VDD a_9707_73807# a_10109_73487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8194 a_41862_58500# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8195 a_37750_13874# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8196 result_out[9] a_1644_66933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8197 a_23390_72234# VDD a_23298_72234# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8198 a_8494_10383# a_7775_10625# a_7931_10357# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8199 VSS a_10055_58791# a_41766_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X82 a_47394_10862# a_12985_16367# a_47886_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X820 VSS a_10515_23975# a_27710_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8200 a_38450_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8201 a_43774_9858# a_12985_19087# a_43378_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8202 VDD a_3983_12015# a_3843_13880# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8203 a_12056_55535# a_10975_55535# a_11709_55777# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8204 a_27710_24918# VSS a_27314_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8205 a_24302_15882# a_12727_13353# a_24794_15484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8206 VSS a_11067_21583# a_24698_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8207 a_12056_65327# a_11141_65327# a_11709_65569# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8208 VSS a_26397_51183# a_32401_49871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8209 a_27806_57496# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X821 a_5265_28157# a_4995_27791# a_5175_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8210 VDD a_37427_47893# a_39127_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8211 a_1849_52271# a_1683_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8212 a_30843_52521# a_28881_52271# a_30625_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8213 VSS a_7571_31599# a_8197_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X8214 VDD VSS a_31330_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8215 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8216 a_17670_16886# a_12727_13353# a_17274_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8217 a_2080_64605# a_1643_64213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8218 a_6373_69679# a_5438_69679# a_6008_69679# VSS sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u M=2
X8219 a_9223_22895# a_5531_22895# a_9135_22895# VSS sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=0p ps=0u w=650000u l=150000u
X822 a_36746_70226# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8220 VSS a_12047_57685# a_11981_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8221 VSS a_11053_62607# a_11801_64015# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X8222 a_32917_35307# a_30757_37455# a_32831_35307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8223 VSS a_12877_16911# a_27710_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8224 VSS a_12981_62313# a_39758_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8225 a_36746_60186# a_36717_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8226 a_35438_58178# a_16746_58180# a_35346_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8227 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8228 a_36746_19898# a_36629_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8229 a_31726_10862# a_12546_22351# a_31330_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X823 a_35438_68218# a_16746_68220# a_35346_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8230 a_6257_23145# a_5085_23047# a_6185_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8231 VSS a_4351_26703# a_9528_25071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8232 a_20027_27221# a_7571_29199# a_20635_27247# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8233 a_18770_59504# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8234 a_19559_43177# a_19596_42919# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X8235 a_10339_14735# a_9865_14441# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8236 VDD a_13620_36519# a_12889_35537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8237 a_16744_40517# a_15775_40229# a_16707_40183# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8238 a_8377_24847# a_5449_25071# a_8031_24527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X8239 VDD a_20103_30287# a_20505_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 a_31822_14480# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8240 vcm_commonmode a_16362_18528# a_27406_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8241 a_37846_22512# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8242 a_40858_8456# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8243 VSS a_2419_48783# a_11569_57711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8244 a_2748_68565# a_2927_68565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8245 a_31422_16520# a_16746_16518# a_31330_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8246 VDD a_11067_67279# a_41370_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8247 VDD a_33939_43439# a_34045_43439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8248 a_42997_47081# a_18979_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8249 a_44474_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X825 a_31726_20902# a_11067_67279# a_31330_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8250 a_41370_61190# a_16362_61190# a_41462_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8251 VDD a_14131_44135# a_13944_43957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8252 a_29718_62194# a_12981_62313# a_29322_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8253 a_30722_58178# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8254 a_2203_51183# a_1757_51183# a_2107_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8255 a_44778_71230# a_39299_48783# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8256 a_43470_69222# a_16746_69224# a_43378_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8257 vcm_commonmode a_16362_66210# a_40458_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8258 VSS a_8933_22583# a_11049_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8259 a_33764_41831# a_32795_41855# a_33668_41831# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X826 a_8222_47414# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X8260 VDD a_3983_16617# a_4630_15823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8261 VDD a_19885_50095# a_20914_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8262 VDD a_12947_8725# a_26310_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8263 VSS a_12985_19087# a_22690_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8264 a_42374_24918# VSS a_42466_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8265 a_2004_42453# a_2012_33927# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8266 a_45878_70548# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8267 a_38358_14878# a_16362_14512# a_38450_14512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8268 VSS a_7896_18695# a_7059_24135# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8269 a_42466_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X827 VSS a_4571_26677# a_8205_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.72e+11p ps=4.36e+06u w=650000u l=150000u
X8270 VDD a_11719_28023# a_14553_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8271 a_48490_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8272 a_45386_60186# a_16362_60186# a_45478_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8273 a_7460_31055# a_6835_31055# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8274 a_30418_63198# a_16746_63200# a_30326_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8275 a_10391_47919# a_9945_47919# a_10295_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8276 a_5737_75369# a_2451_72373# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8277 a_28318_70226# a_16362_70226# a_28410_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8278 a_5320_18231# a_3325_18543# a_5462_18365# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8279 a_18016_46983# a_12447_29199# a_18158_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X828 vcm_commonmode VSS a_40458_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8280 VSS a_12901_66665# a_21686_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8281 a_6757_65327# a_6722_65579# a_6519_65301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8282 VDD a_12985_16367# a_35346_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8283 vcm_commonmode a_16362_65206# a_44474_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8284 VSS a_2744_66103# a_1915_67477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8285 VDD a_7803_55509# a_9280_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.85e+11p ps=5.37e+06u w=1e+06u l=150000u
X8286 VSS a_2099_59861# a_2327_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X8287 VDD a_12985_7663# a_18278_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8288 VDD a_12546_22351# a_48398_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8289 VSS a_28757_27247# a_32507_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X829 VDD a_32327_35839# a_32187_36161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8290 a_4717_48437# a_4499_48841# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8291 a_18278_62194# a_16362_62194# a_18370_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8292 a_22386_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8293 vcm_commonmode a_16362_57174# a_34434_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8294 a_40981_43781# a_39244_41953# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8295 a_1644_74005# a_1591_64239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8296 a_46786_68218# a_12901_66959# a_46390_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8297 a_7873_46653# a_7494_46287# a_7801_46653# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=0p ps=0u w=420000u l=150000u
X8298 a_28909_49871# a_29055_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8299 a_2739_22895# a_2317_28892# a_2376_23047# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X83 a_21382_15516# a_16746_15514# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X830 vcm_commonmode a_16362_18528# a_44474_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8300 vcm_commonmode a_16362_67214# a_17366_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8301 VDD a_1586_66567# a_3983_65327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8302 a_21382_65206# a_16746_65208# a_21290_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8303 a_3141_59887# a_2785_60151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8304 vcm_commonmode a_16362_56170# a_47486_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8305 a_21261_47919# a_21095_47919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8306 a_6817_42255# a_6269_43567# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8307 a_1908_17141# a_2283_15797# a_2229_16143# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8308 a_20286_20902# a_16362_20536# a_20378_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8309 a_23390_23548# a_16746_23546# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X831 VSS a_3949_41935# a_6514_37191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X8310 a_19374_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8311 a_39854_63520# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8312 a_19096_44129# a_18627_44581# a_19500_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8313 a_49798_59182# a_12727_58255# a_49402_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8314 VDD a_12355_15055# a_43378_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8315 a_35438_11500# a_16746_11498# a_35346_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8316 VSS a_12981_59343# a_28714_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8317 a_24394_56170# a_16746_56172# a_24302_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8318 a_25702_17890# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8319 VDD a_12895_13967# a_34342_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X832 a_48890_58500# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8320 a_4885_71855# a_4719_71855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8321 VDD a_31648_43781# a_31552_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8322 a_13049_31627# a_8461_32937# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8323 a_22338_48285# a_21261_47919# a_22176_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8324 a_35346_68218# a_16362_68218# a_35438_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8325 a_24394_8488# a_16746_8486# a_24302_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8326 VDD a_75475_38962# a_76180_38962# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8327 a_10789_74273# a_10571_74031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8328 a_7050_53333# a_17843_48981# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X8329 a_4035_33205# a_4191_33449# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X833 VSS a_23565_38565# a_23599_38007# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8330 a_30816_37253# a_27652_38237# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8331 a_2557_63151# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8332 a_48398_67214# a_16362_67214# a_48490_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8333 a_31171_27412# a_31263_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X8334 VDD a_12981_59343# a_47394_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8335 VDD a_20505_29967# a_22535_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X8336 a_8399_49159# a_8143_48246# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8337 VDD a_6559_59879# a_7901_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8338 a_5785_25321# a_5211_24759# a_5363_25321# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X8339 a_30326_58178# a_10515_22671# a_30818_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X834 a_21686_12870# a_10055_58791# a_21290_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8340 a_28410_55166# VDD a_28318_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8341 a_29718_16886# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8342 a_9735_63669# a_11759_63927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8343 VDD a_1929_10651# a_5775_12649# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8344 a_30722_11866# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8345 a_27314_10862# a_16362_10496# a_27406_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8346 a_43470_22544# a_16746_22542# a_43378_22910# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8347 a_17274_71230# a_12901_66665# a_17766_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8348 a_38358_59182# a_16362_59182# a_38450_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8349 a_42466_57174# a_16746_57176# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X835 a_33734_63198# a_15439_49525# a_33338_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8350 VSS a_1586_9991# a_4075_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8351 a_25398_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8352 a_4427_30511# a_3983_30761# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8353 VDD a_8543_36469# a_8423_39367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8354 a_1586_45431# a_7295_43031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8355 a_42770_64202# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8356 VSS a_24703_35823# a_16510_8760# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X8357 a_34222_43439# a_34045_43439# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8358 VSS a_24055_36415# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X8359 a_40366_21906# a_11067_21583# a_40858_21508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X836 VSS a_10055_58791# a_48794_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8360 a_7755_38991# a_6372_38279# VSS VSS sky130_fd_pr__nfet_01v8 ad=5.6875e+11p pd=4.35e+06u as=0p ps=0u w=650000u l=150000u
X8361 a_40366_17890# a_16362_17524# a_40458_17524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8362 a_2107_45577# a_1591_45205# a_2012_45565# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X8363 VDD a_12447_29199# a_40383_29575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8364 VDD a_33856_44869# a_33760_44869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8365 a_28714_63198# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8366 a_4798_23759# a_4852_23413# a_4627_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X8367 a_26815_42405# a_23567_42035# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X8368 vcm_commonmode a_16362_71230# a_38450_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8369 a_10863_16733# a_10239_16367# a_10755_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X837 VSS a_77972_39480# a_77918_39826# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8370 a_33830_16488# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8371 VSS a_12901_66959# a_18674_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8372 a_22690_67214# a_12727_67753# a_22294_67214# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8373 a_4312_51005# a_3983_50095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8374 a_13390_29575# a_15207_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8375 a_46882_15484# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8376 vcm_commonmode a_16362_10496# a_34434_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8377 a_46786_21906# a_12985_7663# a_46390_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8378 a_17682_50095# a_7050_53333# a_18034_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8379 a_43378_12870# a_12877_16911# a_43870_12472# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X838 a_6619_47607# a_4443_46607# a_6793_47713# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8380 VDD a_10515_22671# a_49402_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8381 vcm_commonmode a_16362_20536# a_17366_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8382 a_8143_48246# a_6831_63303# a_8143_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8383 a_20286_65206# a_16362_65206# a_20378_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8384 a_26310_22910# a_10515_23975# a_26802_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8385 VDD a_1586_18695# a_8123_14741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8386 a_19374_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8387 a_16270_55166# VSS a_16362_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8388 a_30818_20504# a_30764_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8389 VSS a_4578_40455# a_4443_36611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X839 a_7387_69929# a_2686_70223# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.39e+12p pd=1.278e+07u as=0p ps=0u w=1e+06u l=150000u M=2
X8390 a_30418_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8391 a_33338_64202# a_16362_64202# a_33430_64202# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8392 a_36746_13874# a_12877_16911# a_36350_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8393 a_18430_32143# a_17711_32385# a_17867_32117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X8394 a_25879_48169# a_6835_46823# a_25961_47919# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X8395 a_19678_65206# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8396 a_36671_39913# a_35739_39679# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8397 VDD a_7464_39215# a_7847_40847# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8398 vcm_commonmode VSS a_43470_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8399 a_19774_17492# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X84 VDD a_11067_47695# a_12899_3855# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X840 a_18278_55166# a_18602_55312# a_18770_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8400 a_19678_23914# a_10515_23975# a_19282_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8401 VDD a_12877_14441# a_23298_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8402 a_49798_12870# a_10055_58791# a_49402_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8403 a_20778_12472# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8404 a_17274_18894# a_16362_18528# a_17366_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8405 vcm_commonmode a_16362_69222# a_32426_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8406 a_47394_11866# a_10055_58791# a_47886_11468# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8407 VSS a_19591_50943# a_19525_51017# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X8408 a_11710_28335# a_10873_27497# a_11626_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8409 a_37354_68218# a_12727_67753# a_37846_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X841 a_2004_42453# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8410 VSS a_9123_57399# a_3714_58345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8411 a_41862_66532# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8412 a_23298_9858# a_12546_22351# a_23790_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8413 a_36442_60186# a_16746_60188# a_36350_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8414 VDD a_6372_38279# a_7999_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X8415 a_36442_19532# a_16746_19530# a_36350_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8416 a_28056_43781# a_13835_43177# VDD VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8417 a_31330_12870# a_16362_12504# a_31422_12504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8418 a_19374_70226# a_16746_70228# a_19282_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8419 a_49494_18528# a_16746_18526# a_49402_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X842 VDD a_11999_67477# a_11947_68279# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8420 vcm_commonmode a_16362_15516# a_46482_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8421 a_20378_24552# VDD a_20286_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8422 a_24302_66210# a_16362_66210# a_24394_66210# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8423 a_26345_40871# a_26550_40871# a_26508_40969# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8424 a_18413_47919# a_18243_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X8425 a_6921_23555# a_5839_22351# a_6825_23555# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X8426 VSS a_18695_47349# a_18626_47375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X8427 a_24794_11468# a_24740_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8428 a_1803_19087# a_1626_19087# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8429 a_3026_21807# a_2411_19605# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X843 VDD a_7896_18695# a_7059_24135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8430 a_15131_39997# a_14951_39997# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8431 a_42374_62194# a_12355_15055# a_42866_62516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8432 VDD a_5064_65327# a_5239_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8433 VDD a_6260_47919# a_6435_47893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8434 VDD a_38044_44759# a_37857_44501# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8435 a_9364_71311# a_9150_71311# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8436 a_39362_8854# a_12985_19087# a_39854_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8437 VSS a_25221_41281# a_25355_40183# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8438 a_2411_26133# a_2327_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u M=4
X8439 a_46390_19898# a_11067_67279# a_46882_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X844 VSS a_1586_40455# a_3983_48469# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8440 VSS a_2315_24540# a_3529_25731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8441 a_33041_51157# a_33313_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X8442 a_18770_67536# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8443 a_33593_31287# a_27535_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8444 a_49894_8456# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8445 a_45782_8854# a_43270_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8446 a_11183_30761# a_9367_29397# a_11377_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=0p ps=0u w=1e+06u l=150000u
X8447 VDD a_10975_66407# a_22294_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8448 a_48890_56492# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8449 a_43774_71230# a_12947_71576# a_43378_71230# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X845 a_41370_71230# a_16362_71230# a_41462_71230# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8450 a_76346_38962# a_76180_38962# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8451 a_28318_63198# a_12981_62313# a_28810_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8452 a_32826_61512# a_28547_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8453 VDD a_35033_37692# a_34639_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8454 VSS a_2191_68565# a_4719_51183# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8455 a_27406_14512# a_16746_14510# a_27314_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8456 VSS a_10515_23975# a_18674_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8457 a_22690_20902# a_11067_67279# a_22294_20902# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8458 a_32218_49257# a_32134_49159# a_32135_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8459 VDD a_10288_17143# a_10239_16911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X846 a_46786_62194# a_12981_62313# a_46390_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8460 a_23685_29111# a_23734_29941# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8461 VDD a_12257_56623# a_25306_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8462 a_39454_67214# a_16746_67216# a_39362_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8463 vcm_commonmode a_16362_64202# a_36442_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8464 a_47790_70226# a_12901_66665# a_47394_70226# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8465 VSS a_3327_9308# a_9179_13737# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8466 a_29205_34215# a_29513_34428# a_27560_34337# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X8467 a_41766_23914# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8468 a_16746_57176# a_11803_55311# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X8469 a_38358_22910# a_16362_22544# a_38450_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X847 a_32334_10862# a_12985_16367# a_32826_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8470 a_42466_20536# a_16746_20534# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8471 a_28115_34743# a_27183_34789# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X8472 a_8117_30287# a_4248_29967# a_8129_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8473 VSS a_6177_61127# a_5653_60039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8474 a_5239_45717# a_2292_43291# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8475 a_37750_62194# a_12981_62313# a_37354_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8476 a_32730_8854# a_12947_8725# a_32334_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8477 a_10338_19631# a_5535_18012# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8478 VSS a_12895_13967# a_34738_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8479 a_7749_37903# a_6786_37557# a_7761_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X848 VDD a_20635_29415# a_40133_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X8480 a_9468_57487# a_9599_57141# a_9278_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8481 VDD a_13909_35395# a_19500_35303# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8482 vcm_commonmode a_16362_22544# a_32426_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8483 a_1915_21482# a_2007_21237# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8484 a_31330_57174# a_16362_57174# a_31422_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8485 VSS a_12899_10927# a_47790_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8486 a_11611_12252# a_11455_12157# a_11756_12381# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X8487 VSS a_76082_39738# a_75824_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8488 VSS a_1923_59583# a_3905_60797# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8489 a_7299_59887# a_7580_61751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X849 a_26402_7484# VDD a_26310_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8490 a_5135_50069# a_5147_50943# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8491 a_20153_49917# a_19675_49525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8492 a_10526_21807# a_6559_22671# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8493 VSS a_30311_35877# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X8494 a_19416_51017# a_18335_50645# a_19069_50613# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8495 VDD a_9031_54135# a_6236_54421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8496 a_28318_7850# VDD a_28810_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8497 a_35742_14878# a_35601_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8498 a_16746_22542# a_16510_8760# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X8499 a_5823_57961# a_4119_70741# a_5905_57961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 a_28318_9858# a_16362_9492# a_28410_9492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X850 vcm_commonmode a_16362_61190# a_17366_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8500 a_24698_59182# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8501 vcm_commonmode a_16362_8488# a_47486_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8502 a_18674_24918# a_18007_27441# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u M=2
X8503 a_3005_56079# a_2727_56417# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X8504 a_24698_17890# a_12899_11471# a_24302_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8505 a_48794_13874# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8506 a_3578_25625# a_2223_28617# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8507 a_22294_16886# a_12899_11471# a_22786_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8508 a_2557_59709# a_1923_59583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8509 a_49494_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X851 a_29718_72234# VDD a_29322_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8510 VSS a_1915_11092# a_1867_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8511 a_39854_71552# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8512 a_30035_44581# a_29269_44545# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X8513 a_34434_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8514 a_39362_61190# a_16362_61190# a_39454_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8515 a_14830_48463# a_11067_13095# a_14524_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8516 VSS a_11710_58487# a_11981_57487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X8517 vcm_commonmode a_16362_61190# a_21382_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8518 a_5731_40079# a_4314_40821# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8519 a_4472_54991# a_4035_54965# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X852 a_4036_51157# a_4215_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8520 a_6821_26311# a_5085_24759# a_6984_26409# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8521 a_28714_16886# a_12727_13353# a_28318_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8522 VSS a_12727_15529# a_25702_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8523 a_11851_64391# a_11710_58487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X8524 a_27652_38237# a_29943_36965# a_30875_36919# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8525 VDD a_11964_18543# a_12139_18517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8526 a_32334_8854# a_16362_8488# a_32426_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8527 VSS a_2959_47113# a_35337_52093# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X8528 a_16362_61190# a_12907_56399# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X8529 a_7187_20719# a_6743_20969# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X853 a_2629_59709# a_2250_59343# a_2557_59709# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8530 VSS a_10975_66407# a_37750_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8531 a_30326_66210# a_10975_66407# a_30818_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8532 VSS a_6651_31599# a_2235_30503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X8533 a_28410_63198# a_16746_63200# a_28318_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8534 a_41766_64202# a_12355_65103# a_41370_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8535 vcm_commonmode a_16362_60186# a_25398_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8536 a_29814_59504# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8537 vcm_commonmode a_16362_19532# a_25398_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8538 a_35838_23516# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8539 a_35438_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X854 a_30722_68218# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8540 a_23905_28129# a_9529_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8541 a_21686_7850# VDD a_21290_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8542 a_39454_20536# a_16746_20534# a_39362_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8543 a_42466_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8544 VDD a_2989_45717# a_3019_46070# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8545 a_22411_40183# a_21479_40229# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X8546 result_out[8] a_1644_65845# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8547 a_2107_21807# a_1591_21807# a_2012_21807# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X8548 VSS a_20827_37737# a_22127_37737# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X8549 a_42770_72234# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X855 a_10957_57711# a_10791_57711# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8550 a_4043_44343# a_3247_20495# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8551 a_5441_72399# a_5087_72512# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X8552 a_14679_31288# a_10531_31055# a_15212_31375# VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=150000u
X8553 a_36350_15882# a_16362_15516# a_36442_15516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8554 a_39454_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8555 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8556 a_40458_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8557 VSS a_4242_35407# a_4314_40821# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8558 a_18579_27399# a_10873_27497# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8559 a_19877_52245# a_19591_50943# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X856 VSS a_3325_29967# a_4903_29975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8560 a_24302_57174# a_12257_56623# a_24794_57496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8561 a_3391_15797# a_3594_15955# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8562 a_30745_27791# a_18703_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8563 a_25019_47679# a_24844_47753# a_25198_47741# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8564 a_33430_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8565 a_35742_55166# VSS a_35346_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8566 VSS a_1915_45908# a_1867_45743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8567 a_26112_30663# a_14926_31849# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X8568 VSS a_38115_52263# a_39219_52271# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8569 a_1761_34319# a_1591_34319# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X857 VDD a_12901_58799# a_25306_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8570 a_7999_40553# a_7097_40303# a_7905_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X8571 VDD a_24497_47349# a_24387_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8572 a_18674_65206# a_10975_66407# a_18278_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8573 a_46482_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8574 VDD a_42188_43677# a_41289_43421# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X8575 VSS a_12901_66665# a_32730_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8576 a_9123_55223# a_9695_54965# a_9468_55311# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X8577 VDD a_12985_16367# a_46390_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8578 VSS a_2847_21781# a_2781_21807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X8579 VSS a_13957_36121# a_13891_36189# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X858 a_21382_18528# a_16746_18526# a_21290_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8580 VDD a_12901_66959# a_36350_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8581 VDD a_12907_56399# a_16362_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X8582 VDD a_7523_62581# a_7289_62607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8583 a_24698_12870# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8584 a_30418_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8585 VDD a_12985_7663# a_29322_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8586 VDD a_19442_28585# a_19459_29423# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X8587 VSS a_7195_65564# a_7126_65693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8588 a_5169_24643# a_5085_24759# a_5087_24643# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8589 a_17222_27247# a_16865_27511# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X859 a_13413_47375# a_11067_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X8590 VDD a_1586_36727# a_7295_43031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8591 a_49798_62194# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8592 a_2672_21807# a_1591_21807# a_2325_22049# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8593 a_6260_47919# a_5345_47919# a_5913_48161# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X8594 vcm_commonmode a_16362_57174# a_45478_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8595 VSS a_5547_36495# a_5731_37039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8596 VSS a_19245_39747# a_20839_41001# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X8597 vcm_commonmode a_16362_67214# a_28410_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8598 VDD a_12877_16911# a_19282_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8599 a_34342_22910# a_10515_23975# a_34834_22512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X86 VDD a_38077_29941# a_31084_30485# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X860 VDD a_2099_59861# a_2327_27247# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X8600 a_32426_65206# a_16746_65208# a_32334_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8601 a_37846_64524# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8602 a_32887_40767# a_32121_40741# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X8603 a_31330_20902# a_16362_20536# a_31422_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8604 a_39389_52271# a_39219_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8605 VDD a_12981_62313# a_41370_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8606 a_1644_74005# a_1591_64239# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8607 vcm_commonmode a_16362_59182# a_18370_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8608 a_6775_53877# a_22921_52245# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8609 VSS a_12355_15055# a_26706_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X861 VSS a_30375_51335# a_19576_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8610 a_22386_57174# a_16746_57176# a_22294_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8611 a_23694_18894# a_23736_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8612 a_33830_9460# a_32951_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8613 a_2215_36495# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8614 a_3357_67257# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8615 a_30722_60186# a_12981_59343# a_30326_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8616 a_30722_19898# a_12895_13967# a_30326_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8617 a_25204_44869# a_24331_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X8618 a_5903_13967# a_4812_13879# a_5814_13967# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X8619 VSS a_33155_40191# a_33101_40513# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X862 a_18674_10862# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8620 VSS a_6098_73095# a_6713_72765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8621 a_42374_70226# a_12516_7093# a_42866_70548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8622 a_3541_9593# a_1689_10396# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8623 VDD a_12985_19087# a_43378_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8624 a_38358_60186# a_12727_58255# a_38850_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8625 a_46390_68218# a_16362_68218# a_46482_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8626 VDD VSS a_27314_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8627 a_8305_16885# a_8087_17289# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8628 a_5903_13967# a_5959_13621# a_5731_13647# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X8629 a_41597_29967# a_41243_30080# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X863 vcm_commonmode a_16362_9492# a_31422_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8630 VDD a_37427_47893# a_17507_52047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X8631 a_41462_23548# a_16746_23546# a_41370_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8632 VSS a_7005_55223# a_6138_54599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8633 a_21261_47919# a_21095_47919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8634 a_40458_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8635 VDD a_5239_20693# a_3987_19623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X8636 VSS config_2_in[2] a_1591_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X8637 VSS a_18105_40157# a_17797_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8638 a_21737_49249# a_21519_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8639 a_28318_71230# a_12901_66665# a_28810_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X864 VSS a_30891_28309# a_26748_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8640 a_28810_20504# a_28756_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8641 VSS a_9219_71285# a_9150_71311# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=640000u l=150000u
X8642 VSS a_12727_67753# a_43774_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8643 a_40762_65206# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8644 a_28410_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8645 a_40858_17492# a_39673_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8646 a_11709_61217# a_11491_60975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8647 VSS a_12687_34191# a_12793_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8648 a_7865_46805# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8649 a_18770_12472# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X865 a_17927_31573# a_5831_39189# a_18145_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X8650 a_4885_71855# a_4719_71855# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8651 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8652 a_41370_9858# a_16362_9492# a_41462_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8653 a_12713_43011# a_18811_42405# a_19743_42359# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8654 a_10472_26159# a_10244_26159# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X8655 VDD a_12546_22351# a_22294_10862# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8656 vcm_commonmode VSS a_36442_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8657 a_2411_26133# a_2327_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8658 VDD a_6816_19355# a_7911_21379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8659 a_40458_70226# a_16746_70228# a_40366_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X866 a_27747_42359# a_26815_42405# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X8660 a_5533_17455# a_5363_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8661 a_20682_68218# a_12901_66959# a_20286_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8662 VSS a_12901_58799# a_46786_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8663 a_43774_56170# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8664 a_29322_12870# a_16362_12504# a_29414_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8665 a_17274_9858# a_16362_9492# a_17366_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8666 a_44874_16488# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8667 a_41370_13874# a_12727_15529# a_41862_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8668 a_8453_51727# a_7933_51433# a_8381_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8669 VSS a_12901_66959# a_29718_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X867 a_5695_10927# a_5345_10927# a_5600_10927# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8670 a_26706_66210# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8671 a_7162_59575# a_6559_59663# a_7376_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=0p ps=0u w=1e+06u l=150000u
X8672 a_18370_24552# VDD a_18278_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8673 VSS a_11067_13095# a_30722_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8674 a_48490_13508# a_16746_13506# a_48398_13874# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8675 vcm_commonmode a_16362_10496# a_45478_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8676 VDD a_29269_40741# a_30816_41605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X8677 a_27406_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8678 VSS a_20905_32143# a_22062_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8679 a_11115_59317# a_11521_58951# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X868 a_25702_11866# a_12985_16367# a_25306_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8680 a_5601_11471# a_4429_14191# a_5529_11471# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8681 a_5363_30503# a_15548_30761# a_20773_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X8682 VSS a_26397_51183# a_29847_48734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8683 vcm_commonmode a_16362_20536# a_28410_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8684 a_31330_65206# a_16362_65206# a_31422_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8685 a_34738_14878# a_12727_15529# a_34342_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8686 a_9355_32117# a_5346_33775# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X8687 a_23694_59182# a_12727_58255# a_23298_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8688 a_8576_28111# a_4248_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X8689 VSS a_12947_56817# a_20682_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X869 a_20649_36391# a_20957_36604# a_20623_36595# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X8690 a_17766_18496# a_17712_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8691 a_47790_55166# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8692 VSS a_10257_56377# a_10191_56445# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8693 VSS a_14926_31849# a_15925_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8694 VDD a_12727_13353# a_21290_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8695 a_17092_50959# a_14985_51701# a_16992_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X8696 VDD a_14912_27497# a_15599_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.165e+12p ps=6.33e+06u w=1e+06u l=150000u
X8697 a_35346_69222# a_12901_66959# a_35838_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8698 vcm_commonmode a_16362_12504# a_18370_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8699 a_5346_33775# a_4999_33781# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X87 a_24302_63198# a_16362_63198# a_24394_63198# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X870 VSS a_42188_43677# a_42283_42359# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X8700 a_13980_41605# a_13107_41317# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X8701 a_22386_10496# a_16746_10494# a_22294_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8702 a_28318_18894# a_16362_18528# a_28410_18528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8703 VDD a_4124_64391# a_4075_64239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8704 VSS a_33641_29967# a_39115_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X8705 a_48398_68218# a_12727_67753# a_48890_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8706 a_12579_35862# a_12549_35836# a_12507_35862# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X8707 a_1987_33402# a_1867_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8708 a_1815_12342# a_1633_12342# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X8709 a_33826_50075# a_33515_48576# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X871 a_2689_65103# a_1770_14441# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.053e+12p pd=1.104e+07u as=0p ps=0u w=650000u l=150000u M=4
X8710 a_47486_60186# a_16746_60188# a_47394_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8711 a_47486_19532# a_16746_19530# a_47394_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8712 a_22294_67214# a_16362_67214# a_22386_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8713 a_27710_58178# a_12901_58799# a_27314_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8714 a_11521_66567# a_12047_57685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8715 VSS VSS a_24698_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8716 a_26259_47491# a_25015_48437# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8717 VSS a_12683_51329# a_14092_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X8718 a_6927_71855# a_6913_72399# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X8719 a_38850_7452# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X872 a_38299_31055# a_36507_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X8720 a_34738_7850# a_33864_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8721 a_36442_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8722 VSS a_76082_40202# a_75824_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8723 a_19946_51157# a_2840_66103# a_21831_51183# VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u M=2
X8724 a_35458_28879# a_33839_28309# a_35345_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.55e+11p pd=5.31e+06u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X8725 VDD VDD a_48398_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8726 VSS VDD a_44778_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8727 a_25798_68540# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8728 a_32730_17890# a_12899_11471# a_32334_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8729 a_17774_27791# a_9529_28335# a_17691_27791# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X873 a_45386_70226# a_16362_70226# a_45478_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8730 a_21712_43781# a_20743_43493# a_21616_43781# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8731 a_9370_60975# a_7580_61751# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8732 a_12257_56623# a_11619_56615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8733 a_39758_23914# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8734 a_13643_28327# a_35815_31751# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8735 a_9234_32509# a_9135_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8736 VSS a_11067_21583# a_43774_21906# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8737 a_25702_9858# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8738 VDD a_19416_51017# a_19591_50943# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8739 a_46882_57496# a_43267_31055# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X874 VDD a_6444_16367# a_6619_16341# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8740 a_3449_54201# a_2840_53511# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8741 a_41766_72234# VDD a_41370_72234# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8742 VSS a_3016_60949# a_4340_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8743 a_12056_65327# a_10975_65327# a_11709_65569# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X8744 a_29814_67536# a_29760_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8745 a_26310_64202# a_11067_13095# a_26802_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8746 a_40233_27791# a_18979_30287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8747 a_3983_25321# a_3325_18543# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8748 a_30818_62516# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8749 VSS a_12727_15529# a_33734_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X875 a_46882_9460# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8750 a_13957_36121# a_12663_35431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X8751 a_29322_57174# a_16362_57174# a_29414_57174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8752 a_32887_42405# a_32121_42369# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X8753 a_21012_30761# a_21273_30485# a_21231_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X8754 VSS a_12877_16911# a_46786_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8755 a_20682_21906# a_12985_7663# a_20286_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8756 VSS a_4351_67279# a_23193_52245# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8757 a_10045_21379# a_6559_22671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8758 a_2107_71689# a_1757_71317# a_2012_71677# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8759 VDD a_10515_22671# a_23298_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X876 a_37750_64202# a_12355_65103# a_37354_64202# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8760 a_46390_7850# VSS a_46482_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8761 VSS a_10515_23975# a_29718_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8762 a_38754_70226# a_38557_32143# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8763 a_37446_68218# a_16746_68220# a_37354_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8764 a_36350_23914# a_16362_23548# a_36442_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8765 a_36600_49159# a_4351_67279# a_36831_49257# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8766 a_4682_10749# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8767 a_23694_12870# a_10055_58791# a_23298_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8768 a_35742_63198# a_15439_49525# a_35346_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8769 a_1803_20719# a_1626_20719# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X877 a_33734_59182# a_25787_28327# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8770 vcm_commonmode a_16362_23548# a_30418_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8771 VDD a_2021_17973# a_27359_43985# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8772 a_12671_36694# a_12713_36483# a_12671_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8773 a_19684_35077# a_18811_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X8774 a_12219_47158# a_7571_26151# a_11760_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8775 a_43378_71230# a_16362_71230# a_43470_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8776 a_48794_62194# a_12981_62313# a_48398_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8777 a_8271_74953# a_7921_74581# a_8176_74941# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X8778 VSS a_10515_63143# a_12723_14191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X8779 VSS a_12895_13967# a_45782_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X878 a_35838_72556# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8780 a_46482_7484# VDD a_46390_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8781 vcm_commonmode a_16362_61190# a_19374_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8782 a_32730_68218# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8783 a_23390_18528# a_16746_18526# a_23298_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8784 VDD a_11067_21583# a_33338_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8785 a_12831_38543# a_12801_38517# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8786 VDD a_12901_58799# a_27314_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8787 vcm_commonmode a_16362_15516# a_20378_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8788 a_27710_11866# a_12985_16367# a_27314_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8789 a_43319_31029# a_43678_31029# a_43455_31055# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X879 VDD a_12985_7663# a_35346_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8790 VSS a_6607_39991# a_6559_39759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8791 a_15074_50871# a_14983_51157# a_15288_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.7e+11p pd=2.94e+06u as=0p ps=0u w=1e+06u l=150000u
X8792 VSS a_33694_30761# a_33741_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X8793 a_2835_62215# a_3108_62043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X8794 VSS a_10667_60735# a_10601_60809# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8795 a_20378_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8796 vcm_commonmode a_16362_9492# a_27406_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8797 a_47394_70226# a_16362_70226# a_47486_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8798 a_46786_14878# a_43175_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8799 a_15080_32143# a_14354_32117# a_8491_41383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.37e+12p ps=1.274e+07u w=1e+06u l=150000u M=4
X88 a_45782_68218# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X880 VSS a_2012_33927# a_2093_28918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8800 a_7581_74031# a_6098_73095# a_7499_74031# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8801 VDD a_8197_31599# a_11644_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X8802 a_4298_58951# a_7815_49855# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8803 a_37846_72556# a_36613_48169# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8804 a_5043_20214# a_4792_20443# a_4584_20407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8805 VDD a_12985_7663# a_37354_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8806 vcm_commonmode a_16362_14512# a_24394_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8807 VDD a_12901_66665# a_41370_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8808 a_33338_16886# a_12899_11471# a_33830_16488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8809 a_34434_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X881 vcm_commonmode a_16362_14512# a_22386_14512# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8810 a_4139_23145# a_3325_18543# a_4067_23145# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8811 a_32795_29967# a_32544_30083# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X8812 a_37354_62194# a_16362_62194# a_37446_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8813 a_20286_19898# a_11067_67279# a_20778_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8814 a_31422_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8815 a_41462_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8816 VDD a_12889_35537# a_12831_35645# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X8817 a_2417_52513# a_2199_52271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8818 a_4127_50069# a_5135_50069# a_5081_50095# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8819 a_24394_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X882 a_31330_16886# a_12899_11471# a_31822_16488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8820 a_12407_54965# a_12755_53030# a_12689_55311# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X8821 VDD a_7865_46805# a_7895_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8822 VSS a_2163_73085# a_2124_73211# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8823 vcm_commonmode a_16362_66210# a_49494_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8824 a_4906_60431# a_4187_60673# a_4343_60405# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X8825 a_1683_5059# a_1761_2767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8826 a_1881_54447# a_1846_54699# a_1643_54421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8827 a_38450_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8828 a_1915_20394# a_2007_20149# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X8829 VSS a_8753_31055# a_14097_31375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X883 a_16228_28335# a_15599_28585# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X8830 a_12473_37429# a_30991_35307# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X8831 VSS a_12983_63151# a_35742_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8832 a_9326_49334# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X8833 VSS a_2411_26133# a_2369_36861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8834 a_27406_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8835 a_43470_56170# a_16746_56172# a_43378_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8836 a_44778_17890# a_42718_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8837 a_37446_21540# a_16746_21538# a_37354_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8838 a_6905_63151# a_6831_63303# a_6559_63401# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.38e+11p ps=3.64e+06u w=650000u l=150000u
X8839 a_10590_21263# a_10151_21379# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X884 VDD a_13390_29575# a_2787_30503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.62e+12p ps=1.524e+07u w=1e+06u l=150000u M=4
X8840 a_26402_66210# a_16746_66212# a_26310_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8841 a_7577_60137# a_6467_55527# a_7162_60039# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X8842 a_5345_74031# a_5179_74031# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8843 a_25306_21906# a_16362_21540# a_25398_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8844 a_28410_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8845 VDD a_15439_49525# a_35346_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8846 a_2203_9839# a_1757_9839# a_2107_9839# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X8847 VDD a_12899_10927# a_39362_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8848 a_15775_36965# a_13557_37999# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X8849 VDD a_11067_13095# a_12712_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X885 a_38450_65206# a_16746_65208# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8850 a_30975_28023# a_30052_32117# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8851 VDD a_9707_51325# a_9668_51451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8852 VSS a_12899_10927# a_21686_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8853 a_32730_21906# a_32772_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8854 a_29322_20902# a_16362_20536# a_29414_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8855 VSS a_9637_30511# a_10280_31171# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8856 a_12139_18517# a_11964_18543# a_12318_18543# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8857 a_5318_18909# a_4241_18543# a_5156_18543# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8858 a_2464_73309# a_2250_73309# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8859 a_44474_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X886 a_35346_62194# a_16362_62194# a_35438_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8860 a_46786_55166# VSS a_46390_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8861 a_6909_51183# a_5909_51433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8862 VDD a_11130_22869# a_11067_47695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X8863 VDD a_6743_23555# a_7187_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8864 VSS VDD a_30722_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8865 a_41325_30333# a_35815_31751# a_41243_30080# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8866 a_29718_65206# a_10975_66407# a_29322_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8867 a_2369_18543# a_2325_18785# a_2203_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X8868 VDD a_12516_7093# a_34342_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8869 a_22690_13874# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X887 a_25307_51549# a_24683_51183# a_25199_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X8870 a_13107_41317# a_12341_41281# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X8871 VSS a_5291_56765# a_5252_56891# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8872 a_9150_71311# a_9063_71553# a_8746_71443# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X8873 a_23390_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8874 a_34434_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8875 a_3705_37557# a_3487_37961# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X8876 a_47790_63198# a_43362_28879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8877 a_17366_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8878 vcm_commonmode a_16362_58178# a_43470_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8879 a_19678_57174# a_10515_22671# a_19282_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X888 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X8880 a_19967_41781# a_52778_39936# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8881 a_34738_66210# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8882 vcm_commonmode a_16362_68218# a_26402_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8883 a_35838_65528# a_34251_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8884 VDD a_40743_31287# a_31659_31751# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8885 a_45386_22910# a_10515_23975# a_45878_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8886 a_3763_10761# a_3413_10389# a_3668_10749# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X8887 VDD a_1586_36727# a_4259_32687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8888 a_2125_68053# a_1959_68053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8889 a_11759_59575# a_11521_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X889 VSS a_10747_68565# a_8958_65961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8890 a_38450_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8891 a_35346_55166# VSS a_35438_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8892 a_21479_42405# a_19596_42919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X8893 a_2163_59585# a_3295_54421# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X8894 a_6809_27907# a_6773_27805# a_6737_27907# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8895 VDD a_2283_15797# a_2873_13879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8896 VSS a_12981_62313# a_24698_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8897 a_21686_60186# a_17507_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8898 a_10325_67503# a_9135_67503# a_10216_67503# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X8899 a_20378_58178# a_16746_58180# a_20286_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X89 a_36442_18528# a_16746_18526# a_36350_18894# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X890 VSS a_9828_56311# a_9599_57141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8900 a_21686_19898# a_9135_27239# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X8901 a_34434_71230# a_16746_71232# a_34342_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8902 a_8176_74941# a_8059_74746# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8903 a_25417_51425# a_25199_51183# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X8904 a_38850_17492# a_37919_28111# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8905 a_35346_14878# a_12877_14441# a_35838_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8906 VSS a_12985_7663# a_35742_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X8907 a_38754_23914# a_10515_23975# a_38358_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8908 a_9326_49007# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X8909 VDD a_12877_14441# a_42374_15882# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X891 VDD a_11067_67279# a_48398_20902# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8910 a_16707_40183# a_16744_40517# VSS VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X8911 a_15683_39141# a_13097_39631# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X8912 a_18278_24918# a_18007_27441# a_18770_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8913 a_22448_38341# a_21479_38053# a_22411_38007# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X8914 a_22786_22512# a_12341_3311# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8915 a_49402_21906# a_11067_21583# a_49894_21508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8916 a_49402_17890# a_16362_17524# a_49494_17524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8917 VDD a_2847_15039# a_2834_14735# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8918 VDD a_19877_52245# a_20535_51727# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X8919 a_8123_34639# a_4685_37583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X892 VSS a_40139_32143# a_35815_31751# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u M=4
X8920 a_12885_43222# a_12713_43011# a_12671_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X8921 a_38450_70226# a_16746_70228# a_38358_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8922 a_4169_67753# a_3024_67191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8923 a_29915_41959# a_26433_39631# a_30089_41835# VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8924 VSS a_4503_10687# a_4437_10761# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X8925 a_39362_13874# a_12727_15529# a_39854_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8926 a_43870_11468# a_40491_27247# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8927 VSS a_11067_13095# a_28714_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8928 a_36797_27497# a_22291_29415# a_36725_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8929 VDD a_8325_18517# a_8355_18870# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X893 a_20713_39105# a_21387_38591# a_22319_38825# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X8930 a_33830_68540# a_25787_28327# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8931 a_26310_72234# VDD a_26802_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8932 a_26802_21508# a_26748_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8933 a_26402_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8934 a_30818_70548# a_25971_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8935 a_23298_14878# a_16362_14512# a_23390_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8936 VSS a_2775_46025# a_32972_52047# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u M=4
X8937 a_29322_65206# a_16362_65206# a_29414_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8938 VSS a_12215_31573# a_14747_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X8939 a_3425_42313# a_2235_41941# a_3316_42313# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X894 a_18278_72234# VSS a_18370_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8940 VSS a_2411_26133# a_2369_26159# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8941 vcm_commonmode a_16362_17524# a_38450_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8942 a_30326_60186# a_16362_60186# a_30418_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8943 a_52778_39198# a_52590_39198# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X8944 VSS a_12947_56817# a_18674_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8945 a_6786_37557# a_6372_38279# a_7289_38127# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X8946 a_42466_15516# a_16746_15514# a_42374_15882# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8947 VDD a_27560_34337# a_29205_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X8948 a_13275_32463# a_8461_32937# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X8949 a_35307_49871# a_34145_49007# a_35224_49871# VSS sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X895 a_48398_61190# a_16362_61190# a_48490_61190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8950 VDD a_12985_16367# a_20286_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8951 a_45782_9858# a_12985_19087# a_45386_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8952 VDD VSS a_19282_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8953 a_22164_51157# a_22015_51840# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8954 a_10509_72943# a_9353_72399# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8955 a_77568_39738# a_77664_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8956 a_34342_64202# a_11067_13095# a_34834_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8957 a_29814_12472# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8958 a_12231_60949# a_12056_60975# a_12410_60975# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X8959 a_41766_57174# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X896 a_22386_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8960 a_27314_13874# a_16362_13508# a_27406_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8961 VSS a_10590_21263# a_9955_20969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X8962 a_10964_25615# a_10521_25731# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X8963 a_47394_63198# a_12981_62313# a_47886_63520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X8964 VSS a_30052_32117# a_41405_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X8965 a_5490_41365# a_5963_36585# a_7650_35951# VSS sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=0p ps=0u w=650000u l=150000u M=4
X8966 a_31726_68218# a_12901_66959# a_31330_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8967 a_46482_14512# a_16746_14510# a_46390_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8968 vcm_commonmode a_16362_11500# a_43470_11500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8969 a_19678_10862# a_12546_22351# a_19282_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X897 vcm_commonmode a_16362_67214# a_34434_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8970 a_27429_35301# a_27183_34789# a_28056_35077# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8971 vcm_commonmode a_16362_56170# a_32426_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8972 a_42866_19500# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8973 a_29414_24552# VDD a_29322_24918# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8974 vcm_commonmode a_16362_21540# a_26402_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8975 a_8061_58575# a_3295_62083# a_7963_58255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X8976 a_8468_48841# a_7553_48469# a_8121_48437# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X8977 VDD a_2511_60431# a_1923_59583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=4
X8978 VSS a_2473_34293# a_3805_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8979 a_21012_30761# a_20911_31055# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.85e+11p pd=5.37e+06u as=0p ps=0u w=1e+06u l=150000u
X898 a_3339_32463# a_17787_47349# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X8980 a_28441_36389# a_28195_35327# a_29068_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8981 a_19596_40743# a_18627_40767# a_19500_40743# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X8982 VDD a_12983_63151# a_27314_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X8983 a_5438_69679# a_5091_69685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X8984 a_24794_63520# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8985 a_5531_22895# a_5087_23145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X8986 VDD a_2847_49855# a_2834_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8987 a_19374_16520# a_16746_16518# a_19282_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8988 VSS a_11067_23759# a_16362_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u M=2
X8989 a_4151_28879# a_3707_28995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X899 a_32318_48695# a_6831_63303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X8990 a_13620_43047# a_13005_43983# a_13762_42895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X8991 a_7553_48469# a_7387_48469# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X8992 VSS a_10317_55223# a_9695_54965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8993 a_20378_11500# a_16746_11498# a_20286_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X8994 a_27600_36165# a_26631_35877# a_27563_35831# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X8995 a_42866_8456# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8996 a_46390_69222# a_12901_66959# a_46882_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8997 a_5159_43933# a_4535_43567# a_5051_43567# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X8998 VSS a_11760_46983# a_10407_47607# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X8999 a_18674_58178# a_14287_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9 a_27214_28335# a_2787_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.2285e+12p pd=1.288e+07u as=0p ps=0u w=650000u l=150000u M=4
X90 VSS a_24331_38591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X900 VSS a_8509_47673# a_8443_47741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9000 VDD a_5079_35639# a_5153_34025# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X9001 a_20286_68218# a_16362_68218# a_20378_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9002 a_18770_8456# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9003 a_2203_18543# a_1757_18543# a_2107_18543# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9004 VSS a_28757_27247# a_41596_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9005 a_28810_62516# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9006 a_19780_41605# a_18811_41317# a_19743_41271# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9007 a_34434_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9008 a_33338_67214# a_16362_67214# a_33430_67214# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9009 a_10045_29967# a_8273_42479# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X901 a_6614_21237# a_2339_38129# VSS VSS sky130_fd_pr__nfet_01v8 ad=4.225e+11p pd=3.9e+06u as=0p ps=0u w=650000u l=150000u
X9010 a_21519_49007# a_21169_49007# a_21424_49007# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X9011 VDD a_30412_34337# a_29513_34428# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X9012 VDD a_12947_8725# a_28318_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9013 VSS a_12985_19087# a_24698_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9014 a_47486_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9015 a_1644_77813# a_1823_77821# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9016 a_23298_59182# a_16362_59182# a_23390_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9017 a_15957_39655# a_16265_39868# a_15931_39859# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X9018 a_37750_24918# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9019 a_43774_17890# a_12899_11471# a_43378_17890# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X902 a_25263_34473# a_24331_34239# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9020 VSS a_5039_42167# a_14634_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9021 a_26767_50095# a_26321_50095# a_26671_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X9022 VDD a_1923_54591# a_4311_52245# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9023 a_41370_55166# VSS a_41862_55488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9024 VSS a_19531_49007# a_19715_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9025 VSS a_2451_72373# a_3275_73658# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9026 a_22178_30761# a_14646_29423# a_22105_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=9.03e+10p ps=1.27e+06u w=420000u l=150000u
X9027 VDD a_33856_40743# a_33760_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9028 VSS a_13445_51335# a_12755_51562# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9029 vcm_commonmode a_16362_61190# a_40458_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X903 VDD a_23911_35823# a_24017_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9030 a_27314_58178# a_16362_58178# a_27406_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9031 VSS a_5535_18012# a_8753_19319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9032 a_1863_42729# a_1778_42631# a_1645_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9033 vcm_commonmode a_16362_71230# a_23390_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9034 a_47790_16886# a_12727_13353# a_47394_16886# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9035 a_2127_4943# a_1683_5059# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X9036 VDD a_2325_22049# a_2215_22173# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9037 a_7563_46261# a_7407_46529# a_7708_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X9038 VSS a_12727_15529# a_44778_13874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9039 a_41766_10862# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X904 vcm_commonmode a_16362_66210# a_47486_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9040 VDD a_1586_40455# a_1591_44655# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9041 VDD a_12947_71576# a_35346_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9042 a_27314_17890# a_12899_10927# a_27806_17492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9043 a_26310_8854# a_16362_8488# a_26402_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9044 VSS a_12947_23413# a_27710_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9045 a_31822_15484# a_31768_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9046 a_21290_7850# VDD a_21782_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9047 a_31726_21906# a_12985_7663# a_31330_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9048 VSS a_38171_34191# a_38277_34191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9049 VSS a_20359_29199# a_37195_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X905 VDD a_10055_58791# a_38358_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9050 vcm_commonmode a_16362_8488# a_40458_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9051 vcm_commonmode a_16362_60186# a_44474_60186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9052 a_21169_49007# a_21003_49007# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9053 a_18370_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9054 vcm_commonmode a_16362_19532# a_44474_19532# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9055 a_48890_59504# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9056 VSS a_12727_13353# a_17670_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9057 vcm_commonmode a_16362_70226# a_27406_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9058 a_21686_13874# a_12877_16911# a_21290_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9059 a_4956_43567# a_4839_43780# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X906 a_30105_32463# a_18979_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X9060 a_17763_43413# a_17939_43745# a_17891_43805# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9061 VDD a_19311_35823# a_19417_35823# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9062 a_17843_48981# a_17039_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9063 VDD a_6831_63303# a_29220_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.5e+11p ps=5.7e+06u w=1e+06u l=150000u
X9064 a_41370_72234# VSS a_41462_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9065 a_46786_63198# a_15439_49525# a_46390_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9066 a_32334_11866# a_10055_58791# a_32826_11468# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9067 VSS a_7479_54439# a_8219_54447# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9068 a_12901_66665# a_11067_67279# a_12901_66415# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9069 a_22294_68218# a_12727_67753# a_22786_68540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X907 a_36442_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9070 a_26402_8488# a_16746_8486# a_26310_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9071 a_33734_66210# a_12983_63151# a_33338_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9072 vcm_commonmode a_16362_62194# a_17366_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9073 a_18278_58178# a_10515_22671# a_18770_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9074 a_21382_60186# a_16746_60188# a_21290_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9075 a_21382_19532# a_16746_19530# a_21290_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9076 VDD a_12727_58255# a_25306_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9077 VDD a_7624_68021# a_7571_68047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9078 a_18703_29199# a_33694_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X9079 a_18674_11866# a_8491_27023# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X908 a_49402_24918# VSS a_49494_24552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9080 a_8853_61839# a_3295_62083# a_8635_61751# VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9081 VSS a_5749_18297# a_5683_18365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9082 VSS a_18445_46805# a_18379_46831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9083 VDD a_11067_21583# a_44382_22910# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9084 vcm_commonmode a_16362_15516# a_31422_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9085 a_29364_50959# a_6831_63303# a_28789_50613# VSS sky130_fd_pr__nfet_01v8 ad=1.6575e+11p pd=1.81e+06u as=0p ps=0u w=650000u l=150000u
X9086 a_9125_24527# a_8569_25071# a_9043_24527# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9087 VDD a_26523_29199# a_33363_30305# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9088 a_37750_65206# a_10975_66407# a_37354_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9089 VDD a_12727_15529# a_34342_14878# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X909 VDD a_33641_29967# a_40691_30511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.646e+11p ps=2.94e+06u w=420000u l=150000u
X9090 a_9759_67869# a_9135_67503# a_9651_67503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X9091 VSS a_1586_45431# a_1591_45205# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9092 a_35346_63198# a_16362_63198# a_35438_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9093 VDD a_1586_9991# a_1591_14741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9094 a_18856_41831# a_17983_41855# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9095 VDD a_12985_7663# a_48398_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9096 a_12707_26159# a_12263_26409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X9097 a_45478_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9098 a_31114_48169# a_6831_63303# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9099 vcm_commonmode a_16362_68218# a_34434_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 a_3949_41935# a_3491_42239# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=4
X910 a_36579_41271# a_35932_41953# VSS VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u M=2
X9100 a_48398_62194# a_16362_62194# a_48490_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9101 a_31330_19898# a_11067_67279# a_31822_19500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9102 a_9184_49159# a_4298_58951# a_9326_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9103 a_9326_13430# a_1929_12131# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9104 a_4761_45743# a_4717_45985# a_4595_45743# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X9105 VDD a_12877_16911# a_38358_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9106 VDD a_2223_28617# a_2899_27023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9107 a_13081_29199# a_11719_28023# a_12935_31287# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9108 VSS a_18979_30287# a_35357_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X9109 vcm_commonmode a_16362_67214# a_47486_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X911 VSS a_2686_70223# a_4073_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X9110 a_35838_10464# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9111 a_7802_42845# a_6725_42479# a_7640_42479# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9112 VSS a_2589_62839# a_2099_64757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9113 a_8056_13967# a_7841_12167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9114 a_25961_48169# a_25015_48437# a_25879_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.1285e+11p ps=5.04e+06u w=1e+06u l=150000u
X9115 VSS a_10575_62911# a_10509_62985# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X9116 a_49494_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9117 a_25398_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9118 vcm_commonmode a_16362_59182# a_37446_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9119 a_41462_57174# a_16746_57176# a_41370_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X912 a_49494_12504# a_16746_12502# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9120 a_2872_44111# a_2695_44119# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9121 a_42770_18894# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9122 VDD a_5691_36727# a_6930_37583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9123 VSS a_33360_51701# a_32582_51701# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u M=4
X9124 VSS VDD a_28714_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9125 a_24394_67214# a_16746_67216# a_24302_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9126 vcm_commonmode a_16362_64202# a_21382_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9127 a_6177_61127# a_6382_61127# a_6340_61225# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9128 a_26350_28335# a_2787_30503# a_26350_28585# VSS sky130_fd_pr__nfet_01v8 ad=8.775e+11p pd=9.2e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9129 a_10751_59575# a_2840_66103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X913 a_2150_43401# a_1757_43029# a_2040_43401# VSS sky130_fd_pr__nfet_01v8 ad=1.341e+11p pd=1.5e+06u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X9130 a_23298_22910# a_16362_22544# a_23390_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9131 a_2834_45199# a_1757_45205# a_2672_45577# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9132 VDD a_12355_65103# a_33338_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9133 a_25306_9858# a_12546_22351# a_25798_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9134 VDD a_15439_49525# a_46390_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9135 a_22690_62194# a_12981_62313# a_22294_62194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9136 a_5235_71855# a_4885_71855# a_5140_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X9137 a_1642_22583# a_1738_22325# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9138 a_11711_32463# a_10515_32143# a_11711_32143# VSS sky130_fd_pr__nfet_01v8 ad=5.3625e+11p pd=5.55e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9139 VDD a_14985_51701# a_15489_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X914 a_43227_28309# a_18703_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X9140 VSS a_20957_36604# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X9141 VSS a_12993_50345# a_13445_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9142 a_34342_72234# VDD a_34834_72556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9143 VSS a_12899_10927# a_32730_17890# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9144 VSS a_15812_31029# a_7598_36103# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X9145 a_30991_29397# a_31117_28879# a_31422_29423# VSS sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X9146 a_5784_16367# a_5533_17455# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9147 VDD a_31096_38341# a_31000_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9148 a_34834_60508# a_34780_56398# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9149 a_47394_71230# a_12901_66665# a_47886_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X915 a_7050_53333# a_17843_48981# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9150 a_42466_68218# a_16746_68220# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9151 a_4584_20407# a_4792_20443# a_4726_20541# VSS sky130_fd_pr__nfet_01v8 ad=1.995e+11p pd=1.79e+06u as=0p ps=0u w=420000u l=150000u
X9152 a_77086_40693# a_75794_38962# a_76971_38925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u M=2
X9153 a_13183_52047# a_20267_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9154 a_19678_60186# a_19720_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9155 a_18370_58178# a_16746_58180# a_18278_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9156 a_19678_19898# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9157 VDD a_23784_42583# a_23597_42325# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9158 a_20682_14878# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9159 VDD a_2292_43291# a_7708_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X916 a_25398_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9160 a_23577_50095# a_23535_50247# a_23487_50095# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.95e+11p ps=1.9e+06u w=650000u l=150000u
X9161 a_33734_13874# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9162 VSS a_1586_66567# a_3983_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9163 a_24794_71552# a_18151_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9164 a_45478_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9165 VSS a_3983_70767# a_4060_70223# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9166 a_47790_8854# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9167 a_24302_61190# a_16362_61190# a_24394_61190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9168 a_28799_29423# a_23192_27791# a_28703_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9169 VSS a_12901_66959# a_48794_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X917 a_49798_69222# a_12516_7093# a_49402_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9170 a_45782_66210# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9171 vcm_commonmode a_16362_21540# a_34434_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9172 a_43378_23914# a_12947_23413# a_43870_23516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9173 a_43378_19898# a_16362_19532# a_43470_19532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9174 VSS a_2787_30503# a_24632_32259# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9175 a_9326_13103# a_1929_12131# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9176 a_77451_38925# a_76971_38925# sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9177 vcm_commonmode a_16362_20536# a_47486_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9178 VDD a_36507_31573# a_35299_32375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9179 a_28810_70548# a_28756_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X918 a_77285_39738# a_77381_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9180 a_49494_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9181 a_46390_55166# VSS a_46482_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9182 a_42770_59182# a_12727_58255# a_42374_59182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9183 VDD a_12473_42869# a_12885_43222# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9184 a_37459_51183# a_4351_67279# a_37287_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9185 a_36842_18496# a_36629_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9186 a_36746_24918# VSS a_36350_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9187 a_34698_31055# a_33641_29967# a_34395_31287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X9188 a_45478_71230# a_16746_71232# a_45386_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9189 VDD a_12727_13353# a_40366_16886# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X919 VSS a_15548_30761# a_22062_31287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X9190 a_25702_69222# a_12516_7093# a_25306_69222# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9191 VSS a_10975_66407# a_22690_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9192 a_49798_65206# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9193 vcm_commonmode a_16362_12504# a_37446_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9194 a_49894_17492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9195 a_46390_14878# a_12877_14441# a_46882_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9196 a_49798_23914# a_10515_23975# a_49402_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9197 a_20778_23516# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9198 a_7493_12015# a_7841_12167# VSS VSS sky130_fd_pr__nfet_01v8 ad=6.24e+11p pd=5.82e+06u as=0p ps=0u w=650000u l=150000u
X9199 a_20378_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X92 a_2672_45577# a_1757_45205# a_2325_45173# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X920 a_41462_56170# a_16746_56172# a_41370_56170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9200 a_12885_36694# a_12713_36483# a_12671_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X9201 VSS a_14983_51157# a_17092_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9202 a_41462_10496# a_16746_10494# a_41370_10862# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9203 a_47394_18894# a_16362_18528# a_47486_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9204 a_9063_71553# a_9314_69367# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9205 a_32970_31145# a_39272_31573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9206 VSS a_15959_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X9207 a_24394_20536# a_16746_20534# a_24302_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9208 a_2886_47158# a_2656_45895# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9209 a_23626_31573# a_14926_31849# a_23849_30511# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X921 a_42770_17890# a_41967_31375# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9210 a_39758_57174# a_39389_52271# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9211 VDD a_28841_29575# a_41232_28879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9212 a_39758_15882# a_12877_14441# a_39362_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9213 VSS VSS a_43774_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9214 a_25129_48463# a_25015_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9215 a_49494_70226# a_16746_70228# a_49402_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9216 VSS a_12355_65103# a_26706_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9217 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9218 a_20378_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9219 a_7381_35407# a_5963_36585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X922 a_35438_21540# a_16746_21538# a_35346_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9220 VDD a_12899_11471# a_26310_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9221 a_4174_49334# a_2606_41079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9222 a_24394_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9223 a_21290_15882# a_16362_15516# a_21382_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9224 VDD a_2375_29588# a_1895_30138# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X9225 a_44874_68540# a_39299_48783# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9226 a_39454_62194# a_16746_62196# a_39362_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9227 vcm_commonmode a_16362_18528# a_36442_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9228 a_8397_35407# a_6372_38279# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9229 a_40458_16520# a_16746_16518# a_40366_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X923 a_8123_28879# a_6162_28487# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=9.65e+11p pd=7.93e+06u as=0p ps=0u w=1e+06u l=150000u
X9230 a_4328_10761# a_3247_10389# a_3981_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9231 a_20682_55166# VSS a_20286_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9232 a_2451_72373# a_4119_70741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u M=2
X9233 a_7803_11703# a_7203_10383# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9234 VSS a_12947_56817# a_29718_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9235 vcm_commonmode a_16362_8488# a_49494_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9236 a_75794_40594# a_75628_40594# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9237 VDD a_11115_59317# a_11054_59343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X9238 a_31422_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9239 a_18370_11500# a_16746_11498# a_18278_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X924 VSS a_12901_66665# a_28714_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9240 a_27806_13476# a_27752_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9241 a_22097_30287# a_14646_29423# a_20946_30669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9242 VDD a_12985_16367# a_31330_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9243 a_39029_29673# a_32823_29397# a_38436_29941# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9244 VDD a_12895_13967# a_17274_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9245 VDD a_12901_66959# a_21290_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9246 a_48890_67536# a_42985_46831# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9247 a_45386_64202# a_11067_13095# a_45878_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9248 VSS a_26319_41781# a_13576_42589# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9249 a_36442_8488# a_16746_8486# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X925 VDD a_6883_37019# a_7061_34319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9250 VDD a_76648_39738# a_76461_39480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9251 a_16080_28111# a_14273_27791# a_16008_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X9252 a_4864_62581# a_2689_65103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9253 a_12404_34191# a_12227_34191# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9254 a_10679_74397# a_10055_74031# a_10571_74031# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X9255 VSS a_3143_22364# a_4083_22351# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9256 a_2981_28111# a_2473_34293# a_2899_28111# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9257 a_2307_31965# a_1683_31599# a_2199_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X9258 VSS a_5504_37815# a_5449_37191# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9259 vcm_commonmode a_16362_57174# a_30418_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X926 a_22352_44869# a_21479_44581# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X9260 a_10570_25625# a_9669_26703# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9261 a_35346_56170# a_12947_56817# a_35838_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9262 VDD VDD a_41370_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9263 VDD a_10515_22671# a_42374_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9264 VSS a_10515_23975# a_48794_22910# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9265 a_18278_66210# a_10975_66407# a_18770_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9266 a_15097_51183# a_14983_51157# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9267 VSS a_1923_54591# a_5009_56623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9268 VDD a_6608_19319# a_5135_19061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9269 VDD a_12727_67753# a_25306_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X927 a_24394_66210# a_16746_66212# a_24302_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9270 a_22786_64524# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9271 VDD VDD a_17274_7850# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9272 VDD a_29913_43457# a_30356_42919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9273 VSS a_49750_39288# a_51714_39886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X9274 a_25204_40743# a_24331_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X9275 a_18627_40767# a_15397_39631# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X9276 a_19026_31375# a_18162_31055# a_12447_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9277 a_42770_12870# a_10055_58791# a_42374_12870# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9278 a_23694_7850# VDD a_23298_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9279 a_39362_55166# VSS a_39854_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X928 VDD a_1586_36727# a_1683_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9280 a_25702_22910# a_11067_21583# a_25306_22910# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9281 VSS a_12516_7093# a_34738_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9282 VDD a_13669_37429# a_13613_37782# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9283 a_24931_42657# a_12473_42869# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9284 a_5915_35943# a_20027_27221# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X9285 a_11711_67325# a_11521_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9286 VDD a_5767_31573# a_5713_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9287 a_23298_60186# a_12727_58255# a_23790_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9288 VDD a_4625_50613# a_4515_50639# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9289 a_31330_68218# a_16362_68218# a_31422_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X929 a_2325_71285# a_2107_71689# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9290 a_16746_17522# a_16510_8760# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u M=2
X9291 VDD a_13576_40413# a_17797_40517# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9292 a_7624_68021# a_5024_67885# a_7844_68367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9293 VDD a_3339_30503# a_27132_28585# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u M=4
X9294 a_39758_10862# a_39223_32463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9295 a_45478_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9296 a_16762_55488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9297 VDD a_6099_23983# a_5085_23047# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9298 VSS a_12981_59343# a_37750_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9299 a_4065_30761# a_3417_33231# a_3983_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X93 a_31330_11866# a_16362_11500# a_31422_11500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X930 a_39247_38007# a_38315_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9300 a_3070_22390# a_2012_33927# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X9301 VDD a_4495_35925# a_7009_33231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9302 a_4174_49007# a_2606_41079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9303 a_41766_18894# a_12899_10927# a_41370_18894# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9304 a_9361_28335# a_7281_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9305 a_2250_73309# a_2163_73085# a_1846_73195# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9306 a_25398_7484# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9307 a_2325_12533# a_2107_12937# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X9308 a_14361_29967# a_14013_30083# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9309 VDD a_21879_30663# a_21057_30669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X931 a_26402_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9310 a_39503_43957# a_39742_44527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9311 a_2191_68565# a_2847_44629# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9312 a_39362_72234# VSS a_39454_72234# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9313 a_37446_55166# VDD a_37354_55166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9314 a_38754_16886# a_37919_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9315 VSS a_4812_13879# a_5411_12791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9316 a_20914_49551# a_20195_49793# a_20351_49525# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X9317 vcm_commonmode VSS a_21382_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9318 a_43470_70226# a_16746_70228# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9319 VSS a_12877_14441# a_42770_14878# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X932 a_23298_21906# a_16362_21540# a_23390_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9320 a_12579_36189# a_12325_35862# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9321 a_36350_10862# a_16362_10496# a_36442_10496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9322 a_11978_29967# a_8485_29673# a_11886_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X9323 VSS a_12901_58799# a_31726_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9324 VDD VDD a_33338_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9325 a_25306_18894# a_12895_13967# a_25798_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9326 VSS VSS a_25702_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9327 VSS a_7162_60039# a_5749_60039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9328 a_33430_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9329 VDD config_1_in[5] a_1591_16367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X933 VDD a_15439_49525# a_33338_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9330 vcm_commonmode a_16362_15516# a_29414_15516# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9331 VDD a_12947_71576# a_46390_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9332 vcm_commonmode a_16362_9492# a_20378_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9333 vcm_commonmode a_16362_10496# a_30418_10496# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9334 a_16362_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9335 a_18674_60186# a_12981_59343# a_18278_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9336 VDD a_8652_17289# a_8827_17215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9337 a_18674_19898# a_12895_13967# a_18278_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9338 VSS a_9307_30663# a_10870_31599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X9339 a_46482_61190# a_16746_61192# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X934 VDD a_12901_66665# a_29322_70226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9340 VDD a_75199_38962# a_75628_38962# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9341 VDD a_1761_47919# a_28099_42895# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9342 a_29119_42359# a_29513_42333# a_28717_42917# VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=2.4e+11p ps=2.2e+06u w=800000u l=150000u
X9343 VDD a_8836_74953# a_9011_74879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9344 a_30418_9492# a_16746_9490# a_30326_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9345 VDD a_4219_34551# a_3187_34293# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X9346 a_29414_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9347 a_2380_68413# a_2263_68218# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9348 a_32795_41855# a_32029_41829# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X9349 a_12815_19319# a_12672_18115# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X935 a_7461_27247# a_7113_27253# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9350 VSS a_7097_67655# a_5160_68315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9351 a_20286_69222# a_12901_66959# a_20778_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9352 a_44382_21906# a_16362_21540# a_44474_21540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9353 VDD a_12985_19087# a_45386_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9354 a_29322_19898# a_11067_67279# a_29814_19500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9355 a_30311_40229# a_29545_40193# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X9356 a_33338_68218# a_12727_67753# a_33830_68540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9357 a_44778_66210# a_12983_63151# a_44382_66210# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9358 vcm_commonmode a_16362_62194# a_28410_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9359 a_2012_40303# a_1895_40516# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X936 VSS a_1761_52815# a_12559_44527# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9360 a_32426_60186# a_16746_60188# a_32334_60186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9361 a_32426_19532# a_16746_19530# a_32334_19898# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9362 VSS a_13669_37429# a_13613_37782# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9363 a_7039_65469# a_1586_66567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9364 a_13957_36121# a_12663_35431# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9365 a_6993_23555# a_4571_26677# a_6921_23555# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9366 a_25462_27497# a_24768_27247# a_3339_30503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.2245e+11p ps=7.66e+06u w=1e+06u l=150000u M=4
X9367 a_6277_14191# a_5903_13967# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=0p ps=0u w=650000u l=150000u
X9368 a_21382_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9369 a_17366_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X937 a_16510_8760# a_24703_35823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9370 a_25300_38567# a_24331_38591# a_25204_38567# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9371 vcm_commonmode a_16362_69222# a_41462_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9372 a_12481_54447# a_12203_54475# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X9373 VSS a_14926_31849# a_27169_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X9374 VDD a_10299_47607# a_10195_48437# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X9375 a_9184_13255# a_9227_12015# a_9326_13430# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9376 a_48794_65206# a_10975_66407# a_48398_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9377 a_34062_47607# a_24959_30503# a_34257_48169# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9378 VDD a_21049_34717# a_20655_34743# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9379 vcm_commonmode a_16362_64202# a_19374_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X938 a_29414_60186# a_16746_60188# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9380 a_6720_15279# a_5805_15279# a_6373_15521# VSS sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X9381 a_24698_23914# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9382 a_7802_49551# a_6725_49557# a_7640_49929# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9383 a_46390_63198# a_16362_63198# a_46482_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9384 a_2223_28617# a_2847_26133# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9385 a_9135_32143# a_3339_32463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X9386 a_2040_43401# a_1591_43029# a_1945_43023# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X9387 a_43378_9858# a_16362_9492# a_43470_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9388 a_36442_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9389 a_38754_57174# a_10515_22671# a_38358_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X939 VSS a_13809_48463# a_14421_49007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9390 VSS a_11067_13095# a_12895_13967# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9391 a_31822_57496# a_31768_55394# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9392 vcm_commonmode a_16362_68218# a_45478_68218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9393 a_8087_17289# a_7571_16917# a_7992_17277# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X9394 VDD a_7775_10625# a_7736_10499# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9395 a_19282_9858# a_16362_9492# a_19374_9492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9396 VDD a_19004_40413# a_18105_40157# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+11p ps=2.18e+06u w=800000u l=3.83e+06u
X9397 VDD a_12877_16911# a_49402_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9398 VDD a_25517_37455# a_41999_36367# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9399 VSS a_12877_16911# a_31726_12870# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X94 VDD a_5915_35943# a_8397_35407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X940 a_22690_61190# a_12355_15055# a_22294_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9400 a_34359_50639# a_34579_50613# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X9401 VSS a_12981_62313# a_43774_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9402 a_29414_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9403 a_40762_60186# a_39222_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9404 a_40762_19898# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9405 a_2764_31599# a_1683_31599# a_2417_31841# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X9406 a_23694_70226# a_18611_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9407 a_22386_68218# a_16746_68220# a_22294_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9408 vcm_commonmode a_16362_59182# a_48490_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9409 VSS a_9361_28335# a_9529_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u M=6
X941 a_4427_30511# a_3983_30761# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X9410 a_20514_28111# a_15681_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.4735e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X9411 a_21290_23914# a_16362_23548# a_21382_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9412 a_14471_30511# a_10506_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9413 VDD a_13848_44135# a_13661_43957# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9414 a_37354_24918# VSS a_37846_24520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9415 a_77086_40693# a_76346_40594# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=500000u M=2
X9416 VDD a_7390_32693# a_7695_31573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9417 a_30816_39429# a_29943_39141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9418 a_41862_22512# a_40675_27791# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9419 VSS a_43003_30761# a_23395_32463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X942 VDD a_11067_13095# a_12877_14441# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X9420 a_19743_38007# a_18811_38053# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9421 a_6927_40847# a_5885_39759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9422 a_75445_40202# a_75541_40024# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9423 VDD a_12355_65103# a_44382_64202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9424 a_7815_42453# a_7640_42479# a_7994_42479# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9425 a_20682_63198# a_15439_49525# a_20286_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9426 VSS a_33856_44869# a_33819_44535# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X9427 a_26706_61190# a_21371_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9428 a_25398_59182# a_16746_59184# a_25306_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9429 VSS a_10935_11989# a_9491_12297# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X943 a_28599_28023# a_13643_28327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X9430 VSS a_12869_2741# a_12899_2767# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9431 VSS a_12895_13967# a_30722_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9432 a_51714_39886# a_51330_39932# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9433 VDD a_12713_41923# a_16556_40743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9434 VSS a_4792_20443# a_10151_21379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9435 VSS a_4578_40455# a_5594_36727# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.52e+11p ps=2.88e+06u w=420000u l=150000u
X9436 a_2325_49525# a_2107_49929# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9437 VDD a_12257_56623# a_34342_56170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9438 a_11599_61341# a_10975_60975# a_11491_60975# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X9439 VSS a_7377_18012# a_8581_18319# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X944 VSS a_4941_35727# a_6927_39215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X9440 a_45386_72234# VDD a_45878_72556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9441 a_35069_51433# a_35039_51335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6.55e+11p pd=5.31e+06u as=0p ps=0u w=1e+06u l=150000u
X9442 a_6162_28487# a_5211_24759# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u M=2
X9443 a_40050_48463# a_38067_47349# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9444 VSS a_4891_47388# a_23847_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9445 a_42374_14878# a_16362_14512# a_42466_14512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9446 a_32795_39679# a_31280_40517# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X9447 a_10865_72399# a_5877_70197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9448 a_39299_48783# a_16863_29415# a_39127_48463# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X9449 a_45878_60508# a_40050_48463# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X945 a_28410_65206# a_16746_65208# a_28318_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9450 VSS VDD a_46786_7850# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9451 a_17366_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9452 a_5557_74895# a_5441_72399# a_5475_74895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9453 a_29414_58178# a_16746_58180# a_29322_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9454 vcm_commonmode VSS a_26402_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9455 a_39758_9858# a_12985_19087# a_39362_9858# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9456 a_32334_70226# a_16362_70226# a_32426_70226# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9457 VDD a_22448_39429# a_22352_39429# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9458 a_31726_14878# a_31768_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9459 vcm_commonmode a_16362_22544# a_41462_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X946 a_44382_10862# a_16362_10496# a_44474_10496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9460 a_3693_68047# a_3215_68351# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9461 VDD VSS a_38358_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9462 VDD a_6095_44807# a_12203_54475# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9463 a_21611_47919# a_21261_47919# a_21516_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=0p ps=0u w=420000u l=150000u
X9464 a_18770_23516# a_8491_27023# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9465 a_22786_72556# a_17599_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9466 a_18370_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9467 a_11659_66567# a_12231_65301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9468 a_48890_12472# a_42709_29199# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9469 VDD a_12985_7663# a_22294_21906# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X947 a_34342_71230# a_12901_66665# a_34834_71552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9470 VDD a_20881_28111# a_20773_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X9471 a_27710_9858# a_27752_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9472 VSS a_5254_67503# a_7097_67655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9473 VDD a_4328_10761# a_4503_10687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9474 a_22294_62194# a_16362_62194# a_22386_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9475 a_43774_67214# a_41872_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9476 a_10730_28995# a_7841_29673# a_10648_28995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9477 a_12034_58077# a_10957_57711# a_11872_57711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9478 a_34434_17524# a_16746_17522# a_34342_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9479 a_4995_27791# a_3143_22364# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X948 a_8735_15113# a_8289_14741# a_8639_15113# VSS sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X9480 a_6514_37191# a_6883_37019# a_6817_37289# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9481 a_9509_27791# a_6773_27805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9482 a_38754_10862# a_12546_22351# a_38358_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9483 a_2215_51549# a_1591_51183# a_2107_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X9484 a_6060_15279# a_5943_15492# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9485 a_1853_27247# a_1683_27247# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X9486 VDD a_12473_36341# a_12885_36694# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9487 vcm_commonmode a_16362_21540# a_45478_21540# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9488 a_7862_34025# a_6662_34025# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=4
X9489 a_19282_15882# a_16362_15516# a_19374_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X949 a_17322_31171# a_4674_40277# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9490 VDD a_10055_58791# a_25306_12870# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9491 a_5547_21379# a_2317_28892# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X9492 a_2744_46983# a_2959_47113# a_2886_47158# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9493 a_23390_13508# a_16746_13506# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9494 a_48398_7850# VSS a_48490_7484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9495 VSS a_12983_63151# a_20682_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9496 a_43870_63520# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9497 a_38450_16520# a_16746_16518# a_38358_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9498 VDD a_15931_39859# a_15957_39655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9499 vcm_commonmode a_16362_13508# a_35438_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X95 a_3998_15823# a_3911_16065# a_3594_15955# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X950 a_35132_47695# a_15607_46805# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.8675e+11p pd=3.79e+06u as=0p ps=0u w=650000u l=150000u
X9500 a_47886_18496# a_43269_29967# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9501 a_18756_51005# a_6559_59879# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9502 a_6097_16609# a_5879_16367# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9503 vcm_commonmode a_16362_23548# a_18370_23548# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9504 a_4032_49159# a_3325_49551# a_4174_49334# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9505 vcm_commonmode a_16362_12504# a_48490_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9506 a_22386_21540# a_16746_21538# a_22294_21906# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9507 VSS a_3877_57167# a_4220_57685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9508 a_3998_15823# a_3872_15939# a_3594_15955# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X9509 VDD a_6649_25615# a_6782_29967# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X951 VDD a_12713_43011# a_19684_42693# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9510 VDD a_8583_33551# a_19439_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X9511 a_37750_58178# a_36613_48169# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9512 a_27337_38565# a_26447_39141# a_27320_39429# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9513 a_28426_29941# a_20267_30503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9514 a_34977_30511# a_32970_31145# a_34895_30511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9515 VDD a_15439_49525# a_20286_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9516 VDD a_12899_10927# a_24302_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9517 a_48490_7484# VDD a_48398_7850# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9518 a_31543_51335# a_32091_51157# a_31871_51433# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X9519 a_8071_44982# a_7889_44982# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X952 a_3026_9839# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X9520 a_5085_24759# a_6614_21237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9521 a_42866_69544# a_41261_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9522 a_25398_12504# a_16746_12502# a_25306_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9523 a_37446_63198# a_16746_63200# a_37354_63198# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9524 a_6927_56873# a_4119_70741# a_7009_56873# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X9525 a_42374_59182# a_16362_59182# a_42466_59182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9526 VSS a_32823_29397# a_32769_29423# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9527 a_2313_12015# a_1887_12342# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9528 a_17274_61190# a_12981_59343# a_17766_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9529 a_25306_69222# a_16362_69222# a_25398_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X953 a_30722_21906# a_30764_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9530 VSS a_12257_56623# a_27710_57174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9531 vcm_commonmode a_16362_9492# a_29414_9492# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9532 VDD a_17863_44211# a_17889_44007# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.99e+11p ps=4.42e+06u w=420000u l=150000u M=2
X9533 a_24683_27497# a_2235_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.345e+12p pd=1.269e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X9534 VSS a_43319_31029# a_43267_31055# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9535 a_31726_55166# VSS a_31330_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9536 a_5309_25853# a_5087_24643# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X9537 a_15457_47081# a_15607_46805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9538 a_4852_23413# a_3972_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X9539 a_43378_65206# a_12355_65103# a_43870_65528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X954 a_12489_47919# a_9989_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9540 VSS a_3983_12015# a_4065_12879# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9541 a_29414_11500# a_16746_11498# a_29322_11866# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9542 VDD a_12895_13967# a_28318_19898# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9543 a_9445_30761# a_8117_30287# a_9349_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9544 VSS a_12899_2767# a_33734_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9545 a_32730_63198# a_28547_51175# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9546 vcm_commonmode a_16362_71230# a_42466_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9547 VDD a_9276_12167# a_9227_12015# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9548 VSS a_32765_31287# a_31964_30485# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9549 a_29322_68218# a_16362_68218# a_29414_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X955 a_27314_20902# a_16362_20536# a_27406_20536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9550 a_28817_29111# a_38883_29217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X9551 VSS a_1591_72943# a_2169_74913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9552 VSS a_3751_72373# a_4073_72943# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9553 VDD a_12947_8725# a_21290_8854# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9554 a_9577_60437# a_9411_60437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9555 a_4993_32929# a_4775_32687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X9556 VSS a_12947_23413# a_46786_23914# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9557 VDD a_11619_63151# a_9513_65301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9558 a_43774_20902# a_40491_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9559 a_18053_29199# a_15851_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X956 a_38358_69222# a_16362_69222# a_38450_69222# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9560 a_7295_44647# a_17554_30663# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X9561 a_20778_65528# a_16955_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9562 a_46390_56170# a_12947_56817# a_46882_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9563 a_30326_22910# a_10515_23975# a_30818_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9564 VDD a_23395_32463# a_28671_30539# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9565 a_2405_20719# a_2228_20719# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9566 a_23390_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9567 VSS a_12473_36341# a_12892_36367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9568 a_20286_55166# VSS a_20378_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9569 a_10103_48682# a_10195_48437# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X957 VDD a_12981_62313# a_37354_62194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9570 VSS a_12727_13353# a_36746_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9571 VSS a_5085_23047# a_7841_22895# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9572 VSS a_24515_34789# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X9573 a_40762_13874# a_12877_16911# a_40366_13874# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9574 a_1757_38677# a_1591_38677# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9575 a_23790_17492# a_23736_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9576 a_20286_14878# a_12877_14441# a_20778_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9577 VSS a_12985_7663# a_20682_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9578 a_23694_23914# a_10515_23975# a_23298_23914# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9579 VDD a_11902_27497# a_19889_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u M=2
X958 a_33338_57174# a_12257_56623# a_33830_57496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9580 a_2012_30333# a_1895_30138# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9581 VSS a_4191_33449# a_21095_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9582 VDD a_2672_66415# a_2847_66389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9583 a_2928_22583# a_3143_22364# a_3070_22390# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9584 a_2229_16143# a_2004_42453# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9585 a_12412_32143# a_11711_32143# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9586 VSS a_12516_7093# a_45782_70226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9587 a_76648_40202# a_76744_40024# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9588 a_37354_58178# a_10515_22671# a_37846_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9589 a_8367_44343# a_8475_44343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X959 a_42466_67214# a_16746_67216# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9590 a_6985_52815# a_6467_53359# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X9591 a_28756_7638# a_32367_28309# a_32135_28335# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9592 vcm_commonmode VSS a_19374_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9593 a_37750_11866# a_36797_27497# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9594 a_10103_11079# a_9642_10357# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9595 a_19333_48463# a_18907_48502# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9596 vcm_commonmode a_16362_61190# a_49494_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9597 a_23390_70226# a_16746_70228# a_23298_70226# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9598 VSS a_7987_64213# a_7921_64239# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9599 VDD a_16510_8760# a_16746_9490# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u M=2
X96 a_49494_17524# a_16746_17522# a_49402_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X960 a_4119_70741# a_3668_56311# a_4811_65871# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u M=4
X9600 VSS a_12355_15055# a_35742_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9601 a_24302_13874# a_12727_15529# a_24794_13476# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9602 VDD a_10259_10703# a_10661_10383# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9603 a_27806_55488# a_23395_52047# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9604 VSS a_28446_31375# a_36711_29199# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X9605 VSS a_5331_18517# a_4792_20443# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u M=4
X9606 VDD a_4215_51157# a_16219_51183# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9607 a_17670_14878# a_12727_15529# a_17274_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9608 a_26402_61190# a_16746_61192# a_26310_61190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9609 VDD VSS a_36350_24918# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X961 a_44778_55166# VSS a_44382_55166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9610 vcm_commonmode a_16362_17524# a_23390_17524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9611 VDD a_4417_22671# a_4627_23439# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9612 VDD a_7773_63927# a_7539_63695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.5e+11p ps=5.3e+06u w=1e+06u l=150000u
X9613 VSS a_7803_11703# a_7755_11471# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X9614 a_8461_32937# a_6243_30662# a_8389_32937# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X9615 VSS a_12985_16367# a_27710_10862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9616 a_23928_28585# a_23303_28335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=150000u
X9617 VSS a_30835_39783# a_14963_39783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X9618 VSS a_27869_50095# a_28785_47919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9619 a_12132_51005# a_9240_53877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X962 VSS a_26753_37981# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X9620 a_21663_41855# a_20715_41245# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X9621 a_7075_49929# a_6559_49557# a_6980_49917# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X9622 a_24209_48463# a_23767_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9623 a_35687_29199# a_32823_29397# a_35553_29199# VSS sky130_fd_pr__nfet_01v8 ad=2.5025e+11p pd=2.07e+06u as=3.38e+11p ps=2.34e+06u w=650000u l=150000u
X9624 a_11399_71855# a_10883_71855# a_11304_71855# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X9625 VSS a_23567_43123# a_23507_43177# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u M=2
X9626 VSS a_15253_43421# a_14945_43781# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9627 a_15439_49525# a_15575_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X9628 a_32334_63198# a_12981_62313# a_32826_63520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9629 vcm_commonmode a_16362_16520# a_27406_16520# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X963 a_18370_57174# a_16746_57176# a_18278_57174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9630 a_37846_20504# a_36797_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9631 VDD VDD a_44382_72234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9632 a_2727_56417# a_1591_56623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9633 a_37446_16520# a_16746_16518# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9634 a_4712_23759# a_4417_22671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9635 a_5880_41641# a_5490_41365# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u M=4
X9636 a_31422_14512# a_16746_14510# a_31330_14878# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9637 a_30023_41959# a_1761_40847# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9638 a_7725_31599# a_5993_32687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9639 a_8682_41974# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X964 a_19678_18894# a_19720_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9640 VDD a_30052_32117# a_37471_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9641 VSS a_5411_12791# a_5227_13621# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X9642 a_44474_62194# a_16746_62196# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9643 a_43362_28879# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9644 a_26187_48801# a_6835_46823# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9645 a_40383_29575# a_32970_31145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9646 a_6614_10927# a_2292_17179# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9647 a_27406_72234# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9648 vcm_commonmode a_16362_69222# a_39454_69222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9649 a_29718_60186# a_12981_59343# a_29322_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X965 a_24674_31849# a_5363_30503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9650 a_29718_19898# a_12895_13967# a_29322_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9651 a_13692_34191# a_13515_34191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9652 a_43470_67214# a_16746_67216# a_43378_67214# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9653 vcm_commonmode a_16362_64202# a_40458_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9654 a_42374_22910# a_16362_22544# a_42466_22544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9655 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9656 a_38358_12870# a_16362_12504# a_38450_12504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9657 a_24800_41953# a_24331_40767# a_25263_41001# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9658 a_17366_64202# a_16746_64204# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9659 a_34738_61190# a_34780_56398# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X966 VDD a_49984_39288# a_49876_41198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=3.32e+06u w=500000u l=150000u M=4
X9660 a_31330_69222# a_12901_66959# a_31822_69544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9661 a_33430_59182# a_16746_59184# a_33338_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9662 VSS a_75728_39738# a_75541_39480# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9663 vcm_commonmode a_16362_63198# a_26402_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9664 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9665 a_1887_12342# a_1761_11471# a_1815_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9666 VDD a_2606_41079# a_4500_45289# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9667 a_17670_71230# a_13183_52047# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9668 a_16362_69222# a_12907_56399# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X9669 a_6607_39991# a_3949_41935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X967 VSS a_12899_11471# a_23694_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9670 VSS a_35033_42044# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X9671 VDD a_2319_63388# a_2250_63517# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=840000u l=150000u
X9672 VSS a_36116_44765# a_36395_44265# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u M=2
X9673 VDD a_10299_11703# a_9642_10357# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.75e+11p ps=2.95e+06u w=1e+06u l=150000u
X9674 a_4496_18543# a_4379_18756# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9675 a_18811_36965# a_15305_38543# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X9676 a_2417_31841# a_2199_31599# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9677 a_2557_57711# a_1923_54591# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9678 a_18278_60186# a_16362_60186# a_18370_60186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9679 a_32426_21540# a_16746_21538# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X968 a_19743_36919# a_18811_36965# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.52e+11p pd=6.68e+06u as=0p ps=0u w=800000u l=150000u
X9680 VDD a_2847_26133# a_2834_26525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9681 VSS a_2787_32679# a_5767_31573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9682 vcm_commonmode VSS a_34434_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9683 a_11626_28335# a_7571_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9684 a_5925_69929# a_3143_66972# a_6180_69929# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X9685 vcm_commonmode a_16362_65206# a_17366_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9686 a_11163_25321# a_11057_25077# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9687 VDD a_5631_38127# a_7910_38671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9688 a_22690_24918# a_12341_3311# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9689 a_10475_14165# a_10678_14443# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X969 a_20682_13874# a_9503_26151# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9690 a_19282_23914# a_16362_23548# a_19374_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9691 VSS a_37699_27221# a_25744_7638# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9692 VSS a_1761_25615# a_1959_26703# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X9693 a_21856_36513# a_21663_35327# a_22536_35303# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9694 a_36746_58178# a_12901_58799# a_36350_58178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9695 a_17507_30761# a_17554_30663# a_17771_30761# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u M=2
X9696 VDD a_5831_39189# a_7889_44982# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9697 a_47790_9858# a_12985_19087# a_47394_9858# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9698 a_43870_71552# a_41872_29423# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9699 a_19678_68218# a_12901_66959# a_19282_68218# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X97 a_20378_23548# a_16746_23546# a_20286_23914# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X970 a_13390_29575# a_15207_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9700 a_39854_61512# a_39389_52271# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9701 VDD a_3203_17620# a_1895_18756# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X9702 a_28152_40517# a_27183_40229# a_28115_40183# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9703 a_47486_69222# a_16746_69224# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9704 a_49798_57174# a_10515_22671# a_49402_57174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9705 a_2215_23439# a_1591_23445# a_2107_23817# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X9706 VSS a_10471_65002# a_8999_61493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9707 VSS a_12895_13967# a_28714_18894# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9708 a_25702_15882# a_25744_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9709 VDD a_9869_49525# a_9759_49551# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X971 a_9186_54223# a_7155_55509# a_9376_54223# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.6725e+11p ps=3.73e+06u w=650000u l=150000u
X9710 a_5239_65301# a_1923_59583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9711 a_31522_32259# a_27535_30503# a_31440_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9712 a_5791_43541# a_5616_43567# a_5970_43567# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9713 a_28048_52093# a_6467_55527# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X9714 a_16244_34973# a_15775_34239# a_16707_34473# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9715 VDD a_12947_71576# a_20286_71230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9716 a_2325_40545# a_2107_40303# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X9717 VDD a_3020_54135# a_2327_54135# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9718 VSS a_10975_66407# a_41766_66210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9719 a_34342_8854# a_12985_19087# a_34834_8456# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X972 VDD a_14421_49007# a_12516_7093# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=6
X9720 a_3541_19385# a_2143_15271# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9721 VDD a_5800_71855# a_5975_71829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9722 a_2080_58077# a_1643_57685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9723 a_12727_13353# a_11067_13095# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u M=3
X9724 a_29718_14878# a_29760_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9725 vcm_commonmode a_16362_22544# a_39454_22544# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9726 VDD a_2473_34293# a_5253_29673# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9727 a_25687_32259# a_13357_32143# a_25605_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9728 a_43470_20536# a_16746_20534# a_43378_20902# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9729 a_38358_57174# a_16362_57174# a_38450_57174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X973 a_21382_10496# a_16746_10494# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9730 a_44874_8456# a_42718_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9731 a_40762_8854# a_39673_28111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9732 a_23987_39126# a_24029_39355# a_23987_39453# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9733 a_42466_55166# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9734 a_31726_63198# a_15439_49525# a_31330_63198# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9735 VDD a_12899_10927# a_32334_18894# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9736 VDD a_23501_42583# a_18662_43671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9737 a_27239_36341# a_12641_37684# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9738 a_13445_50639# a_12967_50943# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9739 a_33430_12504# a_16746_12502# a_33338_12870# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X974 a_2080_63517# a_1643_63125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9740 VDD a_12899_11471# a_45386_17890# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9741 a_5823_44905# a_5173_44655# a_5905_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X9742 a_42866_14480# a_41967_31375# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9743 a_40366_15882# a_16362_15516# a_40458_15516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9744 a_1887_12015# a_1633_12342# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9745 a_43470_18528# a_16746_18526# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9746 a_10216_67503# a_9301_67503# a_9869_67745# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9747 a_16362_22544# a_11067_23759# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u M=2
X9748 a_25798_24520# a_25744_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9749 VDD a_23172_31573# a_23119_31599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X975 VDD a_2847_26133# a_2223_28617# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u M=2
X9750 VSS a_12985_19087# a_26706_8854# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9751 a_11143_31599# a_10870_31599# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9752 a_2216_28309# a_2847_36799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9753 VSS a_9184_49159# a_7251_50069# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9754 VSS a_12983_63151# a_18674_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9755 VSS a_2007_65002# a_1895_66628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X9756 a_30356_42919# a_29483_42943# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9757 VSS a_6224_73095# a_7581_74031# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9758 a_22690_65206# a_10975_66407# a_22294_65206# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9759 VSS a_12947_56817# a_48794_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X976 a_12126_72221# a_11049_71855# a_11964_71855# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9760 a_77086_40693# VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9761 a_5185_44905# a_1689_10396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9762 a_46882_13476# a_43175_28335# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9763 a_43378_10862# a_12985_16367# a_43870_10464# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9764 VDD VSS a_49402_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9765 VDD a_12901_66959# a_40366_68218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9766 a_20286_63198# a_16362_63198# a_20378_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9767 a_26310_20902# a_12985_7663# a_26802_20504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9768 a_29814_23516# a_29760_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9769 a_29414_19532# a_16746_19530# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X977 a_33734_12870# a_32951_27247# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9770 a_37520_49783# a_4351_67279# a_37751_49667# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9771 a_41766_68218# a_41427_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9772 a_4564_63695# a_4127_63669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9773 a_26310_16886# a_16362_16520# a_26402_16520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9774 a_15681_27247# a_10964_25615# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=2
X9775 VDD a_12901_58799# a_36350_58178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9776 a_30418_14512# a_16746_14510# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9777 a_8304_39465# a_8251_39367# a_8209_39465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X9778 a_7794_53903# a_7764_53877# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=9.65e+11p pd=7.93e+06u as=0p ps=0u w=1e+06u l=150000u
X9779 a_33338_62194# a_16362_62194# a_33430_62194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X978 a_45782_63198# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9780 a_36746_11866# a_12985_16367# a_36350_11866# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9781 VSS a_5831_39189# a_7889_44982# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9782 result_out[5] a_1644_62037# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9783 a_12410_65327# a_1950_59887# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9784 a_33727_39913# a_32795_39679# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9785 a_45478_17524# a_16746_17522# a_45386_17890# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9786 a_25702_56170# a_12257_56623# a_25306_56170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9787 a_19774_15484# a_19720_7638# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9788 a_19678_21906# a_12985_7663# a_19282_21906# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9789 VDD a_12877_16911# a_23298_13874# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X979 vcm_commonmode a_16362_58178# a_41462_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9790 a_49798_10862# a_12546_22351# a_49402_10862# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9791 a_28430_32143# a_14646_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9792 vcm_commonmode a_16362_67214# a_32426_67214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9793 a_20778_10464# a_9503_26151# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9794 VSS a_7244_39189# a_8001_40125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X9795 a_3316_42313# a_2401_41941# a_2969_41909# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X9796 conversion_finished_out a_1644_77813# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u M=2
X9797 a_24673_49007# a_8531_70543# a_23830_49525# VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9798 a_37354_66210# a_10975_66407# a_37846_66532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9799 a_28318_8854# a_16362_8488# a_28410_8488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X98 VDD a_32367_28309# a_28756_7638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.48e+11p ps=2.78e+06u w=700000u l=150000u
X980 a_10883_11177# a_10661_10383# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X9800 a_23298_7850# VDD a_23790_7452# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9801 a_41862_64524# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9802 VDD a_2163_57853# a_2124_57979# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9803 vcm_commonmode a_16362_8488# a_42466_8488# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9804 vcm_commonmode a_16362_59182# a_22386_59182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9805 vcm_commonmode VSS a_16362_24552# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9806 VSS a_2163_56765# a_2124_56891# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9807 a_49494_16520# a_16746_16518# a_49402_16886# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9808 vcm_commonmode a_16362_13508# a_46482_13508# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9809 a_32795_38591# a_32029_38565# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X981 a_10497_10703# a_9484_11989# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X9810 a_25484_37253# a_24515_36965# a_25388_37253# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9811 a_5595_12167# a_5867_11995# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9812 VDD a_2672_39049# a_2847_38975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9813 VDD a_12516_7093# a_17274_69222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9814 VDD a_7580_61751# a_7577_60137# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9815 a_36448_47375# a_26523_28111# a_36275_47695# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.705e+11p ps=3.74e+06u w=650000u l=150000u
X9816 a_34725_37479# a_35033_37692# a_34699_37683# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X9817 VSS a_5595_33205# a_4563_32900# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9818 a_48794_58178# a_42985_46831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9819 VSS a_6435_10901# a_6369_10927# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X982 VSS a_8003_72917# a_9789_73807# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X9820 VDD a_22448_38341# a_22352_38341# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u M=2
X9821 a_42374_60186# a_12727_58255# a_42866_60508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9822 a_2847_69439# a_2672_69513# a_3026_69501# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X9823 a_12139_18517# a_2411_19605# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9824 a_28410_8488# a_16746_8486# a_28318_8854# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9825 VSS a_3911_16065# a_3872_15939# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9826 VSS a_26661_34428# a_26353_34215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9827 a_30415_50871# a_4482_57863# a_30561_50959# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X9828 VDD a_15439_49525# a_31330_63198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9829 VSS a_27359_43985# a_27305_44011# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X983 a_4339_64521# a_10239_57167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9830 a_30743_30287# a_18979_30287# a_30440_31573# VSS sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=0p ps=0u w=650000u l=150000u
X9831 a_6260_10927# a_5179_10927# a_5913_11169# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X9832 VDD a_14361_29967# a_14679_31288# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9833 VSS a_16863_29415# a_40218_27247# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X9834 a_18770_65528# a_14287_51175# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9835 a_7917_13885# a_7917_12265# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X9836 a_8251_39367# a_7910_38671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9837 VSS a_10515_22671# a_25702_58178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9838 VSS a_12901_66665# a_39758_71230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9839 a_35438_66210# a_16746_66212# a_35346_66210# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X984 a_30440_31573# a_30565_30199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9840 a_32334_71230# a_12901_66665# a_32826_71552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9841 a_28318_61190# a_12981_59343# a_28810_61512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9842 a_37446_24552# VDD vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9843 a_41397_30333# a_32823_29397# a_41325_30333# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X9844 a_27417_32509# a_27387_32373# a_27167_32143# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X9845 a_41795_31055# a_20359_29199# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=0p ps=0u w=1e+06u l=150000u
X9846 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X9847 VSS a_7931_10357# a_7862_10383# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9848 VSS a_12985_7663# a_18674_20902# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9849 a_6243_30662# a_5906_28585# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X985 a_7653_20291# a_7377_18012# a_7571_20291# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9850 a_15189_51433# a_14983_51157# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9851 a_33734_61190# a_12355_15055# a_33338_61190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9852 a_19780_41605# a_18811_41317# a_19684_41605# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9853 a_3203_47158# a_2952_46805# a_2744_46983# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X9854 a_30534_49393# a_30525_49551# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9855 a_2656_70197# a_2824_70197# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X9856 a_33761_28111# a_32823_29397# a_33689_28111# VSS sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X9857 vcm_commonmode VSS a_40458_72234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9858 a_39454_65206# a_16746_65208# a_39362_65206# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9859 a_30418_59182# a_16746_59184# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X986 a_47790_7850# a_43269_29967# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9860 a_6792_43719# a_7000_43541# a_6934_43567# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9861 VDD a_1923_54591# a_1643_54421# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9862 a_9276_12167# a_9491_12297# a_9418_12342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X9863 a_44382_18894# a_12895_13967# a_44874_18496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9864 a_41766_21906# a_40675_27791# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9865 VSS VSS a_44778_24918# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9866 a_38358_20902# a_16362_20536# a_38450_20536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9867 a_1849_33237# a_1683_33237# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9868 a_30722_66210# a_25971_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9869 VSS a_40581_31599# a_42941_32143# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X987 a_24302_59182# a_12901_58799# a_24794_59504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9870 a_7829_60431# a_7449_60431# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X9871 vcm_commonmode VSS a_31422_7484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9872 VSS a_7295_44647# a_35765_30287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9873 a_7479_36495# a_7381_35407# a_7561_36495# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9874 a_37750_60186# a_12981_59343# a_37354_60186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9875 a_76082_39738# a_76178_39480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9876 a_37750_19898# a_12895_13967# a_37354_19898# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9877 a_35647_35877# a_33963_35507# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X9878 VSS a_12899_11471# a_34738_16886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9879 vcm_commonmode a_16362_20536# a_32426_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X988 VDD a_12349_25847# a_15681_27497# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u M=2
X9880 a_19459_29423# a_18829_29423# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9881 a_31330_55166# VSS a_31422_55166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9882 a_7295_32259# a_7281_29423# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X9883 a_48490_71230# a_16746_71232# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9884 a_36541_48169# a_19807_28111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9885 VSS a_12727_13353# a_47790_15882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9886 a_21782_18496# a_9135_27239# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9887 a_21686_24918# VSS a_21290_24918# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9888 a_30418_71230# a_16746_71232# a_30326_71230# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9889 a_5135_47414# a_4563_32900# a_4676_47607# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.864e+11p ps=2.68e+06u w=420000u l=150000u
X989 a_2847_40277# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X9890 a_12587_51335# a_2840_66103# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9891 VDD a_12985_19087# a_39362_9858# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9892 vcm_commonmode a_16362_12504# a_22386_12504# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9893 vcm_commonmode a_16362_63198# a_34434_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9894 a_31330_14878# a_12877_14441# a_31822_14480# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9895 a_35346_59182# a_12901_58799# a_35838_59504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9896 a_32334_18894# a_16362_18528# a_32426_18528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9897 a_8857_14709# a_8639_15113# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9898 vcm_commonmode a_16362_62194# a_47486_62194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9899 a_27314_9858# a_12546_22351# a_27806_9460# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X99 VSS a_7519_59575# a_7299_59663# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X990 a_1770_14441# a_1591_14191# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u M=4
X9900 a_48398_58178# a_10515_22671# a_48890_58500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9901 VDD a_7373_40847# a_7999_40553# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9902 a_24698_57174# a_18151_52263# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9903 a_9485_62613# a_9319_62613# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X9904 VSS a_75728_40202# a_75541_40024# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9905 a_5418_45743# a_2292_43291# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9906 a_24698_15882# a_12877_14441# a_24302_15882# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9907 a_48794_11866# a_42709_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9908 VDD a_16012_41959# a_15189_39889# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9909 a_12754_18115# a_10055_58791# a_12672_18115# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X991 vcm_commonmode a_16362_20536# a_34434_20536# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9910 a_9457_71677# a_8575_74853# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9911 a_36442_11500# a_16746_11498# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9912 VSS a_22562_28023# a_22567_27791# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8025e+11p ps=3.77e+06u w=650000u l=150000u
X9913 a_23987_39453# a_23733_39126# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9914 VDD a_11395_62037# a_11299_62215# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X9915 a_24394_62194# a_16746_62196# a_24302_62194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9916 VDD a_4792_20443# a_12353_20969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X9917 VDD a_3983_44655# a_2606_41079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u M=4
X9918 VSS a_4036_51157# a_1586_51335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u M=2
X9919 vcm_commonmode a_16362_18528# a_21382_18528# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X992 a_43378_22910# a_10515_23975# a_43870_22512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9920 a_25798_58500# a_21371_50959# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9921 VDD a_2843_71829# a_5087_72512# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9922 a_28714_14878# a_12727_15529# a_28318_14878# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9923 VSS a_10055_58791# a_25702_11866# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9924 a_20743_43493# a_19780_41605# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.83e+06u
X9925 a_35379_49871# a_2840_66103# a_35307_49871# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X9926 a_2215_40669# a_2411_26133# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9927 VSS config_1_in[11] a_1626_19087# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9928 VSS a_2319_64476# a_2250_64605# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9929 VDD a_75794_38962# a_77451_38925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=4.74e+06u w=500000u l=500000u M=2
X993 a_3983_25321# a_2315_24540# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X9930 a_8540_42167# a_8273_42479# a_8682_41974# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X9931 VSS a_11710_58487# a_11699_58799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X9932 VSS a_1586_40455# a_1591_44655# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9933 a_23593_42919# a_23901_43132# a_23567_43123# VSS sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X9934 a_29322_69222# a_12901_66959# a_29814_69544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9935 VDD a_4191_33449# a_21095_47919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9936 a_12134_69679# a_8575_74853# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X9937 VSS a_11067_13095# a_37750_64202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9938 a_30326_64202# a_11067_13095# a_30818_64524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9939 a_32544_30083# a_26523_29199# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X994 a_36442_58178# a_16746_58180# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9940 a_49798_8854# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X9941 a_35838_21508# a_35601_27497# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9942 a_35438_17524# a_16746_17522# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9943 a_30115_38695# a_1761_43567# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u M=2
X9944 VSS a_10506_29967# a_14013_30083# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9945 a_16556_40743# a_15683_40767# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9946 a_24331_44581# a_22632_42919# VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X9947 a_38358_65206# a_16362_65206# a_38450_65206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9948 a_4871_32687# a_4425_32687# a_4775_32687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9949 a_42466_63198# a_16746_63200# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X995 VDD a_17711_32385# a_17672_32259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9950 a_6934_43894# a_5831_39189# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9951 a_20286_56170# a_12947_56817# a_20778_56492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X9952 a_42770_70226# a_41261_28335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9953 a_41462_68218# a_16746_68220# a_41370_68218# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9954 VDD a_19877_41972# a_13349_37973# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X9955 VSS a_12231_65301# a_12165_65327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9956 VDD a_16228_28335# a_17459_31145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9957 a_24800_35425# a_24331_34239# a_25263_34473# VDD sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9958 a_1757_49557# a_1591_49557# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9959 a_40366_23914# a_16362_23548# a_40458_23548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X996 VDD a_12727_67753# a_49402_67214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9960 VSS a_17222_27247# a_19611_28335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9175e+11p ps=1.89e+06u w=650000u l=150000u
X9961 a_18257_47741# a_18222_47507# a_17787_47349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9962 a_36350_13874# a_16362_13508# a_36442_13508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9963 a_7479_36495# a_7381_35407# a_7561_36815# VSS sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X9964 a_9927_60809# a_9411_60437# a_9832_60797# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X9965 a_10409_18543# a_9983_18870# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9966 a_24302_55166# VSS a_24794_55488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9967 a_45782_61190# a_40050_48463# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9968 a_44474_59182# a_16746_59184# a_44382_59182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9969 vcm_commonmode a_16362_56170# a_41462_56170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X997 VSS a_12981_62313# a_22690_63198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9970 a_4595_20719# a_4149_20719# a_4499_20719# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9971 a_12621_44099# a_21479_44581# a_22352_44869# VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9972 a_28714_71230# a_28756_55394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9973 a_27406_69222# a_16746_69224# a_27314_69222# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9974 a_22836_30287# a_5915_30287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X9975 VDD a_2847_19605# a_2834_19997# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9976 a_33830_24520# a_12899_2767# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9977 a_4972_51017# a_4057_50645# a_4625_50613# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X9978 a_22386_9492# a_16746_9490# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9979 a_26310_24918# VSS a_26402_24552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X998 a_21123_30511# a_21057_30669# a_20821_30511# VSS sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=4.355e+11p ps=3.94e+06u w=650000u l=150000u
X9980 a_2217_35113# a_2011_34837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X9981 VDD a_12983_63151# a_36350_66210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9982 a_6361_44655# a_5823_44905# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9983 a_24698_10862# a_24740_7638# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9984 a_30418_22544# a_16746_22542# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9985 a_11390_21807# a_6559_22671# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u M=4
X9986 a_36442_56170# a_16746_56172# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9987 VSS a_12981_59343# a_22690_61190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9988 a_49798_60186# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9989 a_48490_58178# a_16746_58180# a_48398_58178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X999 a_5839_22351# a_5588_22467# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9990 a_49798_19898# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9991 a_38969_29217# a_38210_30199# a_38883_29217# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9992 a_19374_66210# a_16746_66212# vcm_commonmode VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X9993 vcm_commonmode VSS a_45478_55166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9994 VDD a_12985_16367# a_19282_11866# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X9995 vcm_commonmode a_16362_65206# a_28410_65206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9996 a_23564_31849# a_14646_29423# a_23309_31849# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X9997 a_34342_20902# a_12985_7663# a_34834_20504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X9998 VDD a_3162_43023# a_3339_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8e+11p ps=7.6e+06u w=1e+06u l=150000u M=5
X9999 a_41862_72556# a_41427_52263# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
C0 vcm_commonmode a_17366_55166# 0.84fF
C1 a_16101_31029# a_13390_29575# 0.59fF
C2 a_28410_10496# VDD 0.51fF
C3 a_33155_40191# VDD 0.73fF
C4 a_36613_48169# a_37446_65206# 0.38fF
C5 vcm_commonmode a_48490_64202# 0.87fF
C6 a_2292_43291# a_1586_45431# 0.86fF
C7 a_16891_49220# VDD 0.63fF
C8 a_25398_72234# a_25398_71230# 1.00fF
C9 a_43470_60186# VDD 0.51fF
C10 vcm_commonmode a_35346_10862# 0.31fF
C11 a_12899_3855# a_32772_7638# 0.68fF
C12 a_37446_67214# a_37446_66210# 1.00fF
C13 vcm_commonmode a_27406_23548# 0.87fF
C14 a_10515_63143# a_4495_35925# 0.33fF
C15 a_24394_7484# m3_24296_7346# 2.80fF
C16 vcm_commonmode a_24394_66210# 0.87fF
C17 a_9135_27239# a_21382_17524# 0.38fF
C18 a_16746_61192# a_12981_59343# 0.41fF
C19 a_33430_65206# a_33430_64202# 1.00fF
C20 a_2011_34837# VDD 3.50fF
C21 vcm_commonmode a_36442_19532# 0.87fF
C22 ctopn a_18370_16520# 3.58fF
C23 a_1761_25071# a_12473_42869# 0.79fF
C24 vcm_commonmode a_22294_62194# 0.31fF
C25 a_25787_28327# a_33430_57174# 0.38fF
C26 a_42985_46831# a_12257_56623# 0.40fF
C27 a_23390_15516# VDD 0.51fF
C28 a_17449_46831# VDD 0.62fF
C29 a_38557_32143# a_38450_70226# 0.38fF
C30 a_17366_19532# a_18370_19532# 0.97fF
C31 m3_25300_7346# VDD 0.40fF
C32 a_27406_23548# a_27406_22544# 1.00fF
C33 a_24740_7638# a_12985_19087# 0.41fF
C34 a_13643_28327# a_6459_30511# 0.45fF
C35 a_3854_29977# VDD 0.36fF
C36 vcm_commonmode a_30326_15882# 0.31fF
C37 a_23390_63198# ctopp 3.64fF
C38 a_3780_56347# a_6646_54135# 0.47fF
C39 a_36350_56170# a_36442_56170# 0.32fF
C40 a_21382_71230# VDD 0.58fF
C41 a_41872_29423# a_10515_22671# 0.40fF
C42 a_21382_66210# a_21382_65206# 1.00fF
C43 a_2292_17179# a_7775_10625# 0.33fF
C44 a_22386_14512# a_23390_14512# 0.97fF
C45 a_15683_39141# VDD 1.02fF
C46 a_33430_11500# VDD 0.51fF
C47 a_18915_42089# VDD 0.62fF
C48 a_39222_48169# a_40458_66210# 0.38fF
C49 a_38450_69222# a_39454_69222# 0.97fF
C50 a_29760_7638# a_29414_9492# 0.38fF
C51 ctopn a_17712_7638# 2.36fF
C52 a_4495_35925# a_3607_34639# 1.45fF
C53 a_28756_55394# a_29760_55394# 0.63fF
C54 a_17599_52263# a_34251_52263# 0.35fF
C55 vcm_commonmode a_28318_71230# 0.31fF
C56 a_33430_61190# a_33430_60186# 1.00fF
C57 a_19282_8854# a_19374_8488# 0.32fF
C58 a_37446_24552# VDD 0.60fF
C59 vcm_commonmode a_40366_11866# 0.31fF
C60 a_17366_59182# ctopp 3.43fF
C61 a_48490_64202# a_49494_64202# 0.97fF
C62 a_3247_20495# a_4314_40821# 0.80fF
C63 a_17507_52047# a_2959_47113# 2.31fF
C64 a_39389_52271# a_39454_62194# 0.38fF
C65 vcm_commonmode a_44382_24918# 0.31fF
C66 a_20286_70226# a_20378_70226# 0.32fF
C67 a_4831_58497# a_4792_58371# 0.74fF
C68 a_37354_58178# a_37446_58178# 0.32fF
C69 a_47486_55166# VDD 0.58fF
C70 a_27752_7638# a_12985_16367# 0.41fF
C71 a_45478_22544# a_46482_22544# 0.97fF
C72 a_6835_46823# a_7000_43541# 0.36fF
C73 a_19374_62194# a_19374_61190# 1.00fF
C74 a_14273_27791# VDD 0.51fF
C75 a_39454_57174# VDD 0.51fF
C76 a_36442_65206# a_37446_65206# 0.97fF
C77 vcm_commonmode a_39454_20536# 0.87fF
C78 a_8583_33551# a_32143_35281# 0.76fF
C79 vcm_commonmode a_28410_63198# 0.92fF
C80 a_32426_17524# a_32426_16520# 1.00fF
C81 a_5363_16367# a_5529_16367# 0.69fF
C82 vcm_commonmode a_46390_57174# 0.31fF
C83 a_12355_15055# a_8273_42479# 0.57fF
C84 a_19374_20536# a_19374_19532# 1.00fF
C85 a_27406_23548# a_28410_23548# 0.97fF
C86 a_2840_66103# a_5190_59575# 0.46fF
C87 a_28089_31157# VDD 0.35fF
C88 a_47486_58178# ctopp 3.58fF
C89 a_28410_72234# VDD 1.24fF
C90 a_24394_66210# a_25398_66210# 0.97fF
C91 vcm_commonmode a_22386_59182# 0.87fF
C92 a_31768_55394# a_12727_58255# 0.40fF
C93 a_6725_42479# VDD 0.46fF
C94 a_28883_52031# VDD 0.36fF
C95 a_7925_72399# a_7707_70741# 0.65fF
C96 vcm_commonmode a_33430_72234# 0.69fF
C97 a_19720_7638# a_12727_13353# 0.41fF
C98 a_26550_40871# a_33963_35507# 0.41fF
C99 a_35346_61190# a_35438_61190# 0.32fF
C100 vcm_commonmode a_39454_12504# 0.87fF
C101 a_21382_60186# ctopp 3.59fF
C102 ctopn a_40458_9492# 3.58fF
C103 a_37919_28111# a_38450_23548# 0.38fF
C104 a_24394_68218# VDD 0.51fF
C105 a_27429_35301# VDD 1.42fF
C106 a_24302_7850# VDD 0.62fF
C107 ctopn a_20378_22544# 3.58fF
C108 a_27535_30503# a_20267_30503# 0.32fF
C109 vcm_commonmode a_31330_68218# 0.31fF
C110 a_24394_71230# a_24394_70226# 1.00fF
C111 a_36442_19532# a_37446_19532# 0.97fF
C112 a_46482_23548# a_46482_22544# 1.00fF
C113 a_6559_22671# a_5449_25071# 0.63fF
C114 a_15607_46805# a_32823_29397# 1.20fF
C115 a_8383_27247# VDD 0.62fF
C116 a_7987_64213# a_4339_64521# 0.38fF
C117 a_40458_66210# a_40458_65206# 1.00fF
C118 a_17599_52263# a_8491_57487# 1.41fF
C119 a_41462_14512# a_42466_14512# 0.97fF
C120 a_11067_67279# a_40675_27791# 0.41fF
C121 vcm_commonmode a_34434_21540# 0.87fF
C122 a_6224_73095# a_2952_66139# 0.39fF
C123 a_20378_20536# a_21382_20536# 0.97fF
C124 a_38358_8854# a_38450_8488# 0.32fF
C125 a_11067_13095# a_2959_47113# 0.99fF
C126 a_6515_62037# a_7210_55081# 1.17fF
C127 vcm_commonmode a_39454_17524# 0.87fF
C128 ctopn a_16362_14512# 1.35fF
C129 vcm_commonmode a_26402_60186# 0.87fF
C130 a_38450_13508# VDD 0.51fF
C131 a_39362_70226# a_39454_70226# 0.32fF
C132 a_1761_40847# a_12663_35431# 2.85fF
C133 a_6835_46823# a_7553_48469# 0.35fF
C134 a_38450_62194# a_38450_61190# 1.00fF
C135 a_29414_10496# a_29414_9492# 1.00fF
C136 a_11866_27791# VDD 1.74fF
C137 a_24394_56170# VDD 0.52fF
C138 vcm_commonmode a_45386_13874# 0.31fF
C139 a_19720_7638# a_10515_23975# 0.41fF
C140 a_1586_21959# a_4149_20719# 0.63fF
C141 a_20286_16886# a_20378_16520# 0.32fF
C142 vcm_commonmode a_31330_56170# 0.31fF
C143 ctopn a_21382_23548# 3.40fF
C144 a_26514_47375# VDD 1.59fF
C145 a_5671_21495# a_10543_16580# 0.41fF
C146 a_38450_20536# a_38450_19532# 1.00fF
C147 a_46482_23548# a_47486_23548# 0.97fF
C148 a_30023_41959# a_26433_39631# 0.89fF
C149 a_17366_57174# ctopp 3.24fF
C150 a_43470_66210# a_44474_66210# 0.97fF
C151 ctopn a_30418_19532# 3.59fF
C152 a_41842_27221# a_26523_29199# 0.46fF
C153 a_10506_29967# a_14361_29967# 0.40fF
C154 a_42985_46831# a_10975_66407# 0.40fF
C155 a_33313_51157# VDD 0.64fF
C156 a_40491_27247# a_12727_13353# 0.41fF
C157 a_18370_21540# a_18370_20536# 1.00fF
C158 a_8491_27023# a_12985_16367# 0.41fF
C159 a_23390_61190# VDD 0.51fF
C160 vcm_commonmode a_16362_11500# 4.47fF
C161 a_43175_28335# a_46482_22544# 0.38fF
C162 a_40491_27247# a_43470_23548# 0.38fF
C163 a_20378_12504# a_21382_12504# 0.97fF
C164 a_33486_34191# VDD 0.41fF
C165 vcm_commonmode a_40458_18528# 0.87fF
C166 a_26310_67214# a_26402_67214# 0.32fF
C167 vcm_commonmode a_30326_61190# 0.31fF
C168 a_2143_15271# a_10883_11177# 0.33fF
C169 vcm_commonmode a_20378_24552# 0.84fF
C170 a_43470_71230# a_43470_70226# 1.00fF
C171 a_39299_48783# a_44474_69222# 0.38fF
C172 a_18053_28879# VDD 1.44fF
C173 a_10055_58791# a_31768_7638# 0.41fF
C174 a_31422_62194# ctopp 3.59fF
C175 a_26433_39631# a_1799_29556# 0.52fF
C176 a_26550_40871# a_27263_40871# 0.59fF
C177 a_27406_70226# VDD 0.51fF
C178 vcm_commonmode a_31422_55166# 0.84fF
C179 a_11719_28023# a_9529_28335# 1.61fF
C180 a_18105_40157# VDD 1.03fF
C181 vcm_commonmode a_22386_57174# 0.87fF
C182 a_21187_29415# a_22015_28111# 7.18fF
C183 a_41872_29423# a_12901_66665# 0.40fF
C184 vcm_commonmode a_34342_70226# 0.31fF
C185 a_6816_19355# a_2292_17179# 0.48fF
C186 a_39454_20536# a_40458_20536# 0.97fF
C187 vcm_commonmode a_49494_10496# 0.90fF
C188 a_28410_63198# a_29414_63198# 0.97fF
C189 a_4339_64521# a_10680_52245# 0.42fF
C190 a_4885_71855# VDD 0.50fF
C191 a_37446_71230# ctopp 3.40fF
C192 ctopn a_33430_20536# 3.59fF
C193 a_15253_43421# VDD 0.97fF
C194 a_5682_69367# a_8782_65015# 0.63fF
C195 a_28318_58178# a_28410_58178# 0.32fF
C196 a_23193_52245# VDD 0.68fF
C197 a_3751_72373# a_2843_71829# 0.34fF
C198 a_6559_59663# a_9240_53877# 0.78fF
C199 a_42718_27497# a_12899_11471# 0.41fF
C200 a_2411_19605# a_4075_18543# 0.38fF
C201 a_2787_32679# a_4427_30511# 0.62fF
C202 a_48490_10496# a_48490_9492# 1.00fF
C203 a_23298_9858# a_23390_9492# 0.32fF
C204 a_4889_55535# VDD 0.43fF
C205 a_10055_58791# a_30764_7638# 0.41fF
C206 a_1923_54591# a_5291_56765# 0.35fF
C207 ctopn a_16746_9490# 1.65fF
C208 a_11067_13095# a_8295_47388# 0.37fF
C209 a_40491_27247# a_10515_23975# 0.41fF
C210 a_3339_43023# a_2411_19605# 0.41fF
C211 a_11619_56615# VDD 8.12fF
C212 a_24703_35823# VDD 0.42fF
C213 a_19720_55394# a_6775_53877# 1.13fF
C214 a_1803_20719# a_1586_36727# 1.67fF
C215 a_45478_8488# VDD 0.58fF
C216 vcm_commonmode a_36442_62194# 0.87fF
C217 a_39362_16886# a_39454_16520# 0.32fF
C218 a_32856_48463# a_32227_48169# 0.68fF
C219 a_19807_28111# a_24959_30503# 1.36fF
C220 a_16746_58180# VDD 33.19fF
C221 a_22386_59182# a_23390_59182# 0.97fF
C222 a_2944_64488# VDD 0.88fF
C223 vcm_commonmode a_44474_15516# 0.87fF
C224 ctopn a_33430_12504# 3.59fF
C225 vcm_commonmode a_23298_58178# 0.31fF
C226 a_39389_52271# a_12901_58799# 0.40fF
C227 a_29760_55394# a_29414_59182# 0.38fF
C228 a_41351_39141# VDD 1.09fF
C229 a_1823_66941# a_5291_56765# 0.63fF
C230 a_33430_72234# m3_33332_72146# 2.80fF
C231 a_4351_67279# a_11619_63151# 1.14fF
C232 a_20378_17524# a_21382_17524# 0.97fF
C233 a_16928_36391# a_15968_36061# 0.31fF
C234 a_26397_51183# a_19807_28111# 0.40fF
C235 a_8827_17215# VDD 0.58fF
C236 a_29055_49525# VDD 1.49fF
C237 vcm_commonmode a_42466_71230# 0.86fF
C238 a_5671_21495# a_10409_18543# 0.48fF
C239 a_37446_21540# a_37446_20536# 1.00fF
C240 a_2411_19605# a_1591_23445# 0.35fF
C241 a_24394_24552# a_24394_23548# 1.00fF
C242 a_33430_67214# VDD 0.51fF
C243 a_39454_12504# a_40458_12504# 0.97fF
C244 a_45386_67214# a_45478_67214# 0.32fF
C245 a_41427_52263# a_3339_43023# 0.48fF
C246 ctopn a_28410_21540# 3.59fF
C247 a_1586_45431# a_6725_45205# 0.62fF
C248 vcm_commonmode a_40366_67214# 0.31fF
C249 a_12671_37782# a_12473_37429# 0.31fF
C250 a_2497_53903# VDD 0.44fF
C251 a_21490_28585# VDD 0.31fF
C252 vcm_commonmode a_21382_13508# 0.87fF
C253 a_7571_68047# VDD 0.90fF
C254 a_8017_36495# VDD 0.39fF
C255 a_40458_68218# ctopp 3.59fF
C256 ctopn a_33430_17524# 3.59fF
C257 a_7841_12167# a_5535_18012# 0.67fF
C258 a_30418_9492# VDD 0.51fF
C259 a_25971_52263# a_30418_64202# 0.38fF
C260 a_41261_28335# a_12355_15055# 0.40fF
C261 a_46482_16520# VDD 0.51fF
C262 a_34482_29941# VDD 6.07fF
C263 a_25971_52263# a_12516_7093# 0.40fF
C264 a_32772_7638# a_32426_13508# 0.38fF
C265 a_31330_7850# a_31422_7484# 0.32fF
C266 vcm_commonmode a_37354_9858# 0.31fF
C267 a_21187_29415# a_23736_7638# 0.59fF
C268 a_44474_24552# m3_44376_24414# 2.81fF
C269 a_47486_63198# a_48490_63198# 0.97fF
C270 a_39362_72234# VDD 0.61fF
C271 vcm_commonmode a_17274_22910# 0.33fF
C272 a_28099_42895# VDD 1.68fF
C273 a_21382_18528# a_21382_17524# 1.00fF
C274 a_6646_50639# a_9963_50959# 0.91fF
C275 a_14983_51157# a_17600_50345# 0.33fF
C276 a_5877_70197# a_8485_71855# 0.74fF
C277 a_34434_21540# a_35438_21540# 0.97fF
C278 a_22291_29415# a_29175_28335# 2.04fF
C279 a_6372_38279# a_8123_34319# 0.48fF
C280 a_42374_9858# a_42466_9492# 0.32fF
C281 a_28756_7638# a_28410_22544# 0.38fF
C282 a_25306_64202# a_25398_64202# 0.32fF
C283 vcm_commonmode a_12899_10927# 6.39fF
C284 a_38450_7484# VDD 1.36fF
C285 a_22015_28111# a_26523_28111# 0.77fF
C286 a_8026_13885# VDD 0.33fF
C287 vcm_commonmode a_45478_68218# 0.87fF
C288 a_41462_59182# a_42466_59182# 0.97fF
C289 a_6559_59663# a_4891_47388# 3.33fF
C290 a_24413_39087# a_13097_37455# 0.71fF
C291 a_22294_22910# a_22386_22544# 0.32fF
C292 a_32426_64202# VDD 0.51fF
C293 a_40458_56170# ctopp 3.40fF
C294 a_5438_69679# VDD 0.35fF
C295 a_22386_14512# a_22386_13508# 1.00fF
C296 ctopn a_34434_18528# 3.59fF
C297 a_19559_41001# VDD 0.60fF
C298 a_25787_28327# a_33430_65206# 0.38fF
C299 vcm_commonmode a_39362_64202# 0.31fF
C300 a_39454_17524# a_40458_17524# 0.97fF
C301 a_11067_67279# a_16510_8760# 1.08fF
C302 a_24194_35823# a_16510_8760# 0.31fF
C303 a_22843_29415# a_19807_28111# 0.37fF
C304 a_7640_49929# VDD 0.31fF
C305 a_21382_72234# a_21382_71230# 1.00fF
C306 a_26402_60186# a_27406_60186# 0.97fF
C307 a_43470_24552# a_43470_23548# 1.00fF
C308 a_19807_28111# a_23395_32463# 0.34fF
C309 a_28410_12504# a_28410_11500# 1.00fF
C310 a_14747_31599# VDD 0.38fF
C311 vcm_commonmode a_18278_23914# 0.31fF
C312 a_17366_7484# m3_17268_7346# 2.80fF
C313 a_1683_31599# a_1849_31599# 0.52fF
C314 a_21382_18528# a_22386_18528# 0.97fF
C315 a_1803_20719# a_2007_21237# 0.60fF
C316 a_20378_19532# VDD 0.51fF
C317 a_2787_62063# VDD 0.30fF
C318 a_12641_37684# a_13669_37429# 3.30fF
C319 a_24740_7638# VDD 6.56fF
C320 a_16362_55166# m3_16264_55078# 2.81fF
C321 a_39454_61190# ctopp 3.59fF
C322 ctopn a_43470_10496# 3.59fF
C323 a_41462_69222# VDD 0.51fF
C324 a_31280_36165# VDD 1.60fF
C325 vcm_commonmode a_27314_19898# 0.31fF
C326 vcm_commonmode a_45478_56170# 0.87fF
C327 a_29760_55394# a_29414_57174# 0.38fF
C328 a_41427_52263# a_12257_56623# 0.40fF
C329 a_2235_30503# a_3339_30503# 2.22fF
C330 a_1761_34319# a_38454_34191# 0.49fF
C331 a_21187_29415# a_22291_29415# 1.08fF
C332 a_5345_47919# VDD 0.59fF
C333 a_34780_56398# a_34434_70226# 0.38fF
C334 vcm_commonmode a_48398_69222# 0.31fF
C335 a_48490_22544# VDD 0.54fF
C336 vcm_commonmode a_28410_8488# 0.86fF
C337 a_39454_65206# VDD 0.51fF
C338 a_43362_28879# a_47486_60186# 0.38fF
C339 a_36717_47375# a_10515_22671# 0.40fF
C340 a_12907_56399# a_12727_58255# 0.34fF
C341 a_18278_14878# a_18370_14512# 0.32fF
C342 a_43470_70226# ctopp 3.58fF
C343 a_1591_57711# a_1770_14441# 0.96fF
C344 vcm_commonmode a_46390_65206# 0.31fF
C345 a_34342_69222# a_34434_69222# 0.32fF
C346 a_36717_47375# a_36442_66210# 0.38fF
C347 a_40458_18528# a_40458_17524# 1.00fF
C348 a_8583_33551# a_1761_39215# 0.73fF
C349 a_1761_37039# a_1761_34319# 1.53fF
C350 a_28959_49783# a_27869_50095# 0.35fF
C351 a_24394_72234# a_25398_72234# 0.97fF
C352 a_28318_24918# VDD 0.36fF
C353 a_20359_29199# a_11067_23759# 0.98fF
C354 a_1689_10396# a_2012_33927# 0.86fF
C355 a_44382_64202# a_44474_64202# 0.32fF
C356 ctopn a_38450_15516# 3.59fF
C357 a_9529_28335# a_23051_28023# 0.47fF
C358 a_5449_25071# a_5085_24759# 1.26fF
C359 a_1761_25071# config_2_in[0] 0.93fF
C360 a_34251_52263# a_35438_62194# 0.38fF
C361 vcm_commonmode a_44474_61190# 0.87fF
C362 a_13357_32143# a_22399_32143# 1.18fF
C363 a_44474_14512# VDD 0.51fF
C364 vcm_commonmode a_12983_63151# 6.20fF
C365 a_23390_20536# VDD 0.51fF
C366 a_38358_55166# VDD 0.35fF
C367 a_41370_22910# a_41462_22544# 0.32fF
C368 a_12447_29199# a_28446_31375# 0.44fF
C369 a_6515_62037# a_4482_57863# 0.51fF
C370 a_30418_10496# a_31422_10496# 0.97fF
C371 a_36904_28879# VDD 0.63fF
C372 ctopn a_48490_11500# 3.43fF
C373 a_32334_65206# a_32426_65206# 0.32fF
C374 a_41462_14512# a_41462_13508# 1.00fF
C375 a_20827_37737# VDD 0.64fF
C376 vcm_commonmode a_30326_20902# 0.31fF
C377 a_16362_68218# ctopp 1.35fF
C378 vcm_commonmode a_19282_63198# 0.31fF
C379 a_1761_32143# a_1761_34319# 1.73fF
C380 a_27869_50095# a_12907_27023# 0.32fF
C381 a_17682_50095# a_26218_48981# 0.64fF
C382 vcm_commonmode a_48490_70226# 0.87fF
C383 a_45478_60186# a_46482_60186# 0.97fF
C384 a_49494_23548# VDD 1.14fF
C385 a_32426_58178# ctopp 3.59fF
C386 a_23298_23914# a_23390_23548# 0.32fF
C387 a_30764_7638# a_30418_21540# 0.38fF
C388 a_46482_66210# VDD 0.51fF
C389 a_2004_42453# a_2012_33927# 1.10fF
C390 a_47486_12504# a_47486_11500# 1.00fF
C391 a_12120_29941# VDD 0.42fF
C392 vcm_commonmode a_29414_16520# 0.87fF
C393 a_12725_44527# a_1761_27791# 1.27fF
C394 a_21382_72234# VDD 1.58fF
C395 a_20286_66210# a_20378_66210# 0.32fF
C396 a_18151_52263# a_12727_58255# 0.40fF
C397 a_2787_30503# a_23736_7638# 0.57fF
C398 a_23390_12504# VDD 0.51fF
C399 a_12663_40871# VDD 7.26fF
C400 a_1950_59887# a_10501_65871# 0.42fF
C401 a_34434_70226# a_34434_69222# 1.00fF
C402 a_40458_18528# a_41462_18528# 0.97fF
C403 a_25133_37571# a_12473_36341# 0.55fF
C404 vcm_commonmode a_26402_72234# 0.69fF
C405 a_3339_43023# a_4191_33449# 0.45fF
C406 vcm_commonmode a_30326_12870# 0.31fF
C407 a_20378_24552# a_21382_24552# 0.97fF
C408 a_12907_27023# a_18703_29199# 0.76fF
C409 a_32334_19898# a_32426_19532# 0.32fF
C410 a_18370_21540# VDD 0.52fF
C411 vcm_commonmode a_21382_7484# 0.69fF
C412 a_1761_40847# a_13123_38231# 1.52fF
C413 a_17366_62194# a_18370_62194# 0.97fF
C414 a_33430_11500# a_33430_10496# 1.00fF
C415 a_38436_29941# VDD 0.81fF
C416 a_25971_52263# a_15607_46805# 0.46fF
C417 a_39223_32463# a_12985_7663# 0.41fF
C418 a_16362_56170# ctopp 1.09fF
C419 a_37354_14878# a_37446_14512# 0.32fF
C420 vcm_commonmode a_25306_21906# 0.31fF
C421 a_19374_69222# ctopp 3.59fF
C422 a_3247_10389# VDD 0.44fF
C423 a_32772_7638# a_32426_7484# 0.35fF
C424 a_23390_17524# VDD 0.51fF
C425 a_39389_52271# a_39454_72234# 0.34fF
C426 a_33864_28111# a_34434_15516# 0.38fF
C427 a_3983_59887# VDD 0.31fF
C428 a_5363_30503# a_26413_31055# 0.72fF
C429 a_5254_67503# a_7107_58487# 0.42fF
C430 ctopp m3_34336_55078# 0.36fF
C431 a_28295_31287# VDD 0.38fF
C432 vcm_commonmode a_30326_17890# 0.31fF
C433 a_17366_65206# ctopp 3.43fF
C434 a_1803_19087# a_5098_41641# 0.62fF
C435 a_22386_57174# a_23390_57174# 0.97fF
C436 vcm_commonmode a_17274_60186# 0.33fF
C437 a_25398_15516# a_26402_15516# 0.97fF
C438 a_30788_28487# a_35815_31751# 0.84fF
C439 a_22291_29415# a_26523_28111# 2.32fF
C440 a_23567_44211# VDD 1.52fF
C441 a_1591_19631# VDD 0.41fF
C442 a_9507_53877# VDD 0.41fF
C443 a_35601_27497# a_35438_18528# 0.38fF
C444 a_36107_36965# VDD 0.93fF
C445 a_32823_29397# a_28841_29575# 0.73fF
C446 a_42985_46831# a_48490_58178# 0.38fF
C447 a_17599_52263# a_7479_54439# 0.65fF
C448 a_23390_71230# a_24394_71230# 0.97fF
C449 vcm_commonmode a_24394_69222# 0.87fF
C450 a_44474_59182# VDD 0.51fF
C451 a_3295_54421# a_1923_54591# 0.94fF
C452 a_6831_63303# a_2872_44111# 0.61fF
C453 a_42374_23914# a_42466_23548# 0.32fF
C454 a_35438_11500# a_36442_11500# 0.97fF
C455 a_48490_64202# ctopp 3.43fF
C456 a_14912_27497# a_11430_26159# 0.38fF
C457 a_39362_66210# a_39454_66210# 0.32fF
C458 a_7917_13885# a_8117_12559# 0.34fF
C459 vcm_commonmode a_31422_22544# 0.87fF
C460 a_5199_11791# VDD 0.36fF
C461 a_41427_52263# a_10975_66407# 0.40fF
C462 vcm_commonmode a_22386_65206# 0.87fF
C463 a_24394_18528# VDD 0.51fF
C464 a_19502_51157# VDD 0.93fF
C465 a_9135_25321# VDD 0.31fF
C466 ctopn a_22386_8488# 3.40fF
C467 a_39454_24552# a_40458_24552# 0.97fF
C468 a_1823_66941# a_3295_54421# 0.67fF
C469 vcm_commonmode a_31330_18894# 0.31fF
C470 a_24394_66210# ctopp 3.59fF
C471 a_19720_55394# a_2872_44111# 1.37fF
C472 a_1761_46287# a_12801_38517# 2.96fF
C473 a_39222_48169# a_40458_69222# 0.38fF
C474 a_17274_55166# VDD 0.37fF
C475 a_36442_62194# a_37446_62194# 0.97fF
C476 vcm_commonmode a_27406_14512# 0.87fF
C477 a_29361_38017# VDD 1.42fF
C478 a_11067_67279# a_25744_7638# 0.41fF
C479 vcm_commonmode a_22294_55166# 0.30fF
C480 a_32823_29397# a_30565_30199# 0.62fF
C481 a_33430_10496# VDD 0.51fF
C482 VDD result_out[9] 0.62fF
C483 a_3023_16341# VDD 1.83fF
C484 a_36717_47375# a_12901_66665# 0.40fF
C485 a_35346_20902# a_35438_20536# 0.32fF
C486 a_48490_60186# VDD 0.54fF
C487 vcm_commonmode a_40366_10862# 0.31fF
C488 a_9135_27239# a_21382_21540# 0.38fF
C489 a_24302_63198# a_24394_63198# 0.32fF
C490 a_11719_28023# VDD 3.14fF
C491 a_41462_57174# a_42466_57174# 0.97fF
C492 a_8531_70543# a_4758_45369# 1.07fF
C493 a_44474_15516# a_45478_15516# 0.97fF
C494 vcm_commonmode a_32426_23548# 0.87fF
C495 a_10753_12559# VDD 0.33fF
C496 a_13015_43493# VDD 0.94fF
C497 a_43470_58178# VDD 0.51fF
C498 vcm_commonmode a_29414_66210# 0.87fF
C499 a_12341_3311# a_22386_18528# 0.38fF
C500 a_32772_7638# a_12727_13353# 0.41fF
C501 a_20378_62194# VDD 0.51fF
C502 a_4351_67279# a_8491_57487# 0.55fF
C503 vcm_commonmode a_41462_19532# 0.87fF
C504 ctopn a_23390_16520# 3.59fF
C505 vcm_commonmode a_27314_62194# 0.31fF
C506 a_28410_15516# VDD 0.51fF
C507 a_21095_47919# VDD 0.42fF
C508 a_42466_71230# a_43470_71230# 0.97fF
C509 a_6559_22671# a_8933_22583# 0.67fF
C510 a_18278_59182# a_18370_59182# 0.32fF
C511 a_11067_66191# a_6559_22671# 0.38fF
C512 a_19720_7638# a_19374_19532# 0.38fF
C513 vcm_commonmode a_35346_15882# 0.31fF
C514 a_28410_63198# ctopp 3.64fF
C515 a_43269_29967# a_47486_24552# 0.55fF
C516 a_2223_28617# a_3801_24643# 0.31fF
C517 a_26402_71230# VDD 0.58fF
C518 a_28547_51175# a_12901_58799# 0.40fF
C519 a_21371_50959# a_25398_59182# 0.38fF
C520 a_5831_39189# a_8143_44982# 0.30fF
C521 a_38450_11500# VDD 0.51fF
C522 a_28980_41831# VDD 1.51fF
C523 a_32951_27247# a_33430_9492# 0.38fF
C524 a_16362_17524# a_16746_17522# 2.28fF
C525 vcm_commonmode a_33338_71230# 0.31fF
C526 a_30326_72234# a_30418_72234# 0.32fF
C527 a_9411_60437# a_9577_60437# 0.72fF
C528 a_42466_24552# VDD 0.60fF
C529 vcm_commonmode a_45386_11866# 0.31fF
C530 a_22386_59182# ctopp 3.59fF
C531 a_22386_64202# a_22386_63198# 1.23fF
C532 a_35346_12870# a_35438_12504# 0.32fF
C533 a_9307_30663# VDD 1.41fF
C534 a_4427_30511# a_4571_26677# 1.61fF
C535 a_1757_44655# VDD 0.63fF
C536 a_30418_59182# a_30418_58178# 1.00fF
C537 a_2451_72373# a_1586_69367# 1.09fF
C538 a_40086_28335# VDD 0.45fF
C539 a_44474_57174# VDD 0.51fF
C540 a_2959_47113# a_10680_52245# 0.86fF
C541 a_43267_31055# a_26523_28111# 0.42fF
C542 a_32772_7638# a_10515_23975# 0.40fF
C543 a_12663_39783# a_24029_39355# 0.57fF
C544 a_6095_44807# a_4339_64521# 1.10fF
C545 a_21382_13508# a_22386_13508# 0.97fF
C546 a_12677_36893# VDD 1.02fF
C547 vcm_commonmode a_44474_20536# 0.87fF
C548 a_2235_30503# a_9669_26703# 0.35fF
C549 a_14258_44527# a_12621_44099# 0.37fF
C550 a_2606_41079# a_1761_39215# 0.75fF
C551 a_26267_39631# VDD 0.38fF
C552 a_26402_68218# a_27406_68218# 0.97fF
C553 a_21371_52263# a_26402_64202# 0.38fF
C554 vcm_commonmode a_33430_63198# 0.92fF
C555 a_34251_52263# a_12355_15055# 0.40fF
C556 a_11067_46823# a_5039_42167# 0.93fF
C557 a_18611_52047# a_12516_7093# 8.29fF
C558 a_37919_28111# a_38450_14512# 0.38fF
C559 m3_25300_72146# VDD 0.40fF
C560 a_12355_65103# a_5039_42167# 0.57fF
C561 a_10515_23975# a_16746_22542# 0.41fF
C562 a_19967_41781# a_7841_12167# 0.42fF
C563 a_38450_56170# a_38450_55166# 1.00fF
C564 a_37446_24552# m3_37348_24414# 2.81fF
C565 a_43378_63198# a_43470_63198# 0.32fF
C566 a_34434_57174# a_34434_56170# 1.00fF
C567 a_32334_72234# VDD 0.62fF
C568 vcm_commonmode a_27406_59182# 0.87fF
C569 a_30788_28487# a_33641_29967# 0.37fF
C570 a_33694_30761# a_34759_31029# 0.33fF
C571 a_7295_44647# a_20267_30503# 3.10fF
C572 a_1761_52815# a_7078_36103# 0.45fF
C573 a_12899_10927# a_12899_11471# 23.45fF
C574 a_3891_50645# a_2595_47653# 0.34fF
C575 a_35061_51727# VDD 0.30fF
C576 a_2775_46025# a_7251_50069# 0.31fF
C577 a_31768_7638# a_12877_14441# 0.41fF
C578 a_37919_28111# a_12727_13353# 0.41fF
C579 a_30326_21906# a_30418_21540# 0.32fF
C580 a_8583_33551# a_20359_29199# 0.35fF
C581 vcm_commonmode a_44474_12504# 0.87fF
C582 a_26402_60186# ctopp 3.59fF
C583 ctopn a_45478_9492# 3.58fF
C584 a_39673_28111# a_40458_23548# 0.38fF
C585 a_29414_68218# VDD 0.51fF
C586 a_12725_44527# a_1761_41935# 0.66fF
C587 a_29322_7850# VDD 0.63fF
C588 a_48398_58178# a_48490_58178# 0.32fF
C589 a_18370_16520# a_18370_15516# 1.00fF
C590 ctopn a_25398_22544# 3.58fF
C591 a_7000_43541# a_15009_47919# 0.34fF
C592 a_4429_14191# VDD 1.25fF
C593 vcm_commonmode a_36350_68218# 0.31fF
C594 a_37354_59182# a_37446_59182# 0.32fF
C595 a_28103_38591# VDD 0.91fF
C596 vcm_commonmode a_39454_21540# 0.87fF
C597 a_10659_9813# VDD 0.38fF
C598 a_5363_30503# VDD 9.87fF
C599 a_29760_55394# a_29414_65206# 0.38fF
C600 a_35346_17890# a_35438_17524# 0.32fF
C601 a_17366_72234# a_17366_71230# 1.00fF
C602 a_30764_7638# a_12877_14441# 0.41fF
C603 a_22294_60186# a_22386_60186# 0.32fF
C604 vcm_commonmode a_16362_10496# 4.47fF
C605 a_10975_66407# a_4191_33449# 5.64fF
C606 a_4798_23759# a_5839_22351# 0.40fF
C607 a_2004_42453# a_7841_12167# 1.05fF
C608 a_41462_64202# a_41462_63198# 1.23fF
C609 vcm_commonmode a_44474_17524# 0.87fF
C610 ctopn a_21382_14512# 3.59fF
C611 a_10873_27497# a_11902_27497# 1.33fF
C612 vcm_commonmode a_31422_60186# 0.87fF
C613 a_2216_28309# a_4151_28879# 0.36fF
C614 a_43470_13508# VDD 0.51fF
C615 a_40050_48463# a_45478_68218# 0.38fF
C616 a_17274_18894# a_17366_18528# 0.32fF
C617 a_21371_52263# a_3339_30503# 0.58fF
C618 a_13669_37429# a_25517_37455# 1.22fF
C619 a_4215_51157# a_18501_50645# 0.61fF
C620 a_6467_53359# VDD 0.43fF
C621 a_33430_22544# a_33430_21540# 1.00fF
C622 a_9319_62613# VDD 0.41fF
C623 a_3305_38671# a_5963_36585# 0.36fF
C624 a_29414_56170# VDD 0.52fF
C625 a_37919_28111# a_10515_23975# 0.41fF
C626 a_40458_13508# a_41462_13508# 0.97fF
C627 a_16891_36649# VDD 0.64fF
C628 a_2021_17973# a_1803_20719# 0.91fF
C629 a_11710_58487# a_11619_63151# 0.91fF
C630 a_45478_68218# a_46482_68218# 0.97fF
C631 a_21371_50959# a_25398_57174# 0.38fF
C632 vcm_commonmode a_36350_56170# 0.31fF
C633 a_34780_56398# a_12257_56623# 0.40fF
C634 ctopn a_26402_23548# 3.40fF
C635 a_4629_13647# VDD 1.18fF
C636 a_24959_30503# VDD 10.16fF
C637 a_25971_52263# a_30418_70226# 0.38fF
C638 a_40491_27247# a_43470_14512# 0.38fF
C639 a_2177_53359# a_2007_51701# 0.31fF
C640 a_6775_53877# a_9271_52789# 0.60fF
C641 vcm_commonmode a_19282_8854# 0.31fF
C642 a_22015_28111# a_33641_29967# 0.97fF
C643 a_3247_20495# a_2011_34837# 0.63fF
C644 a_29927_29199# a_35299_32375# 0.30fF
C645 a_3339_43023# a_11067_47695# 0.75fF
C646 a_10680_52245# a_8295_47388# 0.37fF
C647 a_1823_63677# config_2_in[15] 0.51fF
C648 a_12473_42869# a_24029_39355# 0.34fF
C649 a_26402_56170# a_27406_56170# 0.97fF
C650 a_22386_57174# ctopp 3.58fF
C651 a_1761_52815# a_32971_35281# 0.46fF
C652 a_41872_29423# a_43470_60186# 0.38fF
C653 a_29760_55394# a_10515_22671# 0.40fF
C654 a_51422_39932# VDD 0.37fF
C655 ctopn a_35438_19532# 3.59fF
C656 a_28757_27247# a_30891_28309# 0.82fF
C657 a_29119_42359# VDD 0.58fF
C658 a_28547_51175# a_32426_66210# 0.38fF
C659 a_26397_51183# VDD 3.29fF
C660 a_19720_55394# a_18151_52263# 0.79fF
C661 a_49402_21906# a_49494_21540# 0.32fF
C662 a_28410_61190# VDD 0.51fF
C663 vcm_commonmode a_21382_11500# 0.87fF
C664 a_30418_58178# a_30418_57174# 1.00fF
C665 a_9301_67503# VDD 0.62fF
C666 a_4443_46607# a_12381_35836# 0.75fF
C667 vcm_commonmode a_45478_18528# 0.87fF
C668 a_28756_55394# a_28881_52271# 0.39fF
C669 vcm_commonmode a_35346_61190# 0.31fF
C670 a_31768_55394# a_31422_62194# 0.38fF
C671 a_1591_14741# a_1757_14741# 0.75fF
C672 a_37446_16520# a_37446_15516# 1.00fF
C673 vcm_commonmode a_25398_24552# 0.84fF
C674 a_40050_48463# a_45478_56170# 0.38fF
C675 a_11067_46823# a_20267_30503# 0.79fF
C676 a_32772_7638# a_32426_11500# 0.38fF
C677 a_22386_19532# a_22386_18528# 1.00fF
C678 a_24740_7638# a_24394_18528# 0.38fF
C679 a_12546_22351# a_5535_18012# 0.54fF
C680 a_26310_10862# a_26402_10496# 0.32fF
C681 a_23051_28023# VDD 0.58fF
C682 a_36442_62194# ctopp 3.59fF
C683 a_32426_70226# VDD 0.51fF
C684 vcm_commonmode a_35438_55166# 0.84fF
C685 a_30311_40229# VDD 0.90fF
C686 vcm_commonmode a_31768_7638# 10.36fF
C687 vcm_commonmode a_27406_57174# 0.87fF
C688 a_26397_51183# a_26514_47375# 0.31fF
C689 vcm_commonmode a_39362_70226# 0.31fF
C690 a_41370_60186# a_41462_60186# 0.32fF
C691 a_42718_27497# a_12985_7663# 0.41fF
C692 a_27752_7638# a_27406_19532# 0.38fF
C693 a_4674_40277# a_3607_34639# 0.89fF
C694 a_24893_37429# a_24413_39087# 0.38fF
C695 vcm_commonmode a_20286_16886# 0.31fF
C696 a_17366_15516# a_17366_14512# 1.00fF
C697 a_42466_71230# ctopp 3.40fF
C698 ctopn a_38450_20536# 3.59fF
C699 a_28446_31375# a_36507_31573# 0.30fF
C700 a_19780_41605# VDD 1.92fF
C701 a_40050_48463# a_12983_63151# 0.40fF
C702 a_36350_18894# a_36442_18528# 0.32fF
C703 a_25419_50959# VDD 17.49fF
C704 vcm_commonmode a_19374_72234# 0.69fF
C705 a_25398_61190# a_26402_61190# 0.97fF
C706 a_27937_27247# VDD 0.36fF
C707 a_12231_55509# VDD 0.36fF
C708 a_16270_24918# a_16362_24552# 0.32fF
C709 a_33963_35507# VDD 1.67fF
C710 a_43362_28879# a_12981_62313# 0.40fF
C711 vcm_commonmode a_41462_62194# 0.87fF
C712 a_31422_68218# a_31422_67214# 1.00fF
C713 vcm_commonmode a_30764_7638# 10.35fF
C714 a_21382_58178# VDD 0.51fF
C715 a_4339_64521# VDD 10.15fF
C716 a_3339_32463# a_2787_30503# 1.81fF
C717 vcm_commonmode a_49494_15516# 0.90fF
C718 ctopn a_38450_12504# 3.59fF
C719 a_45478_56170# a_46482_56170# 0.97fF
C720 vcm_commonmode a_28318_58178# 0.31fF
C721 a_2099_59861# a_2012_33927# 1.16fF
C722 a_36442_72234# m3_36344_72146# 2.80fF
C723 a_7407_46529# a_7368_46403# 0.74fF
C724 a_12901_66959# a_12727_67753# 23.56fF
C725 vcm_commonmode m2_48260_54946# 0.45fF
C726 a_22843_29415# VDD 13.34fF
C727 vcm_commonmode a_47486_71230# 0.86fF
C728 a_27314_55166# a_27406_55166# 0.32fF
C729 a_28410_8488# a_29414_8488# 0.97fF
C730 a_38450_67214# VDD 0.51fF
C731 a_23395_32463# VDD 5.57fF
C732 a_18278_57174# a_18370_57174# 0.32fF
C733 a_2361_74575# VDD 0.74fF
C734 a_21290_15882# a_21382_15516# 0.32fF
C735 ctopn a_33430_21540# 3.59fF
C736 a_30052_32117# a_28757_27247# 0.62fF
C737 a_3247_20495# VDD 9.31fF
C738 a_29414_70226# a_30418_70226# 0.97fF
C739 vcm_commonmode a_45386_67214# 0.31fF
C740 a_41462_19532# a_41462_18528# 1.00fF
C741 a_9547_54421# VDD 0.40fF
C742 a_6831_63303# a_32318_48695# 0.65fF
C743 a_6607_42167# a_3607_34639# 0.71fF
C744 a_45386_10862# a_45478_10496# 0.32fF
C745 vcm_commonmode a_26402_13508# 0.87fF
C746 a_10515_22671# a_16746_57176# 2.28fF
C747 a_45478_68218# ctopp 3.59fF
C748 ctopn a_38450_17524# 3.59fF
C749 a_1761_22895# a_1803_20719# 1.37fF
C750 a_35438_9492# VDD 0.51fF
C751 a_39299_48783# a_44474_58178# 0.38fF
C752 a_21187_29415# a_12907_27023# 1.19fF
C753 a_19282_71230# a_19374_71230# 0.32fF
C754 a_34780_56398# a_8531_70543# 0.35fF
C755 a_27406_60186# a_27406_59182# 1.00fF
C756 a_9955_21807# VDD 1.18fF
C757 vcm_commonmode a_42374_9858# 0.31fF
C758 a_33864_28111# a_34434_20536# 0.38fF
C759 a_15607_46805# a_28757_27247# 2.59fF
C760 a_12981_62313# a_16746_62196# 2.28fF
C761 a_31330_11866# a_31422_11500# 0.32fF
C762 a_12357_37999# a_13837_39860# 0.67fF
C763 a_41872_29423# VDD 8.20fF
C764 a_36442_15516# a_36442_14512# 1.00fF
C765 vcm_commonmode a_22294_22910# 0.31fF
C766 a_38784_42589# VDD 1.29fF
C767 a_34780_56398# a_10975_66407# 0.40fF
C768 a_28547_51175# a_2840_66103# 1.85fF
C769 a_13123_38231# a_1761_34319# 1.59fF
C770 vcm_commonmode a_42985_46831# 9.74fF
C771 a_44474_61190# a_45478_61190# 0.97fF
C772 a_21382_9492# a_21382_8488# 1.00fF
C773 a_11067_67279# a_9989_46831# 0.36fF
C774 a_35346_24918# a_35438_24552# 0.32fF
C775 a_25744_7638# a_25398_23548# 0.38fF
C776 a_8491_27023# a_18370_23548# 0.36fF
C777 a_3339_32463# a_7749_37903# 0.42fF
C778 a_31959_34751# VDD 0.53fF
C779 a_18662_43671# a_16152_43677# 2.10fF
C780 a_43470_7484# VDD 1.23fF
C781 a_36717_47375# a_36442_69222# 0.38fF
C782 a_33864_28111# a_34434_12504# 0.38fF
C783 a_27167_52271# a_27333_52271# 0.66fF
C784 a_37446_64202# VDD 0.51fF
C785 a_32334_62194# a_32426_62194# 0.32fF
C786 a_41334_29575# VDD 0.87fF
C787 a_9135_56623# VDD 0.71fF
C788 vcm_commonmode a_18278_14878# 0.31fF
C789 a_45478_56170# ctopp 3.40fF
C790 a_6180_69929# VDD 0.35fF
C791 ctopn a_39454_18528# 3.59fF
C792 a_27263_40871# VDD 0.53fF
C793 vcm_commonmode a_44382_64202# 0.31fF
C794 a_35438_69222# a_35438_68218# 1.00fF
C795 a_2143_15271# a_10317_13647# 0.54fF
C796 a_29760_55394# a_12901_66665# 0.40fF
C797 a_45386_55166# a_45478_55166# 0.32fF
C798 a_25398_8488# a_25398_7484# 1.00fF
C799 a_47486_8488# a_48490_8488# 0.97fF
C800 a_16362_23548# VDD 2.47fF
C801 a_37354_57174# a_37446_57174# 0.32fF
C802 a_40366_15882# a_40458_15516# 0.32fF
C803 vcm_commonmode a_23298_23914# 0.31fF
C804 a_19410_43439# VDD 1.36fF
C805 a_48490_70226# a_49494_70226# 0.97fF
C806 vcm_commonmode a_20286_66210# 0.31fF
C807 a_18370_58178# a_19374_58178# 0.97fF
C808 a_25398_19532# VDD 0.51fF
C809 a_33864_28111# a_34434_17524# 0.38fF
C810 a_44474_61190# ctopp 3.59fF
C811 ctopn a_48490_10496# 3.43fF
C812 a_12889_39889# a_1799_29556# 1.50fF
C813 a_46482_69222# VDD 0.51fF
C814 a_2944_64488# a_4339_64521# 0.61fF
C815 a_12549_35836# VDD 2.41fF
C816 vcm_commonmode a_32334_19898# 0.31fF
C817 a_12983_63151# ctopp 3.23fF
C818 a_29414_16520# a_30418_16520# 0.97fF
C819 a_6662_34025# a_7862_34025# 0.48fF
C820 a_16510_8760# a_22399_32143# 0.46fF
C821 a_38358_71230# a_38450_71230# 0.32fF
C822 a_4482_57863# a_17682_50095# 1.35fF
C823 a_4674_57685# VDD 1.31fF
C824 a_46482_60186# a_46482_59182# 1.00fF
C825 vcm_commonmode a_33430_8488# 0.86fF
C826 a_44474_65206# VDD 0.51fF
C827 a_5831_39189# a_8461_32937# 0.86fF
C828 a_35438_63198# a_35438_62194# 1.00fF
C829 a_1591_29973# VDD 0.42fF
C830 a_17507_52047# a_21382_59182# 0.38fF
C831 a_21371_50959# a_12901_58799# 0.40fF
C832 a_48490_70226# ctopp 3.42fF
C833 a_15189_39889# VDD 1.56fF
C834 a_13097_36367# a_12381_35836# 2.70fF
C835 a_9963_50959# VDD 2.54fF
C836 a_40458_9492# a_40458_8488# 1.00fF
C837 a_33338_24918# VDD 0.36fF
C838 ctopn a_43470_15516# 3.59fF
C839 a_38557_32143# a_38115_52263# 0.86fF
C840 a_12549_44212# a_12641_42036# 0.46fF
C841 a_35438_67214# a_36442_67214# 0.97fF
C842 vcm_commonmode a_49494_61190# 0.91fF
C843 a_7155_55509# a_7387_64239# 0.34fF
C844 a_5915_35943# a_15661_29199# 0.40fF
C845 a_20905_32143# a_14646_29423# 0.53fF
C846 a_2235_30503# a_16101_31029# 0.63fF
C847 a_1915_35015# a_3325_29967# 0.31fF
C848 a_12907_27023# a_26523_28111# 2.32fF
C849 a_49494_14512# VDD 1.12fF
C850 vcm_commonmode a_21382_67214# 0.87fF
C851 a_4075_18543# a_4241_18543# 0.50fF
C852 a_28410_20536# VDD 0.51fF
C853 a_43378_55166# VDD 0.35fF
C854 a_17366_63198# VDD 0.63fF
C855 a_12641_37684# a_13837_38772# 2.52fF
C856 VDD result_out[2] 0.52fF
C857 a_11067_66191# a_12869_2741# 0.47fF
C858 a_3339_43023# a_8583_33551# 27.64fF
C859 a_17274_13874# a_17366_13508# 0.32fF
C860 vcm_commonmode a_35346_20902# 0.31fF
C861 ctopn a_12877_16911# 3.23fF
C862 a_12725_44527# a_15193_44005# 0.50fF
C863 a_8423_39367# VDD 0.60fF
C864 a_28756_55394# a_12355_15055# 0.40fF
C865 a_22294_68218# a_22386_68218# 0.32fF
C866 a_17599_52263# a_22386_64202# 0.38fF
C867 vcm_commonmode a_24302_63198# 0.31fF
C868 a_3607_34639# a_3187_34293# 0.37fF
C869 a_22843_29415# a_34482_29941# 6.72fF
C870 a_20161_48463# VDD 0.41fF
C871 a_4758_45369# a_7368_46403# 0.60fF
C872 a_6361_57711# VDD 0.57fF
C873 a_21382_7484# a_22386_7484# 0.97fF
C874 a_44474_8488# a_44474_7484# 1.00fF
C875 vcm_commonmode a_18370_9492# 0.88fF
C876 a_30418_24552# m3_30320_24414# 2.81fF
C877 a_18162_31055# VDD 0.99fF
C878 vcm_commonmode a_34434_16520# 0.87fF
C879 ctopn a_20378_13508# 3.59fF
C880 a_16955_52047# a_20359_29199# 0.30fF
C881 a_9529_28335# a_17712_7638# 0.76fF
C882 a_25306_72234# VDD 0.62fF
C883 vcm_commonmode a_18278_59182# 0.31fF
C884 a_28410_12504# VDD 0.51fF
C885 a_2689_65103# a_5024_67885# 0.42fF
C886 ctopn a_28756_7638# 2.62fF
C887 a_49402_62194# VDD 0.31fF
C888 a_32426_9492# a_33430_9492# 0.97fF
C889 a_12371_53903# VDD 0.39fF
C890 vcm_commonmode a_35346_12870# 0.31fF
C891 a_33430_13508# a_33430_12504# 1.00fF
C892 a_23901_35516# VDD 1.06fF
C893 a_1768_16367# a_1823_54973# 1.14fF
C894 a_48490_16520# a_49494_16520# 0.97fF
C895 ctopn a_16362_22544# 1.33fF
C896 a_1683_33237# a_1849_33237# 0.72fF
C897 a_3063_19087# a_1895_18756# 0.45fF
C898 a_2143_15271# a_9983_18870# 0.31fF
C899 a_23390_21540# VDD 0.51fF
C900 vcm_commonmode a_26402_7484# 0.69fF
C901 a_17712_7638# a_12985_19087# 0.40fF
C902 vcm_commonmode a_30326_21906# 0.31fF
C903 a_11067_67279# a_36629_27791# 0.41fF
C904 a_24394_69222# ctopp 3.59fF
C905 a_26919_41271# VDD 0.64fF
C906 vcm_commonmode a_20378_64202# 0.87fF
C907 a_21371_50959# a_25398_65206# 0.38fF
C908 a_25971_52263# a_26523_29199# 1.64fF
C909 vcm_commonmode a_48398_58178# 0.31fF
C910 a_28410_17524# VDD 0.51fF
C911 a_49402_24918# VDD 0.47fF
C912 a_1591_23445# a_1757_23445# 0.42fF
C913 ctopp m3_48968_55078# 0.38fF
C914 a_35299_32375# VDD 1.07fF
C915 vcm_commonmode a_35346_17890# 0.31fF
C916 a_22386_65206# ctopp 3.59fF
C917 a_5345_74031# VDD 0.59fF
C918 a_23390_67214# a_23390_66210# 1.00fF
C919 vcm_commonmode a_22294_60186# 0.31fF
C920 a_7939_30503# a_6459_30511# 0.46fF
C921 a_1586_45431# a_1761_44111# 0.38fF
C922 a_24800_43041# VDD 3.97fF
C923 a_41427_52263# a_41462_68218# 0.38fF
C924 a_2143_15271# VDD 13.69fF
C925 a_6098_73095# a_7499_74031# 0.34fF
C926 a_10515_63143# a_5039_42167# 0.86fF
C927 a_43270_27791# a_45478_24552# 0.63fF
C928 a_19374_65206# a_19374_64202# 1.00fF
C929 a_4429_14191# a_5199_11791# 0.35fF
C930 a_36350_13874# a_36442_13508# 0.32fF
C931 a_1761_44111# a_13005_43983# 1.18fF
C932 a_41370_68218# a_41462_68218# 0.32fF
C933 a_17507_52047# a_21382_57174# 0.38fF
C934 a_23395_52047# a_12257_56623# 0.40fF
C935 a_5915_30287# a_14625_30761# 0.61fF
C936 a_2292_43291# a_4443_46607# 0.73fF
C937 a_20359_29199# a_15607_46805# 9.40fF
C938 a_7959_15279# VDD 0.41fF
C939 a_24209_48463# VDD 0.42fF
C940 vcm_commonmode a_29414_69222# 0.87fF
C941 a_21371_52263# a_26402_70226# 0.38fF
C942 a_43175_28335# a_46482_13508# 0.38fF
C943 a_49494_59182# VDD 1.22fF
C944 a_40458_7484# a_41462_7484# 0.97fF
C945 a_3016_60949# a_3325_49551# 0.30fF
C946 a_29760_55394# a_19807_28111# 0.83fF
C947 a_11602_25071# a_12707_26159# 0.46fF
C948 a_28817_29111# a_17712_7638# 0.52fF
C949 a_22294_56170# a_22386_56170# 0.32fF
C950 a_17599_52263# a_10515_22671# 0.40fF
C951 a_39389_52271# a_39454_60186# 0.38fF
C952 vcm_commonmode a_36442_22544# 0.87fF
C953 a_28756_55394# a_28410_66210# 0.38fF
C954 a_24394_69222# a_25398_69222# 0.97fF
C955 vcm_commonmode a_27406_65206# 0.87fF
C956 a_6883_37019# a_3607_34639# 0.70fF
C957 a_29414_18528# VDD 0.51fF
C958 a_24683_51183# VDD 0.44fF
C959 a_17366_72234# a_18370_72234# 0.97fF
C960 a_11251_59879# a_12683_51329# 0.43fF
C961 a_12641_37684# a_13005_35823# 1.90fF
C962 a_19374_61190# a_19374_60186# 1.00fF
C963 a_2007_23957# VDD 0.43fF
C964 ctopn a_27406_8488# 3.40fF
C965 a_8491_41383# a_5915_35943# 2.89fF
C966 a_34434_64202# a_35438_64202# 0.97fF
C967 a_26661_34428# VDD 0.84fF
C968 a_10055_58791# a_11067_23759# 0.34fF
C969 vcm_commonmode a_36350_18894# 0.31fF
C970 a_29414_66210# ctopp 3.59fF
C971 a_17507_52047# a_28881_52271# 0.33fF
C972 a_23928_28585# a_23192_27791# 0.87fF
C973 a_23395_52047# a_27406_62194# 0.38fF
C974 vcm_commonmode a_16270_24918# 0.33fF
C975 a_41427_52263# a_41462_56170# 0.38fF
C976 a_2235_30503# a_14926_31849# 1.10fF
C977 a_6224_73095# a_6515_67477# 0.47fF
C978 a_20378_55166# VDD 0.60fF
C979 a_31422_22544# a_32426_22544# 0.97fF
C980 a_31768_7638# a_12899_11471# 0.41fF
C981 a_9424_60949# a_7210_55081# 0.30fF
C982 vcm_commonmode a_32426_14512# 0.87fF
C983 a_17488_48731# a_7841_12167# 2.26fF
C984 a_22386_65206# a_23390_65206# 0.97fF
C985 a_37733_37477# VDD 1.81fF
C986 vcm_commonmode a_27314_55166# 0.30fF
C987 a_38450_10496# VDD 0.51fF
C988 a_18370_17524# a_18370_16520# 1.00fF
C989 vcm_commonmode a_18278_57174# 0.31fF
C990 a_36464_49783# VDD 0.34fF
C991 a_1950_59887# a_5682_69367# 0.63fF
C992 vcm_commonmode a_45386_10862# 0.31fF
C993 a_22386_56170# a_22386_55166# 1.00fF
C994 a_3016_60949# a_5252_56891# 0.60fF
C995 a_21371_50959# a_27869_50095# 0.35fF
C996 a_42466_67214# a_42466_66210# 1.00fF
C997 vcm_commonmode a_37446_23548# 0.87fF
C998 a_10055_58791# a_16362_12504# 1.27fF
C999 vcm_commonmode a_34434_66210# 0.87fF
C1000 a_38557_32143# a_12983_63151# 0.40fF
C1001 a_15505_52521# VDD 0.38fF
C1002 a_1923_73087# a_4719_71855# 0.57fF
C1003 a_36797_27497# a_12877_16911# 0.41fF
C1004 a_30764_7638# a_12899_11471# 0.41fF
C1005 a_25398_62194# VDD 0.51fF
C1006 a_21290_61190# a_21382_61190# 0.32fF
C1007 a_38450_65206# a_38450_64202# 1.00fF
C1008 vcm_commonmode a_46482_19532# 0.87fF
C1009 ctopn a_28410_16520# 3.59fF
C1010 vcm_commonmode a_32334_62194# 0.31fF
C1011 a_39222_48169# a_12981_62313# 0.40fF
C1012 a_33430_15516# VDD 0.51fF
C1013 a_22386_19532# a_23390_19532# 0.97fF
C1014 a_39223_32463# a_39454_8488# 0.38fF
C1015 a_10590_21263# VDD 0.59fF
C1016 a_32426_23548# a_32426_22544# 1.00fF
C1017 a_6138_54599# a_6236_54421# 0.30fF
C1018 vcm_commonmode a_40366_15882# 0.31fF
C1019 a_33430_63198# ctopp 3.64fF
C1020 a_41370_56170# a_41462_56170# 0.32fF
C1021 a_31422_71230# VDD 0.58fF
C1022 a_26402_66210# a_26402_65206# 1.00fF
C1023 a_27406_14512# a_28410_14512# 0.97fF
C1024 a_32029_38565# VDD 1.98fF
C1025 a_11067_13095# a_5449_25071# 0.63fF
C1026 a_43470_11500# VDD 0.51fF
C1027 a_33727_42089# VDD 0.64fF
C1028 a_43470_69222# a_44474_69222# 0.97fF
C1029 a_13097_35279# a_14735_35805# 0.34fF
C1030 a_2596_16911# VDD 0.43fF
C1031 vcm_commonmode a_38358_71230# 0.31fF
C1032 a_28547_51175# a_32426_72234# 0.35fF
C1033 a_38450_61190# a_38450_60186# 1.00fF
C1034 a_7210_55081# a_8199_58229# 0.37fF
C1035 a_24302_8854# a_24394_8488# 0.32fF
C1036 a_47486_24552# VDD 0.58fF
C1037 a_27406_59182# ctopp 3.59fF
C1038 a_27535_30503# a_31964_30485# 0.32fF
C1039 a_12631_28585# a_14471_28585# 0.50fF
C1040 a_16746_15514# a_12877_14441# 2.28fF
C1041 a_23395_32463# a_28295_31287# 0.35fF
C1042 a_1586_45431# a_4842_45467# 0.31fF
C1043 a_25306_70226# a_25398_70226# 0.32fF
C1044 a_41261_28335# a_12727_67753# 0.40fF
C1045 a_2339_38129# a_3143_22364# 0.35fF
C1046 a_42374_58178# a_42466_58178# 0.32fF
C1047 a_35601_27497# a_12899_10927# 0.41fF
C1048 a_7295_44647# a_17554_30663# 0.39fF
C1049 a_24394_62194# a_24394_61190# 1.00fF
C1050 a_49494_57174# VDD 1.10fF
C1051 vcm_commonmode a_17274_13874# 0.33fF
C1052 a_3325_18543# a_2411_19605# 0.77fF
C1053 a_41462_65206# a_42466_65206# 0.97fF
C1054 vcm_commonmode a_49494_20536# 0.90fF
C1055 a_35739_39679# VDD 0.94fF
C1056 vcm_commonmode a_38450_63198# 0.92fF
C1057 a_37446_17524# a_37446_16520# 1.00fF
C1058 a_22015_28111# a_16863_29415# 7.37fF
C1059 a_17507_52047# a_4351_67279# 0.44fF
C1060 a_24394_20536# a_24394_19532# 1.00fF
C1061 a_28756_7638# a_28410_13508# 0.38fF
C1062 a_39673_28111# a_40458_14512# 0.38fF
C1063 a_12341_3311# a_5535_18012# 0.43fF
C1064 a_32426_23548# a_33430_23548# 0.97fF
C1065 a_12357_37999# a_12889_39889# 0.36fF
C1066 a_36717_47375# VDD 6.91fF
C1067 vcm_commonmode a_32426_59182# 0.87fF
C1068 a_29414_66210# a_30418_66210# 0.97fF
C1069 a_12985_19087# a_16746_9490# 2.28fF
C1070 a_3339_30503# a_6752_29941# 0.37fF
C1071 vcm_commonmode m3_16264_66122# 3.21fF
C1072 a_23395_52047# a_10975_66407# 0.40fF
C1073 vcm_commonmode a_41427_52263# 10.02fF
C1074 a_12355_15055# a_8491_41383# 1.82fF
C1075 a_2775_46025# a_17682_50095# 1.20fF
C1076 a_2959_47113# VDD 18.90fF
C1077 a_3339_43023# a_2606_41079# 1.31fF
C1078 a_40366_61190# a_40458_61190# 0.32fF
C1079 vcm_commonmode a_49494_12504# 0.90fF
C1080 a_31422_60186# ctopp 3.59fF
C1081 a_34434_68218# VDD 0.51fF
C1082 a_10975_66407# a_8491_27023# 2.39fF
C1083 a_34342_7850# VDD 0.62fF
C1084 a_19410_43439# a_12663_40871# 1.71fF
C1085 a_24800_43041# a_28099_42895# 0.57fF
C1086 a_43267_31055# a_46482_63198# 0.42fF
C1087 ctopn a_30418_22544# 3.58fF
C1088 a_27535_30503# a_12447_29199# 0.43fF
C1089 a_5039_42167# a_7571_26151# 1.97fF
C1090 a_28547_51175# a_32426_69222# 0.38fF
C1091 a_29414_71230# a_29414_70226# 1.00fF
C1092 a_5682_69367# a_2952_66139# 0.51fF
C1093 a_39299_48783# a_12901_66959# 0.40fF
C1094 vcm_commonmode a_41370_68218# 0.31fF
C1095 a_41462_19532# a_42466_19532# 0.97fF
C1096 a_29760_7638# a_29414_19532# 0.38fF
C1097 a_23736_7638# a_12727_15529# 0.41fF
C1098 a_10055_58791# a_27752_7638# 0.41fF
C1099 a_12801_38517# a_12663_39783# 0.77fF
C1100 a_5208_70063# VDD 1.27fF
C1101 a_45478_66210# a_45478_65206# 1.00fF
C1102 a_46482_14512# a_47486_14512# 0.97fF
C1103 a_39799_38825# VDD 0.63fF
C1104 vcm_commonmode a_44474_21540# 0.87fF
C1105 a_6459_30511# a_12340_29967# 0.39fF
C1106 a_28757_27247# a_28841_29575# 0.66fF
C1107 a_43175_28335# a_46482_7484# 0.34fF
C1108 a_43267_31055# a_43362_28879# 3.67fF
C1109 a_17599_52263# a_12901_66665# 0.40fF
C1110 a_4482_57863# a_29361_51727# 0.47fF
C1111 a_25398_20536# a_26402_20536# 0.97fF
C1112 a_43378_8854# a_43470_8488# 0.32fF
C1113 vcm_commonmode a_21382_10496# 0.87fF
C1114 a_1768_16367# VDD 6.28fF
C1115 vcm_commonmode a_49494_17524# 0.91fF
C1116 ctopn a_26402_14512# 3.59fF
C1117 a_12263_4391# a_10964_25615# 0.82fF
C1118 a_12713_43011# a_12473_41781# 2.05fF
C1119 a_9353_72399# VDD 0.95fF
C1120 vcm_commonmode a_36442_60186# 0.87fF
C1121 a_30052_32117# a_28446_31375# 0.33fF
C1122 a_48490_13508# VDD 0.54fF
C1123 a_44382_70226# a_44474_70226# 0.32fF
C1124 a_32772_7638# a_32426_10496# 0.38fF
C1125 a_14983_51157# a_13445_50639# 0.79fF
C1126 a_16362_19532# VDD 2.47fF
C1127 a_6831_63303# a_26218_48981# 0.62fF
C1128 a_43470_62194# a_43470_61190# 1.00fF
C1129 a_34434_10496# a_34434_9492# 1.00fF
C1130 a_34434_56170# VDD 0.52fF
C1131 a_26748_7638# a_26402_23548# 0.38fF
C1132 a_31768_55394# a_31422_55166# 0.46fF
C1133 a_17366_8488# VDD 0.64fF
C1134 a_3339_43023# a_5595_33205# 1.66fF
C1135 a_4351_67279# a_11067_13095# 0.44fF
C1136 a_25306_16886# a_25398_16520# 0.32fF
C1137 vcm_commonmode a_41370_56170# 0.31fF
C1138 ctopn a_31422_23548# 3.40fF
C1139 a_38067_47349# VDD 0.62fF
C1140 a_43470_20536# a_43470_19532# 1.00fF
C1141 vcm_commonmode a_24302_8854# 0.31fF
C1142 vcm_commonmode a_16746_15514# 5.36fF
C1143 a_11067_63143# a_3339_43023# 0.83fF
C1144 a_27406_57174# ctopp 3.58fF
C1145 a_48490_66210# a_49494_66210# 0.97fF
C1146 a_14287_51175# a_12901_58799# 0.40fF
C1147 ctopn a_40458_19532# 3.59fF
C1148 vcm_commonmode m3_16264_13370# 3.21fF
C1149 a_2235_30503# a_22577_29111# 0.45fF
C1150 a_28757_27247# a_30565_30199# 0.48fF
C1151 a_42985_46831# a_12355_65103# 0.40fF
C1152 a_23298_72234# a_23390_72234# 0.32fF
C1153 a_23390_21540# a_23390_20536# 1.00fF
C1154 a_30764_7638# a_30418_16520# 0.38fF
C1155 a_33430_61190# VDD 0.51fF
C1156 vcm_commonmode a_26402_11500# 0.87fF
C1157 a_41872_29423# a_43470_58178# 0.38fF
C1158 a_4443_46607# a_1761_35407# 0.48fF
C1159 a_25398_12504# a_26402_12504# 0.97fF
C1160 a_1849_33237# VDD 0.62fF
C1161 a_36392_43677# a_32327_40191# 0.54fF
C1162 a_31330_67214# a_31422_67214# 0.32fF
C1163 vcm_commonmode a_40366_61190# 0.31fF
C1164 vcm_commonmode a_30418_24552# 0.84fF
C1165 a_3983_45743# VDD 0.46fF
C1166 a_48490_71230# a_48490_70226# 1.00fF
C1167 a_8295_47388# VDD 13.32fF
C1168 a_4075_63151# VDD 0.33fF
C1169 a_13643_28327# a_9529_28335# 0.67fF
C1170 a_41462_62194# ctopp 3.59fF
C1171 a_18151_52263# a_4674_40277# 4.10fF
C1172 a_39222_48169# a_37557_32463# 0.91fF
C1173 a_37446_70226# VDD 0.51fF
C1174 vcm_commonmode a_40458_55166# 0.84fF
C1175 a_51714_39886# VDD 0.57fF
C1176 a_14287_51175# a_18370_64202# 0.38fF
C1177 a_17507_52047# a_12355_15055# 0.40fF
C1178 vcm_commonmode a_32426_57174# 0.87fF
C1179 a_18370_16520# VDD 0.52fF
C1180 vcm_commonmode a_44382_70226# 0.31fF
C1181 a_44474_20536# a_45478_20536# 0.97fF
C1182 a_17274_7850# a_17366_7484# 0.32fF
C1183 a_39223_32463# a_12727_13353# 0.41fF
C1184 VDD config_1_in[1] 0.89fF
C1185 a_23390_24552# m3_23292_24414# 2.81fF
C1186 a_33430_63198# a_34434_63198# 0.97fF
C1187 vcm_commonmode a_25306_16886# 0.31fF
C1188 a_13576_42589# a_12641_42036# 3.10fF
C1189 a_18278_72234# VDD 0.62fF
C1190 ctopp m2_48260_54946# 1.14fF
C1191 a_47486_71230# ctopp 3.39fF
C1192 ctopn a_43470_20536# 3.59fF
C1193 a_30679_43493# VDD 1.05fF
C1194 a_33338_58178# a_33430_58178# 0.32fF
C1195 a_25133_37571# a_1761_30511# 1.57fF
C1196 a_6559_59879# a_11711_50645# 0.63fF
C1197 a_20378_21540# a_21382_21540# 0.97fF
C1198 a_22015_28111# a_19720_7638# 0.37fF
C1199 a_28318_9858# a_28410_9492# 0.32fF
C1200 a_17712_7638# VDD 7.53fF
C1201 a_4035_54965# VDD 0.38fF
C1202 a_10055_58791# a_8491_27023# 0.42fF
C1203 a_12549_44212# a_16152_43677# 1.75fF
C1204 vcm_commonmode a_46482_62194# 0.87fF
C1205 a_44382_16886# a_44474_16520# 0.32fF
C1206 a_7841_12167# a_10873_27497# 0.46fF
C1207 a_16863_29415# a_22291_29415# 1.15fF
C1208 vcm_commonmode a_17366_68218# 1.83fF
C1209 a_2419_48783# a_1586_45431# 0.31fF
C1210 a_26402_58178# VDD 0.51fF
C1211 a_27406_59182# a_28410_59182# 0.97fF
C1212 a_13669_38517# a_15305_38543# 0.43fF
C1213 a_2840_66103# a_2419_48783# 0.45fF
C1214 a_11067_67279# a_16746_19530# 0.41fF
C1215 ctopn a_43470_12504# 3.59fF
C1216 vcm_commonmode a_33338_58178# 0.31fF
C1217 a_75199_38962# VDD 0.44fF
C1218 a_39454_72234# m3_39356_72146# 2.80fF
C1219 a_15775_41317# VDD 1.00fF
C1220 a_17507_52047# a_21382_65206# 0.38fF
C1221 VDD config_2_in[2] 0.97fF
C1222 a_28756_7638# a_28410_7484# 0.35fF
C1223 a_25398_17524# a_26402_17524# 0.97fF
C1224 a_2011_34837# a_1915_35015# 1.99fF
C1225 a_25419_50959# a_24959_30503# 1.42fF
C1226 a_42466_21540# a_42466_20536# 1.00fF
C1227 a_2191_68565# a_1761_25071# 0.69fF
C1228 a_29414_24552# a_29414_23548# 1.00fF
C1229 a_43470_67214# VDD 0.51fF
C1230 a_44474_12504# a_45478_12504# 0.97fF
C1231 a_14646_29423# VDD 4.28fF
C1232 a_39223_32463# a_10515_23975# 0.41fF
C1233 a_42985_46831# ctopp 2.48fF
C1234 ctopn a_38450_21540# 3.59fF
C1235 a_17488_48731# a_5831_39189# 0.49fF
C1236 a_4443_46607# a_3339_32463# 2.62fF
C1237 a_18703_29199# a_18979_30287# 1.92fF
C1238 a_19096_44129# VDD 1.53fF
C1239 a_36613_48169# a_37446_68218# 0.38fF
C1240 a_12473_37429# a_13669_37429# 0.82fF
C1241 VDD config_2_in[11] 1.06fF
C1242 a_1823_53885# VDD 1.55fF
C1243 a_21187_29415# a_30975_28023# 0.39fF
C1244 a_22291_29415# a_23685_29111# 0.32fF
C1245 a_13643_28327# a_28817_29111# 0.77fF
C1246 vcm_commonmode a_31422_13508# 0.87fF
C1247 a_11067_13095# a_12355_15055# 0.69fF
C1248 a_27183_36965# VDD 1.02fF
C1249 ctopn a_43470_17524# 3.59fF
C1250 a_40458_9492# VDD 0.51fF
C1251 a_16955_52047# a_12257_56623# 0.40fF
C1252 vcm_commonmode a_17366_56170# 1.83fF
C1253 vcm_commonmode a_20286_69222# 0.31fF
C1254 a_17599_52263# a_22386_70226# 0.38fF
C1255 a_25744_7638# a_25398_14512# 0.38fF
C1256 a_8491_27023# a_18370_14512# 0.38fF
C1257 a_36350_7850# a_36442_7484# 0.32fF
C1258 a_20378_22544# VDD 0.51fF
C1259 vcm_commonmode a_47394_9858# 0.31fF
C1260 a_24959_30503# a_23395_32463# 2.64fF
C1261 a_11183_30761# VDD 0.55fF
C1262 a_17599_52263# a_19807_28111# 0.56fF
C1263 a_11619_56615# a_8295_47388# 3.25fF
C1264 a_34251_52263# a_35438_60186# 0.38fF
C1265 a_3024_67191# a_9643_63125# 0.39fF
C1266 a_4812_13879# a_5227_13621# 0.52fF
C1267 vcm_commonmode a_27314_22910# 0.31fF
C1268 ctopn a_12895_13967# 3.23fF
C1269 a_3247_20495# a_4629_13647# 0.44fF
C1270 a_2235_41941# VDD 0.50fF
C1271 a_18151_52263# a_24394_66210# 0.38fF
C1272 a_20286_69222# a_20378_69222# 0.32fF
C1273 vcm_commonmode a_18278_65206# 0.31fF
C1274 a_26402_18528# a_26402_17524# 1.00fF
C1275 a_1761_30511# a_12473_36341# 1.91fF
C1276 a_39454_21540# a_40458_21540# 0.97fF
C1277 a_9135_27239# a_21382_16520# 0.38fF
C1278 a_47394_9858# a_47486_9492# 0.32fF
C1279 a_9260_25045# VDD 0.56fF
C1280 a_30326_64202# a_30418_64202# 0.32fF
C1281 a_48490_7484# VDD 1.28fF
C1282 vcm_commonmode a_12981_59343# 6.23fF
C1283 a_18611_52047# a_23390_62194# 0.38fF
C1284 a_36613_48169# a_37446_56170# 0.38fF
C1285 a_34482_29941# a_38067_47349# 0.32fF
C1286 a_16362_14512# VDD 2.47fF
C1287 a_46482_59182# a_47486_59182# 0.97fF
C1288 a_27314_22910# a_27406_22544# 0.32fF
C1289 a_42466_64202# VDD 0.51fF
C1290 a_3305_38671# a_6786_37557# 0.73fF
C1291 a_2589_55535# VDD 0.79fF
C1292 vcm_commonmode a_23298_14878# 0.31fF
C1293 ctopn a_20378_11500# 3.59fF
C1294 a_18278_65206# a_18370_65206# 0.32fF
C1295 a_27406_14512# a_27406_13508# 1.00fF
C1296 a_11067_67279# a_29760_7638# 0.41fF
C1297 ctopn a_44474_18528# 3.59fF
C1298 a_75794_40594# VDD 0.83fF
C1299 a_3024_67191# a_8772_63927# 0.57fF
C1300 vcm_commonmode a_49402_64202# 0.30fF
C1301 a_44474_17524# a_45478_17524# 0.97fF
C1302 vcm_commonmode a_20378_70226# 0.87fF
C1303 a_37446_58178# vcm_commonmode 0.87fF
C1304 a_6559_22671# a_4528_26159# 1.62fF
C1305 a_31422_60186# a_32426_60186# 0.97fF
C1306 a_21382_23548# VDD 0.52fF
C1307 a_10515_22671# a_7841_22895# 0.42fF
C1308 a_4891_47388# a_12659_54965# 2.00fF
C1309 a_33864_28111# a_34434_21540# 0.38fF
C1310 a_18370_66210# VDD 0.52fF
C1311 a_33430_12504# a_33430_11500# 1.00fF
C1312 vcm_commonmode a_28318_23914# 0.31fF
C1313 a_1761_49007# a_14258_44527# 2.21fF
C1314 a_35463_44031# VDD 0.83fF
C1315 a_31768_55394# a_12983_63151# 0.40fF
C1316 a_20378_70226# a_20378_69222# 1.00fF
C1317 vcm_commonmode a_25306_66210# 0.31fF
C1318 a_26402_18528# a_27406_18528# 0.97fF
C1319 a_25419_50959# a_22843_29415# 0.82fF
C1320 a_30418_19532# VDD 0.51fF
C1321 a_13643_28327# a_37699_27221# 0.44fF
C1322 a_12981_59343# a_16362_61190# 19.89fF
C1323 a_25419_50959# a_23395_32463# 0.39fF
C1324 a_1915_35015# VDD 4.79fF
C1325 vcm_commonmode a_37354_19898# 0.31fF
C1326 a_21382_67214# ctopp 3.59fF
C1327 a_13716_43047# a_12357_37999# 0.40fF
C1328 a_25787_28327# a_12981_62313# 0.40fF
C1329 a_2143_15271# a_10753_12559# 0.40fF
C1330 a_19439_47919# VDD 0.40fF
C1331 a_13183_52047# a_12901_66959# 0.40fF
C1332 a_18278_19898# a_18370_19532# 0.32fF
C1333 vcm_commonmode a_38450_8488# 0.86fF
C1334 a_49494_65206# VDD 1.12fF
C1335 a_19807_28111# a_30790_30663# 0.58fF
C1336 a_19374_11500# a_19374_10496# 1.00fF
C1337 a_4248_29967# VDD 2.90fF
C1338 a_3949_41935# a_4685_37583# 1.56fF
C1339 a_23298_14878# a_23390_14512# 0.32fF
C1340 a_5831_39189# a_1761_25071# 0.39fF
C1341 a_21663_41855# VDD 0.88fF
C1342 a_39362_69222# a_39454_69222# 0.32fF
C1343 a_45478_18528# a_45478_17524# 1.00fF
C1344 a_39673_28111# a_12727_15529# 0.41fF
C1345 a_38358_24918# VDD 0.36fF
C1346 a_49402_64202# a_49494_64202# 0.32fF
C1347 a_2235_31055# VDD 0.48fF
C1348 ctopn a_48490_15516# 3.43fF
C1349 a_1803_19087# a_2411_26133# 1.05fF
C1350 a_3024_67191# a_5595_63125# 0.79fF
C1351 a_7815_45503# VDD 0.60fF
C1352 vcm_commonmode a_26402_67214# 0.87fF
C1353 a_34251_52263# a_12727_67753# 0.40fF
C1354 a_43175_28335# a_46482_11500# 0.38fF
C1355 a_33430_20536# VDD 0.51fF
C1356 a_49402_55166# VDD 0.48fF
C1357 a_2775_46025# a_29361_51727# 0.41fF
C1358 a_46390_22910# a_46482_22544# 0.32fF
C1359 a_26748_7638# a_12877_16911# 0.41fF
C1360 a_22386_63198# VDD 0.57fF
C1361 a_12641_37684# a_13909_38659# 0.96fF
C1362 a_35438_10496# a_36442_10496# 0.97fF
C1363 a_12263_4391# a_11067_21583# 1.62fF
C1364 a_37354_65206# a_37446_65206# 0.32fF
C1365 a_10975_66407# a_11067_63143# 2.55fF
C1366 a_46482_14512# a_46482_13508# 1.00fF
C1367 a_34699_37683# VDD 1.33fF
C1368 vcm_commonmode a_40366_20902# 0.31fF
C1369 a_16746_9490# VDD 33.20fF
C1370 vcm_commonmode a_29322_63198# 0.31fF
C1371 a_17039_51157# a_7571_29199# 0.62fF
C1372 a_16746_59184# VDD 33.20fF
C1373 a_4674_40277# a_5211_24759# 0.40fF
C1374 vcm_commonmode a_23390_9492# 0.87fF
C1375 a_11067_23759# a_12877_14441# 0.35fF
C1376 a_28318_23914# a_28410_23548# 0.32fF
C1377 a_19807_28111# a_19626_31751# 2.33fF
C1378 a_8491_41383# a_4811_34855# 0.52fF
C1379 a_21382_11500# a_22386_11500# 0.97fF
C1380 a_29667_31055# VDD 0.30fF
C1381 vcm_commonmode a_39454_16520# 0.87fF
C1382 a_20378_64202# ctopp 3.59fF
C1383 ctopn a_25398_13508# 3.59fF
C1384 a_29760_55394# VDD 7.20fF
C1385 vcm_commonmode a_23298_59182# 0.31fF
C1386 a_25306_66210# a_25398_66210# 0.32fF
C1387 a_2411_18517# a_11179_9981# 0.36fF
C1388 a_33430_12504# VDD 0.51fF
C1389 a_39454_70226# a_39454_69222# 1.00fF
C1390 a_14287_51175# a_2840_66103# 0.33fF
C1391 a_16955_52047# a_10975_66407# 0.40fF
C1392 a_45478_18528# a_46482_18528# 0.97fF
C1393 vcm_commonmode a_34780_56398# 10.02fF
C1394 a_3295_62083# a_6559_59663# 0.44fF
C1395 vcm_commonmode a_40366_12870# 0.31fF
C1396 a_25398_24552# a_26402_24552# 0.97fF
C1397 a_29127_35561# VDD 0.63fF
C1398 a_41261_28335# a_42466_63198# 0.42fF
C1399 a_2004_42453# a_3063_19087# 0.64fF
C1400 a_1591_14191# VDD 0.43fF
C1401 a_13413_47375# VDD 0.62fF
C1402 a_28756_55394# a_28410_69222# 0.38fF
C1403 a_36613_48169# a_12901_66959# 0.40fF
C1404 a_1586_9991# a_4075_18543# 0.44fF
C1405 a_37354_19898# a_37446_19532# 0.32fF
C1406 a_28410_21540# VDD 0.51fF
C1407 vcm_commonmode a_31422_7484# 0.69fF
C1408 config_2_in[1] rst_n 0.53fF
C1409 a_36797_27497# a_12895_13967# 0.41fF
C1410 a_3339_43023# a_1586_9991# 0.78fF
C1411 a_4314_40821# a_5915_35943# 0.40fF
C1412 a_2787_32679# a_5993_32687# 1.06fF
C1413 a_22386_62194# a_23390_62194# 0.97fF
C1414 a_38450_11500# a_38450_10496# 1.00fF
C1415 a_46482_58178# VDD 0.51fF
C1416 a_43362_28879# a_12907_27023# 0.35fF
C1417 a_42374_14878# a_42466_14512# 0.32fF
C1418 vcm_commonmode a_35346_21906# 0.31fF
C1419 a_29414_69222# ctopp 3.59fF
C1420 vcm_commonmode a_25398_64202# 0.87fF
C1421 a_2411_18517# a_8123_14741# 0.39fF
C1422 a_12381_35836# a_1761_32143# 1.45fF
C1423 a_33430_17524# VDD 0.51fF
C1424 a_29147_50069# VDD 0.38fF
C1425 a_42466_72234# a_43470_72234# 0.97fF
C1426 a_21290_20902# a_21382_20536# 0.32fF
C1427 a_20378_60186# VDD 0.51fF
C1428 a_35438_55166# a_36442_55166# 0.97fF
C1429 a_41967_31375# a_12899_10927# 0.41fF
C1430 vcm_commonmode a_40366_17890# 0.31fF
C1431 a_27406_65206# ctopp 3.59fF
C1432 a_27406_57174# a_28410_57174# 0.97fF
C1433 a_10055_74031# VDD 0.49fF
C1434 vcm_commonmode a_27314_60186# 0.31fF
C1435 a_30418_15516# a_31422_15516# 0.97fF
C1436 a_49494_8488# m3_49396_8350# 2.78fF
C1437 a_7939_30503# a_22151_29941# 0.34fF
C1438 a_33819_44535# VDD 0.59fF
C1439 a_3325_69135# a_4307_67477# 0.81fF
C1440 a_14293_37455# a_17585_37477# 0.54fF
C1441 a_4312_19061# VDD 0.32fF
C1442 a_4792_20443# a_5535_18012# 1.02fF
C1443 a_7803_55509# a_7764_53877# 0.79fF
C1444 a_9503_26151# a_20378_24552# 0.46fF
C1445 a_7215_36201# VDD 0.67fF
C1446 a_23395_52047# a_27406_55166# 0.47fF
C1447 a_1761_22895# a_13067_38517# 1.00fF
C1448 a_34251_52263# a_12899_2767# 0.53fF
C1449 a_16587_49007# a_16753_49007# 0.69fF
C1450 vcm_commonmode a_34434_69222# 0.87fF
C1451 a_28410_71230# a_29414_71230# 0.97fF
C1452 a_2099_59861# a_1923_54591# 2.17fF
C1453 vcm_commonmode a_12947_8725# 4.77fF
C1454 a_47394_23914# a_47486_23548# 0.32fF
C1455 a_2411_26133# a_2971_37589# 0.36fF
C1456 a_40458_11500# a_41462_11500# 0.97fF
C1457 a_44382_66210# a_44474_66210# 0.32fF
C1458 a_11067_66191# a_11067_13095# 1.55fF
C1459 vcm_commonmode a_41462_22544# 0.87fF
C1460 a_5831_39189# a_2787_32679# 0.83fF
C1461 a_9455_11079# VDD 0.38fF
C1462 a_41427_52263# a_12355_65103# 0.40fF
C1463 vcm_commonmode a_32426_65206# 0.87fF
C1464 a_34434_18528# VDD 0.51fF
C1465 a_42718_27497# a_12727_13353# 0.41fF
C1466 vcm_commonmode a_17274_11866# 0.33fF
C1467 ctopn a_32426_8488# 3.40fF
C1468 a_19720_7638# a_19374_22544# 0.38fF
C1469 a_31768_7638# a_12985_7663# 0.41fF
C1470 a_44474_24552# a_45478_24552# 0.97fF
C1471 a_22015_28111# a_2235_30503# 0.49fF
C1472 a_21290_12870# a_21382_12504# 0.32fF
C1473 vcm_commonmode a_41370_18894# 0.31fF
C1474 a_34434_66210# ctopp 3.59fF
C1475 a_14287_51175# a_12755_51562# 0.31fF
C1476 a_23192_27791# a_27752_7638# 0.56fF
C1477 vcm_commonmode a_21290_24918# 0.31fF
C1478 a_1761_52815# a_2411_26133# 0.71fF
C1479 a_1761_46287# VDD 5.94fF
C1480 a_28756_7638# a_28410_11500# 0.38fF
C1481 vcm_commonmode a_11067_23759# 5.78fF
C1482 a_12901_58799# a_16362_58178# 1.15fF
C1483 a_7933_51433# a_8051_52047# 0.39fF
C1484 a_8625_20175# VDD 0.60fF
C1485 a_25398_55166# VDD 0.60fF
C1486 a_33864_28111# a_12899_10927# 0.41fF
C1487 a_10680_52245# a_28881_52271# 0.41fF
C1488 a_41462_62194# a_42466_62194# 0.97fF
C1489 a_12355_15055# a_10515_22671# 0.35fF
C1490 a_16746_57176# VDD 33.20fF
C1491 vcm_commonmode a_37446_14512# 0.87fF
C1492 a_4571_26677# a_4528_26159# 1.21fF
C1493 vcm_commonmode a_16362_20536# 4.47fF
C1494 a_28446_31375# a_28841_29575# 0.32fF
C1495 a_7571_29199# a_8273_42479# 0.37fF
C1496 a_43470_10496# VDD 0.51fF
C1497 a_16707_40183# VDD 0.61fF
C1498 vcm_commonmode a_23298_57174# 0.31fF
C1499 a_13643_28327# VDD 14.37fF
C1500 a_40366_20902# a_40458_20536# 0.32fF
C1501 a_12727_58255# a_11251_59879# 0.42fF
C1502 a_30764_7638# a_12985_7663# 0.41fF
C1503 a_16362_24552# m3_16264_24414# 2.81fF
C1504 a_29322_63198# a_29414_63198# 0.32fF
C1505 a_10873_27497# a_8935_27791# 0.39fF
C1506 a_1761_43567# a_3305_38671# 0.53fF
C1507 a_20378_57174# a_20378_56170# 1.00fF
C1508 a_46482_57174# a_47486_57174# 0.97fF
C1509 a_5024_67885# a_7773_63927# 1.06fF
C1510 vcm_commonmode a_42466_23548# 0.87fF
C1511 vcm_commonmode a_39454_66210# 0.87fF
C1512 a_3339_43023# a_2339_38129# 1.14fF
C1513 a_23141_52521# VDD 0.38fF
C1514 a_16362_21540# a_16746_21538# 2.28fF
C1515 a_27752_7638# a_12877_14441# 0.41fF
C1516 a_30418_62194# VDD 0.51fF
C1517 a_8583_33551# a_27535_30503# 1.33fF
C1518 vcm_commonmode a_16362_12504# 4.47fF
C1519 ctopn a_17366_9492# 3.42fF
C1520 a_42718_27497# a_10515_23975# 0.41fF
C1521 a_2263_68218# VDD 0.62fF
C1522 a_26631_35877# VDD 1.05fF
C1523 ctopn a_33430_16520# 3.59fF
C1524 a_5449_25071# a_5085_23047# 0.31fF
C1525 vcm_commonmode a_37354_62194# 0.31fF
C1526 a_7862_34025# a_3339_30503# 0.75fF
C1527 a_38450_15516# VDD 0.51fF
C1528 a_34062_47607# VDD 0.35fF
C1529 a_47486_71230# a_48490_71230# 0.97fF
C1530 a_23298_59182# a_23390_59182# 0.32fF
C1531 a_42709_29199# a_12899_10927# 0.40fF
C1532 a_43269_29967# a_12877_16911# 0.41fF
C1533 a_23195_29967# VDD 0.97fF
C1534 vcm_commonmode a_45386_15882# 0.31fF
C1535 a_38450_63198# ctopp 3.64fF
C1536 a_36442_71230# VDD 0.58fF
C1537 a_39247_39095# VDD 0.63fF
C1538 a_48490_11500# VDD 0.55fF
C1539 a_12341_41281# VDD 1.61fF
C1540 a_21290_17890# a_21382_17524# 0.32fF
C1541 a_12381_35836# a_12663_35431# 2.56fF
C1542 a_23535_50247# a_23631_50069# 0.37fF
C1543 vcm_commonmode a_43378_71230# 0.31fF
C1544 a_3667_60405# VDD 0.35fF
C1545 a_18979_30287# a_29175_28335# 0.35fF
C1546 a_32426_59182# ctopp 3.59fF
C1547 a_12869_2741# a_12899_2767# 4.65fF
C1548 a_27406_64202# a_27406_63198# 1.23fF
C1549 a_40366_12870# a_40458_12504# 0.32fF
C1550 vcm_commonmode a_16746_17522# 5.36fF
C1551 a_41427_52263# ctopp 2.62fF
C1552 a_2235_30503# a_23736_7638# 0.36fF
C1553 a_25787_28327# a_33430_68218# 0.38fF
C1554 a_35438_59182# a_35438_58178# 1.00fF
C1555 a_14985_51701# a_14983_51157# 1.62fF
C1556 a_37534_51701# a_37459_51183# 0.74fF
C1557 a_19374_22544# a_19374_21540# 1.00fF
C1558 a_9503_26151# a_12899_10927# 0.41fF
C1559 a_13643_28327# a_18053_28879# 1.43fF
C1560 vcm_commonmode a_22294_13874# 0.31fF
C1561 a_9503_68841# VDD 0.64fF
C1562 a_26402_13508# a_27406_13508# 0.97fF
C1563 a_5449_25071# a_6162_28487# 0.32fF
C1564 a_8782_65015# a_5254_67503# 1.16fF
C1565 vcm_commonmode a_43470_63198# 0.92fF
C1566 a_31422_68218# a_32426_68218# 0.97fF
C1567 a_3247_20495# a_2143_15271# 0.76fF
C1568 a_2971_48463# VDD 0.38fF
C1569 a_9314_69367# a_9319_69141# 0.54fF
C1570 a_42985_46831# a_48490_71230# 0.38fF
C1571 a_14287_51175# a_18370_70226# 0.38fF
C1572 a_2847_21781# VDD 0.48fF
C1573 m3_49396_69134# VDD 0.34fF
C1574 a_12869_2741# a_10964_25615# 0.37fF
C1575 a_6559_22671# a_5993_32687# 0.51fF
C1576 a_43470_56170# a_43470_55166# 1.00fF
C1577 a_48398_63198# a_48490_63198# 0.32fF
C1578 a_13909_41923# a_19967_41781# 0.57fF
C1579 a_39454_57174# a_39454_56170# 1.00fF
C1580 a_1923_59583# a_7039_65469# 0.51fF
C1581 vcm_commonmode a_37446_59182# 0.87fF
C1582 a_31768_55394# a_31422_60186# 0.38fF
C1583 a_7295_44647# a_12447_29199# 5.16fF
C1584 a_28717_42917# VDD 1.57fF
C1585 a_43362_28879# a_47486_67214# 0.38fF
C1586 a_16955_52047# a_20378_66210# 0.38fF
C1587 a_12907_56399# a_12983_63151# 0.39fF
C1588 a_35346_21906# a_35438_21540# 0.32fF
C1589 a_7571_29199# a_10873_27497# 0.85fF
C1590 a_6831_63303# a_4482_57863# 2.83fF
C1591 a_36442_60186# ctopp 3.59fF
C1592 a_39454_68218# VDD 0.51fF
C1593 a_20655_34743# VDD 0.59fF
C1594 vcm_commonmode a_17366_18528# 1.82fF
C1595 a_12357_37999# a_32327_40191# 2.65fF
C1596 a_39362_7850# VDD 0.62fF
C1597 a_19720_55394# a_19374_62194# 0.38fF
C1598 a_23390_16520# a_23390_15516# 1.00fF
C1599 a_25787_28327# a_33430_56170# 0.36fF
C1600 ctopn a_35438_22544# 3.58fF
C1601 a_21187_29415# a_18979_30287# 1.53fF
C1602 a_8583_33551# inn_analog 1.53fF
C1603 vcm_commonmode a_46390_68218# 0.31fF
C1604 a_42374_59182# a_42466_59182# 0.32fF
C1605 a_19576_51701# a_4215_51157# 0.33fF
C1606 a_32951_27247# a_33430_19532# 0.38fF
C1607 a_1823_76181# a_4119_70741# 0.53fF
C1608 a_18127_35797# a_13097_37455# 0.73fF
C1609 vcm_commonmode a_49494_21540# 0.90fF
C1610 a_21233_40956# VDD 0.85fF
C1611 a_40366_17890# a_40458_17524# 0.32fF
C1612 vcm_commonmode a_27752_7638# 10.35fF
C1613 a_5915_30287# a_20905_32143# 0.30fF
C1614 a_1586_40455# a_1591_49557# 0.32fF
C1615 a_4191_33449# a_11067_46823# 0.57fF
C1616 a_9135_49557# VDD 0.44fF
C1617 a_48398_72234# a_48490_72234# 0.32fF
C1618 a_21371_52263# a_11803_55311# 0.50fF
C1619 a_8491_27023# a_12877_14441# 0.41fF
C1620 a_26748_7638# a_26402_14512# 0.38fF
C1621 a_27314_60186# a_27406_60186# 0.32fF
C1622 vcm_commonmode a_26402_10496# 0.87fF
C1623 a_46482_64202# a_46482_63198# 1.23fF
C1624 a_16087_31751# VDD 0.44fF
C1625 ctopn a_31422_14512# 3.59fF
C1626 a_12263_4391# a_9135_27239# 1.38fF
C1627 a_12641_43124# a_14293_41807# 0.39fF
C1628 a_40050_48463# a_12981_59343# 0.40fF
C1629 a_1950_59887# a_9411_60437# 0.38fF
C1630 vcm_commonmode a_41462_60186# 0.87fF
C1631 a_6559_22671# a_5831_39189# 0.63fF
C1632 a_15959_44031# VDD 0.95fF
C1633 a_18151_52263# a_12983_63151# 0.40fF
C1634 a_22294_18894# a_22386_18528# 0.32fF
C1635 a_16219_51183# a_16385_51183# 0.40fF
C1636 a_2959_47113# a_26397_51183# 0.79fF
C1637 a_6559_59879# a_13445_50639# 1.80fF
C1638 a_38450_22544# a_38450_21540# 1.00fF
C1639 a_1952_60431# VDD 3.96fF
C1640 a_11619_3303# VDD 10.06fF
C1641 a_39454_56170# VDD 0.52fF
C1642 a_27752_7638# a_27406_22544# 0.38fF
C1643 a_45478_13508# a_46482_13508# 0.97fF
C1644 a_22386_8488# VDD 0.58fF
C1645 a_17366_68218# a_17366_67214# 1.00fF
C1646 a_21371_52263# a_12981_62313# 0.40fF
C1647 vcm_commonmode a_46390_56170# 0.31fF
C1648 ctopn a_36442_23548# 3.40fF
C1649 a_21003_49007# a_21169_49007# 0.39fF
C1650 vcm_commonmode a_29322_8854# 0.31fF
C1651 m3_49396_16382# VDD 0.35fF
C1652 vcm_commonmode a_21382_15516# 0.87fF
C1653 a_31422_56170# a_32426_56170# 0.97fF
C1654 a_32426_57174# ctopp 3.58fF
C1655 a_12809_71285# VDD 0.36fF
C1656 a_11803_55311# a_12727_58255# 1.07fF
C1657 a_42165_36367# VDD 1.62fF
C1658 ctopn a_45478_19532# 3.59fF
C1659 a_28446_31375# a_26523_29199# 0.44fF
C1660 a_5490_41365# VDD 1.24fF
C1661 a_2595_47653# VDD 2.50fF
C1662 a_21371_50959# a_25398_72234# 0.34fF
C1663 vcm_commonmode a_19374_71230# 0.86fF
C1664 a_32772_7638# a_32426_15516# 0.38fF
C1665 a_38450_61190# VDD 0.51fF
C1666 vcm_commonmode a_31422_11500# 0.87fF
C1667 a_35438_58178# a_35438_57174# 1.00fF
C1668 a_5252_56891# a_5291_56765# 0.46fF
C1669 a_8782_65015# a_8999_61493# 0.35fF
C1670 vcm_commonmode a_45386_61190# 0.31fF
C1671 a_42466_16520# a_42466_15516# 1.00fF
C1672 vcm_commonmode a_35438_24552# 0.84fF
C1673 a_49494_9492# m3_49396_9354# 2.78fF
C1674 a_28756_55394# a_12727_67753# 0.40fF
C1675 vcm_commonmode a_17274_67214# 0.33fF
C1676 a_27406_19532# a_27406_18528# 1.00fF
C1677 a_11145_60431# VDD 0.72fF
C1678 a_21187_29415# a_25269_27791# 0.49fF
C1679 a_12907_27023# a_23685_29111# 0.50fF
C1680 a_31330_10862# a_31422_10496# 0.32fF
C1681 a_46482_62194# ctopp 3.59fF
C1682 a_42466_70226# VDD 0.51fF
C1683 a_17366_68218# ctopp 3.43fF
C1684 vcm_commonmode a_45478_55166# 0.84fF
C1685 a_4941_35727# VDD 0.69fF
C1686 a_13183_52047# a_6835_46823# 0.51fF
C1687 vcm_commonmode a_37446_57174# 0.87fF
C1688 a_1586_40455# a_4240_48981# 0.52fF
C1689 a_23390_16520# VDD 0.51fF
C1690 vcm_commonmode a_49402_70226# 0.30fF
C1691 a_1689_10396# a_3143_22364# 0.32fF
C1692 a_46390_60186# a_46482_60186# 0.32fF
C1693 a_4339_64521# a_2959_47113# 0.44fF
C1694 a_11067_66191# a_10515_22671# 6.91fF
C1695 a_17274_11866# a_17366_11500# 0.32fF
C1696 vcm_commonmode a_30326_16886# 0.31fF
C1697 a_36717_47375# a_22843_29415# 0.55fF
C1698 a_17599_52263# VDD 16.21fF
C1699 a_22386_15516# a_22386_14512# 1.00fF
C1700 ctopn a_48490_20536# 3.43fF
C1701 a_46482_7484# m3_46384_7346# 2.80fF
C1702 a_26523_28111# a_18979_30287# 0.49fF
C1703 a_35493_43421# VDD 0.82fF
C1704 a_41370_18894# a_41462_18528# 0.32fF
C1705 a_3987_19623# a_8015_21807# 0.49fF
C1706 vcm_commonmode a_23395_52047# 10.02fF
C1707 a_30418_61190# a_31422_61190# 0.97fF
C1708 a_43470_55166# m3_43372_55078# 2.81fF
C1709 a_21290_24918# a_21382_24552# 0.32fF
C1710 a_15959_35327# VDD 1.04fF
C1711 a_12725_44527# a_27271_37455# 0.31fF
C1712 a_36442_68218# a_36442_67214# 1.00fF
C1713 a_38557_32143# a_38450_63198# 0.42fF
C1714 vcm_commonmode a_8491_27023# 10.30fF
C1715 vcm_commonmode a_8583_33551# 9.60fF
C1716 a_25971_52263# a_12901_66959# 0.40fF
C1717 vcm_commonmode a_22386_68218# 0.87fF
C1718 a_18151_52263# a_24394_69222# 0.38fF
C1719 a_31422_58178# VDD 0.51fF
C1720 a_3987_19623# a_5211_24759# 0.83fF
C1721 a_18278_62194# a_18370_62194# 0.32fF
C1722 a_40323_29967# VDD 0.51fF
C1723 ctopn a_48490_12504# 3.43fF
C1724 a_39222_48169# a_12907_27023# 0.53fF
C1725 a_17366_56170# ctopp 0.37fF
C1726 a_7580_61751# a_6467_55527# 0.50fF
C1727 a_11067_67279# a_19720_7638# 0.41fF
C1728 a_42466_72234# m3_42368_72146# 2.80fF
C1729 a_20655_41271# VDD 0.59fF
C1730 a_21382_69222# a_21382_68218# 1.00fF
C1731 a_14831_50095# a_26662_48981# 0.33fF
C1732 a_17600_50345# VDD 0.73fF
C1733 a_38557_32143# a_41427_52263# 1.91fF
C1734 a_25787_28327# a_43267_31055# 3.84fF
C1735 a_16362_20536# a_16746_20534# 2.28fF
C1736 a_5749_60039# VDD 0.40fF
C1737 a_1689_10396# a_2317_28892# 1.19fF
C1738 a_33430_8488# a_34434_8488# 0.97fF
C1739 a_48490_67214# VDD 0.54fF
C1740 a_1586_36727# a_1757_38677# 0.51fF
C1741 a_23298_57174# a_23390_57174# 0.32fF
C1742 a_2292_17179# a_1591_12565# 0.34fF
C1743 a_26310_15882# a_26402_15516# 0.32fF
C1744 ctopn a_43470_21540# 3.59fF
C1745 a_4811_34855# a_21012_30761# 0.57fF
C1746 a_28152_44869# VDD 1.52fF
C1747 a_2952_66139# a_4307_67477# 0.84fF
C1748 a_34434_70226# a_35438_70226# 0.97fF
C1749 a_46482_19532# a_46482_18528# 1.00fF
C1750 a_2899_28111# VDD 0.38fF
C1751 vcm_commonmode a_36442_13508# 0.87fF
C1752 a_45478_59182# a_45478_58178# 1.00fF
C1753 a_12981_59343# ctopp 3.23fF
C1754 ctopn a_20378_10496# 3.59fF
C1755 a_18370_69222# VDD 0.52fF
C1756 ctopn a_48490_17524# 3.43fF
C1757 a_18611_52047# a_23390_55166# 0.46fF
C1758 a_45478_9492# VDD 0.51fF
C1759 a_4443_46607# a_6372_38279# 1.00fF
C1760 vcm_commonmode a_22386_56170# 0.87fF
C1761 a_5915_30287# a_8753_31055# 0.46fF
C1762 a_24302_71230# a_24394_71230# 0.32fF
C1763 vcm_commonmode a_25306_69222# 0.31fF
C1764 a_32426_60186# a_32426_59182# 1.00fF
C1765 a_20713_39105# a_21479_39141# 0.31fF
C1766 a_25398_22544# VDD 0.51fF
C1767 a_26748_7638# a_12895_13967# 0.41fF
C1768 a_28756_7638# a_12985_19087# 0.41fF
C1769 a_16746_65208# VDD 33.19fF
C1770 a_21382_63198# a_21382_62194# 1.00fF
C1771 a_36350_11866# a_36442_11500# 0.32fF
C1772 a_30790_30663# VDD 0.83fF
C1773 a_41462_15516# a_41462_14512# 1.00fF
C1774 vcm_commonmode a_32334_22910# 0.31fF
C1775 a_20378_70226# ctopp 3.58fF
C1776 a_2473_34293# a_3301_27791# 0.62fF
C1777 a_37446_58178# ctopp 3.59fF
C1778 vcm_commonmode a_23298_65206# 0.31fF
C1779 a_34780_56398# a_12355_65103# 0.40fF
C1780 a_12473_36341# a_12641_36596# 0.39fF
C1781 a_18335_50645# a_18501_50645# 0.51fF
C1782 a_23487_50095# VDD 0.53fF
C1783 a_1586_69367# a_1757_71317# 0.61fF
C1784 a_12907_27023# a_19720_7638# 0.85fF
C1785 a_20635_29415# a_36797_27497# 0.49fF
C1786 a_26402_9492# a_26402_8488# 1.00fF
C1787 a_11069_23983# VDD 0.45fF
C1788 a_40366_24918# a_40458_24552# 0.32fF
C1789 a_11067_23759# a_12899_11471# 0.35fF
C1790 a_16362_12504# a_16746_12502# 2.28fF
C1791 a_12355_15055# a_6162_28487# 0.33fF
C1792 a_18611_52047# a_19576_51701# 0.96fF
C1793 vcm_commonmode a_21382_61190# 0.87fF
C1794 a_21382_67214# a_22386_67214# 0.97fF
C1795 a_21382_14512# VDD 0.51fF
C1796 a_47486_64202# VDD 0.51fF
C1797 a_18979_30287# a_30440_31573# 0.43fF
C1798 a_37354_62194# a_37446_62194# 0.32fF
C1799 vcm_commonmode a_28318_14878# 0.31fF
C1800 ctopn a_25398_11500# 3.59fF
C1801 a_31096_38341# VDD 1.56fF
C1802 a_11067_67279# a_40491_27247# 0.41fF
C1803 VDD dummypin[2] 0.90fF
C1804 a_40458_69222# a_40458_68218# 1.00fF
C1805 a_42718_27497# a_44474_8488# 0.38fF
C1806 a_7841_12167# a_6459_30511# 0.44fF
C1807 a_3301_16617# VDD 0.49fF
C1808 vcm_commonmode a_25398_70226# 0.87fF
C1809 a_1923_54591# a_9707_51325# 0.35fF
C1810 a_49402_60186# VDD 0.31fF
C1811 a_42466_58178# vcm_commonmode 0.87fF
C1812 a_8273_42479# a_6649_25615# 0.53fF
C1813 a_30418_8488# a_30418_7484# 1.00fF
C1814 a_26402_23548# VDD 0.52fF
C1815 a_23390_66210# VDD 0.51fF
C1816 a_19807_28111# a_31659_31751# 0.81fF
C1817 a_19626_31751# VDD 2.34fF
C1818 a_40585_42369# a_41351_42405# 0.37fF
C1819 a_42374_57174# a_42466_57174# 0.32fF
C1820 a_45386_15882# a_45478_15516# 0.32fF
C1821 vcm_commonmode a_33338_23914# 0.31fF
C1822 a_1593_42479# VDD 0.40fF
C1823 vcm_commonmode a_30326_66210# 0.31fF
C1824 a_43175_28335# a_46482_10496# 0.38fF
C1825 VDD conversion_finished_out 0.68fF
C1826 a_23390_58178# a_24394_58178# 0.97fF
C1827 a_13123_38231# a_12381_35836# 0.35fF
C1828 a_35438_19532# VDD 0.51fF
C1829 a_8491_41383# a_37527_29397# 0.36fF
C1830 a_18370_9492# a_19374_9492# 0.97fF
C1831 a_11430_26159# VDD 1.10fF
C1832 a_26402_55166# m3_26304_55078# 2.81fF
C1833 a_19374_13508# a_19374_12504# 1.00fF
C1834 vcm_commonmode a_42374_19898# 0.31fF
C1835 a_26402_67214# ctopp 3.59fF
C1836 a_34434_16520# a_35438_16520# 0.97fF
C1837 a_43378_71230# a_43470_71230# 0.32fF
C1838 vcm_commonmode a_43470_8488# 0.86fF
C1839 m3_42368_7346# VDD 0.33fF
C1840 a_40458_63198# a_40458_62194# 1.00fF
C1841 a_6831_63303# a_2775_46025# 1.61fF
C1842 a_11866_27791# a_11430_26159# 0.51fF
C1843 a_13835_41001# a_12801_38517# 0.39fF
C1844 a_22411_39095# VDD 0.60fF
C1845 a_16746_17522# a_12899_11471# 2.28fF
C1846 a_45478_9492# a_45478_8488# 1.00fF
C1847 a_43378_24918# VDD 0.36fF
C1848 a_11711_32143# VDD 0.51fF
C1849 a_45478_58178# a_45478_57174# 1.00fF
C1850 a_11521_66567# a_10975_66407# 0.44fF
C1851 a_40458_67214# a_41462_67214# 0.97fF
C1852 a_34780_56398# ctopp 2.62fF
C1853 vcm_commonmode a_31422_67214# 0.87fF
C1854 a_29760_55394# a_29414_68218# 0.38fF
C1855 a_11067_47695# a_11067_46823# 1.49fF
C1856 a_4215_51157# a_17039_51157# 1.80fF
C1857 a_38450_20536# VDD 0.51fF
C1858 a_2559_52789# config_2_in[15] 0.33fF
C1859 a_27406_63198# VDD 0.57fF
C1860 a_1761_50639# a_35196_35425# 0.39fF
C1861 a_22294_13874# a_22386_13508# 0.32fF
C1862 vcm_commonmode a_45386_20902# 0.31fF
C1863 a_12641_37684# VDD 6.30fF
C1864 a_27314_68218# a_27406_68218# 0.32fF
C1865 vcm_commonmode a_34342_63198# 0.31fF
C1866 a_5915_35943# a_8753_31055# 0.37fF
C1867 a_39299_48783# a_44474_71230# 0.38fF
C1868 a_21382_59182# VDD 0.51fF
C1869 a_49494_18528# m3_49396_18390# 2.78fF
C1870 a_49494_8488# a_49494_7484# 1.00fF
C1871 a_26402_7484# a_27406_7484# 0.97fF
C1872 vcm_commonmode a_28410_9492# 0.87fF
C1873 a_3339_32463# a_2235_30503# 1.43fF
C1874 a_7773_63927# a_7210_55081# 0.87fF
C1875 vcm_commonmode a_44474_16520# 0.87fF
C1876 a_25398_64202# ctopp 3.59fF
C1877 ctopn a_30418_13508# 3.59fF
C1878 a_23395_52047# a_27406_60186# 0.38fF
C1879 vcm_commonmode a_28318_59182# 0.31fF
C1880 a_2235_30503# a_7841_29673# 0.39fF
C1881 a_4811_34855# a_32167_29611# 0.41fF
C1882 a_33694_30761# a_32823_29397# 0.33fF
C1883 a_7862_34025# a_20505_29967# 0.54fF
C1884 a_4443_46607# a_1761_44111# 0.38fF
C1885 a_38450_12504# VDD 0.51fF
C1886 a_41872_29423# a_43470_67214# 0.38fF
C1887 a_1761_37039# a_1761_35407# 1.27fF
C1888 a_12473_37429# a_13005_35823# 0.76fF
C1889 a_37446_9492# a_38450_9492# 0.97fF
C1890 vcm_commonmode a_45386_12870# 0.31fF
C1891 a_20378_64202# a_21382_64202# 0.97fF
C1892 a_38450_13508# a_38450_12504# 1.00fF
C1893 a_14076_35077# VDD 1.36fF
C1894 a_29760_55394# a_29414_56170# 0.38fF
C1895 a_5959_13621# VDD 0.53fF
C1896 a_25019_47679# VDD 0.35fF
C1897 a_1950_59887# a_7580_61751# 0.39fF
C1898 a_33430_21540# VDD 0.51fF
C1899 vcm_commonmode a_36442_7484# 0.68fF
C1900 a_27752_7638# a_12899_11471# 0.41fF
C1901 a_17366_22544# a_18370_22544# 0.97fF
C1902 a_31768_7638# a_31422_24552# 0.47fF
C1903 a_7803_55509# a_7676_61493# 0.31fF
C1904 vcm_commonmode a_40366_21906# 0.31fF
C1905 a_34434_69222# ctopp 3.59fF
C1906 a_11140_10107# VDD 0.63fF
C1907 vcm_commonmode a_30418_64202# 0.87fF
C1908 a_1761_35407# a_1761_32143# 0.51fF
C1909 a_38450_17524# VDD 0.51fF
C1910 vcm_commonmode a_12516_7093# 6.33fF
C1911 a_25398_60186# VDD 0.51fF
C1912 vcm_commonmode a_17274_10862# 0.33fF
C1913 a_43269_29967# a_12895_13967# 0.41fF
C1914 vcm_commonmode a_45386_17890# 0.31fF
C1915 a_32426_65206# ctopp 3.59fF
C1916 a_8003_72917# VDD 1.91fF
C1917 a_28410_67214# a_28410_66210# 1.00fF
C1918 vcm_commonmode a_32334_60186# 0.31fF
C1919 a_38557_32143# a_12981_59343# 0.40fF
C1920 a_28756_7638# a_28410_10496# 0.38fF
C1921 a_2775_46025# a_12993_50345# 0.51fF
C1922 a_13669_39605# a_13097_37455# 2.74fF
C1923 a_24394_65206# a_24394_64202# 1.00fF
C1924 a_41370_13874# a_41462_13508# 0.32fF
C1925 a_18197_36604# VDD 0.92fF
C1926 vcm_commonmode a_18370_19532# 0.88fF
C1927 a_1803_20719# a_13716_43047# 1.46fF
C1928 a_46390_68218# a_46482_68218# 0.32fF
C1929 a_19720_55394# a_12981_62313# 0.40fF
C1930 a_5399_13255# VDD 1.17fF
C1931 vcm_commonmode a_39454_69222# 0.87fF
C1932 a_6775_53877# a_10503_52828# 0.37fF
C1933 a_45478_7484# a_46482_7484# 0.97fF
C1934 a_4758_45369# a_6775_53877# 1.40fF
C1935 a_18370_23548# a_18370_22544# 1.00fF
C1936 a_28547_51175# a_16863_29415# 5.91fF
C1937 a_12473_42869# a_13909_39747# 0.46fF
C1938 a_27314_56170# a_27406_56170# 0.32fF
C1939 a_1591_71317# VDD 0.37fF
C1940 a_52778_39936# VDD 1.16fF
C1941 vcm_commonmode a_46482_22544# 0.87fF
C1942 a_10531_31055# a_13353_30511# 0.63fF
C1943 vcm_commonmode a_37446_65206# 0.87fF
C1944 a_29414_69222# a_30418_69222# 0.97fF
C1945 a_39454_18528# VDD 0.51fF
C1946 a_24394_61190# a_24394_60186# 1.00fF
C1947 a_19374_24552# VDD 0.60fF
C1948 vcm_commonmode a_22294_11866# 0.31fF
C1949 ctopn a_37446_8488# 3.40fF
C1950 a_4443_46607# a_12621_36091# 10.65fF
C1951 a_39454_64202# a_40458_64202# 0.97fF
C1952 a_11521_66567# a_10055_58791# 0.35fF
C1953 vcm_commonmode a_46390_18894# 0.31fF
C1954 a_39454_66210# ctopp 3.59fF
C1955 vcm_commonmode a_26310_24918# 0.31fF
C1956 a_17507_52047# a_12727_67753# 0.40fF
C1957 a_30418_55166# VDD 0.60fF
C1958 a_10515_63143# a_4191_33449# 0.55fF
C1959 a_36442_22544# a_37446_22544# 0.97fF
C1960 a_12447_29199# a_9405_31599# 0.48fF
C1961 a_2021_22325# a_5993_32687# 0.47fF
C1962 a_21382_57174# VDD 0.51fF
C1963 vcm_commonmode a_42466_14512# 0.87fF
C1964 a_27406_65206# a_28410_65206# 0.97fF
C1965 a_5915_30287# VDD 9.83fF
C1966 vcm_commonmode a_21382_20536# 0.87fF
C1967 vcm_commonmode a_36350_55166# 0.30fF
C1968 a_48490_10496# VDD 0.54fF
C1969 a_23390_17524# a_23390_16520# 1.00fF
C1970 vcm_commonmode a_28318_57174# 0.31fF
C1971 a_7000_43541# VDD 5.84fF
C1972 a_1950_59887# a_8531_70543# 0.31fF
C1973 a_4891_47388# a_5135_50069# 0.45fF
C1974 a_2124_59459# VDD 0.44fF
C1975 a_32772_7638# a_32426_20536# 0.38fF
C1976 a_18370_23548# a_19374_23548# 0.97fF
C1977 VDD config_1_in[14] 1.06fF
C1978 a_27406_56170# a_27406_55166# 1.00fF
C1979 a_5449_25071# VDD 1.44fF
C1980 a_1761_41935# a_13909_41923# 0.81fF
C1981 a_47486_67214# a_47486_66210# 1.00fF
C1982 vcm_commonmode a_47486_23548# 0.87fF
C1983 a_39454_7484# m3_39356_7346# 2.80fF
C1984 a_21712_43781# VDD 1.71fF
C1985 vcm_commonmode a_44474_66210# 0.87fF
C1986 a_28881_52271# VDD 4.40fF
C1987 vcm_commonmode a_16955_52047# 10.02fF
C1988 a_8491_27023# a_12899_11471# 0.41fF
C1989 a_35438_62194# VDD 0.51fF
C1990 a_26310_61190# a_26402_61190# 0.32fF
C1991 a_36442_55166# m3_36344_55078# 2.81fF
C1992 vcm_commonmode a_21382_12504# 0.87fF
C1993 ctopn a_22386_9492# 3.58fF
C1994 a_1799_29556# a_1761_27791# 2.10fF
C1995 a_43470_65206# a_43470_64202# 1.00fF
C1996 ctopn a_38450_16520# 3.59fF
C1997 a_40050_48463# a_45478_55166# 0.63fF
C1998 a_34780_56398# a_34434_63198# 0.42fF
C1999 vcm_commonmode a_42374_62194# 0.31fF
C2000 a_13643_28327# a_24959_30503# 0.47fF
C2001 a_43470_15516# VDD 0.51fF
C2002 a_16955_52047# a_20378_69222# 0.38fF
C2003 a_18611_52047# a_12901_66959# 0.40fF
C2004 a_27406_19532# a_28410_19532# 0.97fF
C2005 a_32772_7638# a_32426_12504# 0.38fF
C2006 a_5239_20693# VDD 0.53fF
C2007 a_37446_23548# a_37446_22544# 1.00fF
C2008 a_20635_29415# a_21012_30761# 0.56fF
C2009 a_43470_63198# ctopp 3.64fF
C2010 a_25787_28327# a_12907_27023# 0.58fF
C2011 a_10873_27497# a_12341_3311# 0.70fF
C2012 a_1761_41935# a_1761_39215# 0.87fF
C2013 a_23789_39100# a_24561_41583# 0.39fF
C2014 a_46390_56170# a_46482_56170# 0.32fF
C2015 a_41462_71230# VDD 0.58fF
C2016 a_31422_66210# a_31422_65206# 1.00fF
C2017 a_32426_14512# a_33430_14512# 0.97fF
C2018 vcm_commonmode a_16746_21538# 5.36fF
C2019 a_5831_39189# a_2021_22325# 0.47fF
C2020 a_5885_39759# VDD 0.69fF
C2021 a_48490_69222# a_49494_69222# 0.97fF
C2022 a_34251_52263# a_32823_29397# 1.26fF
C2023 a_13097_36367# a_13669_35253# 5.52fF
C2024 a_12877_16911# VDD 7.21fF
C2025 a_35438_72234# a_36442_72234# 0.97fF
C2026 a_23395_52047# a_40050_48463# 0.58fF
C2027 a_25971_52263# a_41261_28335# 9.18fF
C2028 vcm_commonmode a_48398_71230# 0.31fF
C2029 a_43470_61190# a_43470_60186# 1.00fF
C2030 a_29322_8854# a_29414_8488# 0.32fF
C2031 a_7841_22895# VDD 1.37fF
C2032 a_37446_59182# ctopp 3.59fF
C2033 a_2840_53511# a_2952_53333# 0.39fF
C2034 a_29760_7638# a_29414_22544# 0.38fF
C2035 vcm_commonmode a_21382_17524# 0.87fF
C2036 a_38557_32143# a_37534_51701# 0.31fF
C2037 a_12357_37999# a_19967_41781# 0.42fF
C2038 a_5779_75093# VDD 0.35fF
C2039 a_12983_63151# a_16362_66210# 1.15fF
C2040 a_20378_13508# VDD 0.51fF
C2041 a_30326_70226# a_30418_70226# 0.32fF
C2042 a_2451_72373# a_9314_69367# 0.35fF
C2043 a_32772_7638# a_32426_17524# 0.38fF
C2044 a_18979_30287# a_33641_29967# 0.35fF
C2045 a_29414_62194# a_29414_61190# 1.00fF
C2046 a_20378_10496# a_20378_9492# 1.00fF
C2047 a_28756_7638# VDD 6.32fF
C2048 a_2099_59861# a_3143_22364# 0.39fF
C2049 vcm_commonmode a_27314_13874# 0.31fF
C2050 a_46482_65206# a_47486_65206# 0.97fF
C2051 a_19780_37253# VDD 1.73fF
C2052 a_19720_55394# a_19374_55166# 0.46fF
C2053 vcm_commonmode a_48490_63198# 0.92fF
C2054 a_42466_17524# a_42466_16520# 1.00fF
C2055 a_21187_29415# a_18703_29199# 0.84fF
C2056 a_7553_48469# VDD 0.31fF
C2057 a_29414_20536# a_29414_19532# 1.00fF
C2058 a_16362_22544# VDD 2.47fF
C2059 a_37446_23548# a_38450_23548# 0.97fF
C2060 a_12869_2741# a_9135_27239# 3.05fF
C2061 a_43470_72234# VDD 1.23fF
C2062 a_43267_31055# a_12727_58255# 0.40fF
C2063 a_34434_66210# a_35438_66210# 0.97fF
C2064 vcm_commonmode a_42466_59182# 0.87fF
C2065 a_5039_42167# a_1803_19087# 1.38fF
C2066 a_39431_43177# VDD 0.62fF
C2067 a_23395_52047# a_12355_65103# 0.40fF
C2068 a_12869_2741# a_7571_29199# 0.84fF
C2069 vcm_commonmode a_48490_72234# 0.68fF
C2070 a_33864_28111# a_34434_16520# 0.38fF
C2071 a_8500_58799# VDD 0.51fF
C2072 a_8583_33551# a_11067_46823# 0.46fF
C2073 a_45386_61190# a_45478_61190# 0.32fF
C2074 a_41462_60186# ctopp 3.59fF
C2075 a_44474_68218# VDD 0.51fF
C2076 a_4443_46607# a_12473_36341# 0.92fF
C2077 a_19807_28111# a_4811_34855# 0.70fF
C2078 a_30875_34743# VDD 0.64fF
C2079 vcm_commonmode a_22386_18528# 0.87fF
C2080 a_44382_7850# VDD 0.62fF
C2081 a_17274_67214# a_17366_67214# 0.32fF
C2082 ctopn a_40458_22544# 3.58fF
C2083 a_34434_71230# a_34434_70226# 1.00fF
C2084 a_46482_19532# a_47486_19532# 0.97fF
C2085 a_27167_52271# a_2872_44111# 0.73fF
C2086 a_41335_29423# VDD 0.33fF
C2087 a_4351_67279# VDD 13.14fF
C2088 a_5915_35943# VDD 6.62fF
C2089 a_12663_39783# VDD 3.20fF
C2090 a_36797_27497# a_37446_8488# 0.38fF
C2091 a_12381_35836# a_31131_35281# 0.42fF
C2092 a_2686_70223# a_5682_69367# 0.41fF
C2093 a_30418_20536# a_31422_20536# 0.97fF
C2094 a_48398_8854# a_48490_8488# 0.32fF
C2095 vcm_commonmode a_31422_10496# 0.87fF
C2096 vcm_commonmode a_77086_40693# 138.80fF
C2097 a_19374_63198# a_20378_63198# 0.97fF
C2098 ctopn a_36442_14512# 3.59fF
C2099 vcm_commonmode a_46482_60186# 0.87fF
C2100 a_19374_71230# ctopp 3.40fF
C2101 a_49402_70226# a_49494_70226# 0.32fF
C2102 a_19282_58178# a_19374_58178# 0.32fF
C2103 a_48490_62194# a_48490_61190# 1.00fF
C2104 a_39454_10496# a_39454_9492# 1.00fF
C2105 a_19374_55166# m3_19276_55078# 2.81fF
C2106 a_44474_56170# VDD 0.52fF
C2107 a_11067_66191# a_12985_19087# 1.08fF
C2108 a_13097_39631# a_14293_39631# 0.39fF
C2109 a_8491_41383# a_7841_12167# 1.76fF
C2110 a_11067_67279# a_11480_23957# 1.06fF
C2111 a_11067_23759# a_9955_20969# 0.83fF
C2112 a_1761_44111# a_18662_43671# 1.12fF
C2113 a_1761_25071# a_36392_43677# 0.46fF
C2114 a_27406_8488# VDD 0.58fF
C2115 vcm_commonmode a_18370_62194# 0.88fF
C2116 a_30326_16886# a_30418_16520# 0.32fF
C2117 ctopn a_41462_23548# 3.40fF
C2118 a_2419_48783# a_7251_50069# 0.78fF
C2119 a_4891_47388# a_17682_50095# 0.48fF
C2120 a_48490_20536# a_48490_19532# 1.00fF
C2121 a_3339_43023# a_1689_10396# 1.62fF
C2122 vcm_commonmode a_34342_8854# 0.31fF
C2123 m3_16264_8350# VDD 0.30fF
C2124 a_2959_47113# a_8295_47388# 1.19fF
C2125 a_1757_29973# VDD 0.64fF
C2126 vcm_commonmode a_26402_15516# 0.87fF
C2127 a_24800_41953# a_25221_41281# 0.47fF
C2128 a_1761_41935# a_3759_39991# 0.65fF
C2129 a_37446_57174# ctopp 3.58fF
C2130 a_11067_67279# a_32772_7638# 0.41fF
C2131 a_11711_50645# VDD 0.43fF
C2132 vcm_commonmode a_24394_71230# 0.86fF
C2133 a_28410_21540# a_28410_20536# 1.00fF
C2134 a_43470_61190# VDD 0.51fF
C2135 vcm_commonmode a_36442_11500# 0.87fF
C2136 a_30418_12504# a_31422_12504# 0.97fF
C2137 a_1761_46287# a_27263_40871# 0.41fF
C2138 a_36350_67214# a_36442_67214# 0.32fF
C2139 vcm_commonmode a_40458_24552# 0.84fF
C2140 a_23395_52047# ctopp 3.20fF
C2141 a_7862_34025# a_14926_31849# 1.49fF
C2142 a_7939_30503# a_8753_31055# 1.99fF
C2143 a_18703_29199# a_26523_28111# 1.73fF
C2144 vcm_commonmode a_22294_67214# 0.31fF
C2145 a_21371_50959# a_25398_68218# 0.38fF
C2146 a_4215_51157# a_9707_51325# 0.62fF
C2147 VDD inp_analog 5.27fF
C2148 a_21371_52263# a_3339_32463# 3.75fF
C2149 a_8583_33551# ctopp 2.54fF
C2150 a_47486_70226# VDD 0.51fF
C2151 a_25517_37455# VDD 4.32fF
C2152 a_22386_68218# ctopp 3.59fF
C2153 a_14258_44527# a_13984_43781# 0.45fF
C2154 a_1761_8751# VDD 1.11fF
C2155 vcm_commonmode a_42466_57174# 0.87fF
C2156 a_17682_50095# a_28524_47919# 0.58fF
C2157 a_28410_16520# VDD 0.51fF
C2158 a_39222_48169# a_40458_71230# 0.38fF
C2159 a_1586_69367# a_1775_67503# 0.33fF
C2160 a_6880_58773# VDD 0.49fF
C2161 a_22294_7850# a_22386_7484# 0.32fF
C2162 vcm_commonmode a_19282_9858# 0.31fF
C2163 a_38450_63198# a_39454_63198# 0.97fF
C2164 vcm_commonmode a_35346_16886# 0.31fF
C2165 a_18611_52047# a_23390_60186# 0.38fF
C2166 a_18539_47617# a_18500_47491# 0.42fF
C2167 a_12473_42869# VDD 8.68fF
C2168 a_39389_52271# a_39454_67214# 0.38fF
C2169 a_11943_69367# a_12039_69367# 0.36fF
C2170 a_4351_67279# a_11619_56615# 0.46fF
C2171 a_11619_56615# a_5915_35943# 0.37fF
C2172 a_25398_21540# a_26402_21540# 0.97fF
C2173 a_33338_9858# a_33430_9492# 0.32fF
C2174 a_1959_26703# VDD 0.50fF
C2175 a_12755_53030# VDD 1.31fF
C2176 a_20378_7484# VDD 1.24fF
C2177 a_49402_16886# a_49494_16520# 0.32fF
C2178 a_21371_50959# a_25398_56170# 0.38fF
C2179 ctopn a_11067_21583# 3.22fF
C2180 a_14634_47349# VDD 0.36fF
C2181 vcm_commonmode a_27406_68218# 0.87fF
C2182 a_36442_58178# VDD 0.51fF
C2183 a_6559_59663# a_3714_58345# 0.45fF
C2184 a_32426_59182# a_33430_59182# 0.97fF
C2185 a_1823_76181# a_6271_72943# 0.51fF
C2186 a_12355_15055# VDD 15.53fF
C2187 a_17599_52263# a_24959_30503# 6.35fF
C2188 a_7369_24233# a_9669_26703# 0.55fF
C2189 a_1761_41935# a_1799_29556# 0.62fF
C2190 a_22386_56170# ctopp 3.40fF
C2191 a_11067_67279# a_37919_28111# 0.41fF
C2192 ctopn a_16746_18526# 1.68fF
C2193 a_45478_72234# m3_45380_72146# 2.80fF
C2194 a_31004_40743# VDD 1.84fF
C2195 vcm_commonmode a_21290_64202# 0.31fF
C2196 a_40675_27791# a_41462_8488# 0.38fF
C2197 a_30418_17524# a_31422_17524# 0.97fF
C2198 a_17712_7638# a_17366_8488# 0.38fF
C2199 a_1761_50639# a_5039_42167# 0.82fF
C2200 a_41370_72234# a_41462_72234# 0.32fF
C2201 a_47486_21540# a_47486_20536# 1.00fF
C2202 a_16746_60188# VDD 33.19fF
C2203 a_17366_60186# a_18370_60186# 0.97fF
C2204 a_33430_55166# a_34434_55166# 0.97fF
C2205 a_34434_24552# a_34434_23548# 1.00fF
C2206 a_19374_12504# a_19374_11500# 1.00fF
C2207 a_31659_31751# VDD 1.23fF
C2208 a_1923_73087# VDD 6.81fF
C2209 a_31768_55394# a_12981_59343# 0.40fF
C2210 a_1586_18695# a_11179_9981# 0.48fF
C2211 ctopn a_48490_21540# 3.43fF
C2212 a_4351_67279# a_7571_68047# 0.54fF
C2213 a_13097_37455# a_16152_37601# 0.94fF
C2214 a_10786_19881# VDD 0.44fF
C2215 a_31768_7638# a_12727_13353# 0.41fF
C2216 a_24740_7638# a_12877_16911# 0.41fF
C2217 a_6831_63303# a_5190_59575# 0.41fF
C2218 a_7461_27247# VDD 0.81fF
C2219 vcm_commonmode a_41462_13508# 0.87fF
C2220 a_21382_61190# ctopp 3.59fF
C2221 ctopn a_25398_10496# 3.59fF
C2222 a_4351_26703# a_7203_24527# 0.55fF
C2223 a_23390_69222# VDD 0.51fF
C2224 a_12713_36483# VDD 2.26fF
C2225 vcm_commonmode a_27406_56170# 0.87fF
C2226 a_49494_11500# m3_49396_11362# 2.78fF
C2227 a_10673_15055# VDD 0.30fF
C2228 vcm_commonmode a_30326_69222# 0.31fF
C2229 a_40050_48463# a_12516_7093# 0.40fF
C2230 a_19720_7638# a_19374_13508# 0.38fF
C2231 a_6559_59663# a_7519_59575# 0.30fF
C2232 a_41370_7850# a_41462_7484# 0.32fF
C2233 a_30418_22544# VDD 0.51fF
C2234 a_21382_65206# VDD 0.51fF
C2235 a_4427_30511# VDD 1.92fF
C2236 a_11067_23759# a_12985_7663# 0.34fF
C2237 a_19967_41781# a_38011_42035# 0.83fF
C2238 a_13067_38517# a_39836_38567# 0.34fF
C2239 a_7917_13885# a_1929_12131# 0.32fF
C2240 vcm_commonmode a_37354_22910# 0.31fF
C2241 a_25398_70226# ctopp 3.58fF
C2242 a_3063_9295# VDD 0.61fF
C2243 a_42466_58178# ctopp 3.59fF
C2244 a_12283_42359# VDD 0.62fF
C2245 vcm_commonmode a_28318_65206# 0.31fF
C2246 a_25306_69222# a_25398_69222# 0.32fF
C2247 a_1586_18695# a_8123_14741# 0.53fF
C2248 a_31422_18528# a_31422_17524# 1.00fF
C2249 a_12473_36341# a_13097_36367# 0.39fF
C2250 a_14287_51175# a_18370_72234# 0.34fF
C2251 a_12985_7663# a_16362_20536# 19.89fF
C2252 a_44474_21540# a_45478_21540# 0.97fF
C2253 a_30764_7638# a_12727_13353# 0.41fF
C2254 a_35346_64202# a_35438_64202# 0.32fF
C2255 a_25263_34473# VDD 0.59fF
C2256 ctopn a_20378_15516# 3.59fF
C2257 vcm_commonmode a_26402_61190# 0.87fF
C2258 a_26402_14512# VDD 0.51fF
C2259 a_11251_59879# a_4674_40277# 1.88fF
C2260 a_13909_38659# a_12473_37429# 1.21fF
C2261 a_11067_63143# a_12899_11471# 0.41fF
C2262 a_21290_55166# VDD 0.35fF
C2263 a_32334_22910# a_32426_22544# 0.32fF
C2264 a_21382_10496# a_22386_10496# 0.97fF
C2265 vcm_commonmode a_33338_14878# 0.31fF
C2266 ctopn a_30418_11500# 3.59fF
C2267 a_31768_7638# a_10515_23975# 0.41fF
C2268 a_23298_65206# a_23390_65206# 0.32fF
C2269 a_32426_14512# a_32426_13508# 1.00fF
C2270 a_13183_52047# a_17366_64202# 0.38fF
C2271 a_12516_7093# a_12355_65103# 0.75fF
C2272 ctopn a_34434_24552# 0.65fF
C2273 a_49494_12504# m3_49396_12366# 2.78fF
C2274 vcm_commonmode a_30418_70226# 0.87fF
C2275 a_26523_28111# a_25744_7638# 0.82fF
C2276 a_8273_42479# a_8485_29673# 0.77fF
C2277 a_36442_60186# a_37446_60186# 0.97fF
C2278 a_31422_23548# VDD 0.52fF
C2279 a_28410_66210# VDD 0.51fF
C2280 a_38450_12504# a_38450_11500# 1.00fF
C2281 a_3247_20495# a_4941_35727# 1.47fF
C2282 a_16362_72234# VDD 1.77fF
C2283 a_10975_66407# a_16746_66212# 0.41fF
C2284 a_11619_56615# a_12355_15055# 1.86fF
C2285 vcm_commonmode a_38358_23914# 0.31fF
C2286 a_32426_7484# m3_32328_7346# 2.80fF
C2287 a_10935_11989# VDD 0.38fF
C2288 vcm_commonmode a_35346_66210# 0.31fF
C2289 a_25398_70226# a_25398_69222# 1.00fF
C2290 a_31422_18528# a_32426_18528# 0.97fF
C2291 a_13123_38231# a_1761_35407# 1.01fF
C2292 a_2872_44111# a_4191_33449# 0.42fF
C2293 a_40458_19532# VDD 0.51fF
C2294 a_1923_54591# a_2124_56891# 0.43fF
C2295 a_30764_7638# a_10515_23975# 0.41fF
C2296 a_2012_68565# VDD 0.30fF
C2297 a_15968_36061# VDD 2.72fF
C2298 vcm_commonmode a_47394_19898# 0.31fF
C2299 a_2315_24540# config_1_in[15] 0.46fF
C2300 a_31422_67214# ctopp 3.59fF
C2301 a_41427_52263# a_41462_55166# 0.47fF
C2302 a_25971_52263# a_30418_63198# 0.42fF
C2303 a_1768_16367# a_1915_35015# 0.61fF
C2304 a_23298_19898# a_23390_19532# 0.32fF
C2305 a_11887_19087# VDD 0.49fF
C2306 vcm_commonmode a_48490_8488# 0.85fF
C2307 a_12907_27023# a_16228_28335# 0.43fF
C2308 a_6515_62037# a_6559_59663# 0.32fF
C2309 a_6417_62215# a_6467_55527# 0.36fF
C2310 a_24394_11500# a_24394_10496# 1.00fF
C2311 a_15799_29941# VDD 0.72fF
C2312 a_13183_52047# a_26465_48463# 0.53fF
C2313 a_49494_66210# m3_49396_66122# 2.78fF
C2314 vcm_commonmode a_19374_58178# 0.87fF
C2315 a_28318_14878# a_28410_14512# 0.32fF
C2316 a_34639_42089# VDD 0.59fF
C2317 a_44382_69222# a_44474_69222# 0.32fF
C2318 a_3339_43023# a_1761_27791# 0.98fF
C2319 a_25971_52263# a_34251_52263# 1.16fF
C2320 a_28547_51175# a_25787_28327# 4.27fF
C2321 a_43175_28335# a_46482_15516# 0.38fF
C2322 a_12447_29199# a_12899_3855# 2.01fF
C2323 a_2787_32679# a_2317_28892# 0.37fF
C2324 a_22386_55166# a_23390_55166# 0.97fF
C2325 a_36797_27497# a_11067_21583# 0.41fF
C2326 a_3339_32463# a_4495_35925# 0.69fF
C2327 a_26417_47919# a_27393_47919# 0.62fF
C2328 a_15607_46805# a_7295_44647# 0.48fF
C2329 vcm_commonmode a_36442_67214# 0.87fF
C2330 a_43470_20536# VDD 0.51fF
C2331 a_32426_63198# VDD 0.57fF
C2332 a_40458_10496# a_41462_10496# 0.97fF
C2333 a_1591_69141# VDD 0.49fF
C2334 a_42374_65206# a_42466_65206# 0.32fF
C2335 a_4242_35407# VDD 0.53fF
C2336 a_14926_31849# a_23298_28487# 0.34fF
C2337 a_34699_38771# VDD 1.61fF
C2338 vcm_commonmode a_39362_63198# 0.31fF
C2339 a_5915_35943# a_12120_29941# 0.43fF
C2340 a_19807_28111# a_20635_29415# 0.89fF
C2341 a_12947_71576# a_16362_71230# 1.13fF
C2342 a_26402_59182# VDD 0.51fF
C2343 vcm_commonmode a_33430_9492# 0.87fF
C2344 m3_42368_72146# VDD 0.33fF
C2345 a_33338_23914# a_33430_23548# 0.32fF
C2346 a_7387_64239# VDD 0.86fF
C2347 a_12907_27023# a_38239_32375# 0.71fF
C2348 a_27535_30503# a_26523_29199# 0.37fF
C2349 a_8123_56399# a_2872_44111# 1.28fF
C2350 a_26402_11500# a_27406_11500# 0.97fF
C2351 a_34759_31029# VDD 3.18fF
C2352 vcm_commonmode a_49494_16520# 0.90fF
C2353 a_30418_64202# ctopp 3.59fF
C2354 ctopn a_35438_13508# 3.59fF
C2355 a_13909_41923# a_14293_41807# 1.71fF
C2356 a_2411_26133# config_2_in[3] 0.50fF
C2357 a_36442_72234# VDD 1.25fF
C2358 vcm_commonmode a_33338_59182# 0.31fF
C2359 a_39389_52271# a_12727_58255# 0.40fF
C2360 a_30326_66210# a_30418_66210# 0.32fF
C2361 a_4429_14191# a_5959_13621# 0.45fF
C2362 a_12516_7093# ctopp 3.23fF
C2363 a_8197_31599# a_10531_31055# 0.71fF
C2364 vcm_commonmode m3_16264_65118# 3.21fF
C2365 a_5831_39189# a_8491_41383# 2.72fF
C2366 a_43470_12504# VDD 0.51fF
C2367 a_23901_43132# VDD 1.05fF
C2368 a_44474_70226# a_44474_69222# 1.00fF
C2369 a_16955_52047# a_12355_65103# 0.40fF
C2370 a_5963_36585# a_7598_36103# 0.35fF
C2371 a_11067_47695# a_7571_26151# 0.99fF
C2372 a_37926_51727# VDD 0.44fF
C2373 vcm_commonmode a_41462_72234# 0.69fF
C2374 a_30418_24552# a_31422_24552# 0.97fF
C2375 a_27752_7638# a_12985_7663# 0.41fF
C2376 a_5211_24759# a_4798_23759# 0.79fF
C2377 a_4674_40277# a_5691_36727# 1.07fF
C2378 a_7939_30503# VDD 6.45fF
C2379 a_17507_52047# a_10687_52553# 1.09fF
C2380 a_18151_52263# a_4758_45369# 0.85fF
C2381 a_3843_13880# VDD 0.62fF
C2382 a_34763_47349# VDD 0.33fF
C2383 a_42374_19898# a_42466_19532# 0.32fF
C2384 a_38450_21540# VDD 0.51fF
C2385 vcm_commonmode a_41462_7484# 0.69fF
C2386 a_27406_62194# a_28410_62194# 0.97fF
C2387 a_43470_11500# a_43470_10496# 1.00fF
C2388 a_11602_25071# a_9751_25071# 0.48fF
C2389 a_47394_14878# a_47486_14512# 0.32fF
C2390 a_12191_37999# VDD 0.40fF
C2391 vcm_commonmode a_45386_21906# 0.31fF
C2392 a_39454_69222# ctopp 3.59fF
C2393 vcm_commonmode a_35438_64202# 0.87fF
C2394 a_8782_65015# a_3024_67191# 0.49fF
C2395 a_19720_7638# a_19374_7484# 0.34fF
C2396 a_2292_17179# a_3911_16065# 0.37fF
C2397 a_43470_17524# VDD 0.51fF
C2398 a_26310_20902# a_26402_20536# 0.32fF
C2399 a_27752_7638# a_27406_13508# 0.38fF
C2400 a_30418_60186# VDD 0.51fF
C2401 a_40458_55166# a_41462_55166# 0.97fF
C2402 a_8933_22583# VDD 2.05fF
C2403 vcm_commonmode a_22294_10862# 0.31fF
C2404 a_11067_66191# VDD 10.34fF
C2405 a_11067_46823# a_30052_32117# 1.51fF
C2406 a_12357_37999# a_13669_38517# 4.68fF
C2407 a_3417_31599# VDD 0.56fF
C2408 a_11619_56615# a_11887_19087# 0.84fF
C2409 a_37446_65206# ctopp 3.59fF
C2410 a_2787_32679# a_1799_29556# 0.83fF
C2411 a_32426_57174# a_33430_57174# 0.97fF
C2412 vcm_commonmode a_37354_60186# 0.31fF
C2413 a_35438_15516# a_36442_15516# 0.97fF
C2414 a_25321_29673# a_14926_31849# 0.40fF
C2415 a_8171_43541# VDD 0.47fF
C2416 a_12895_13967# VDD 7.04fF
C2417 a_6224_73095# a_6453_71855# 0.39fF
C2418 a_1586_69367# a_2843_71829# 0.88fF
C2419 a_35601_27497# a_35438_24552# 0.46fF
C2420 a_5682_69367# a_8491_57487# 0.75fF
C2421 a_1954_61677# a_1775_60663# 0.53fF
C2422 a_24987_36649# VDD 0.66fF
C2423 vcm_commonmode a_23390_19532# 0.87fF
C2424 a_1803_20719# a_4535_43567# 0.36fF
C2425 a_11067_46823# a_15607_46805# 0.80fF
C2426 a_33430_71230# a_34434_71230# 0.97fF
C2427 vcm_commonmode a_44474_69222# 0.87fF
C2428 a_4311_58229# VDD 0.38fF
C2429 a_45478_11500# a_46482_11500# 0.97fF
C2430 vcm_commonmode a_17274_15882# 0.33fF
C2431 a_9024_71427# VDD 0.45fF
C2432 a_49402_66210# a_49494_66210# 0.32fF
C2433 a_8197_31599# a_11812_30511# 0.58fF
C2434 vcm_commonmode m3_16264_12366# 3.21fF
C2435 a_20378_11500# VDD 0.51fF
C2436 a_15193_41781# VDD 1.03fF
C2437 a_1950_59887# a_8999_61493# 0.48fF
C2438 vcm_commonmode a_42466_65206# 0.87fF
C2439 ctopn a_9135_27239# 2.62fF
C2440 a_44474_18528# VDD 0.51fF
C2441 a_9314_69367# a_9063_71553# 0.34fF
C2442 a_28756_7638# a_28410_15516# 0.38fF
C2443 a_24394_24552# VDD 0.60fF
C2444 vcm_commonmode a_27314_11866# 0.31fF
C2445 ctopn a_42466_8488# 3.40fF
C2446 a_26310_12870# a_26402_12504# 0.32fF
C2447 a_44474_66210# ctopp 3.59fF
C2448 vcm_commonmode a_31330_24918# 0.31fF
C2449 a_16955_52047# ctopp 2.62fF
C2450 a_16863_29415# a_18979_30287# 1.01fF
C2451 a_4149_45743# VDD 0.63fF
C2452 a_17507_52047# a_21382_68218# 0.38fF
C2453 a_1591_18543# a_1895_18756# 0.62fF
C2454 a_21382_59182# a_21382_58178# 1.00fF
C2455 a_34434_55166# VDD 0.60fF
C2456 a_5497_63303# VDD 0.93fF
C2457 a_5363_30503# a_5915_30287# 0.74fF
C2458 a_46482_62194# a_47486_62194# 0.97fF
C2459 a_28305_28879# VDD 1.85fF
C2460 a_26402_57174# VDD 0.51fF
C2461 vcm_commonmode a_47486_14512# 0.87fF
C2462 a_14293_37455# VDD 1.05fF
C2463 vcm_commonmode a_26402_20536# 0.87fF
C2464 vcm_commonmode a_41370_55166# 0.30fF
C2465 a_49984_39288# VDD 0.59fF
C2466 a_17366_68218# a_18370_68218# 0.97fF
C2467 vcm_commonmode a_33338_57174# 0.31fF
C2468 a_5915_35943# a_11719_28023# 0.37fF
C2469 a_36717_47375# a_36442_71230# 0.38fF
C2470 a_45386_20902# a_45478_20536# 0.32fF
C2471 a_8491_27023# a_12985_7663# 0.41fF
C2472 VDD config_1_in[9] 1.03fF
C2473 a_1923_59583# a_2163_59585# 0.38fF
C2474 a_34342_63198# a_34434_63198# 0.32fF
C2475 a_12591_31029# VDD 0.45fF
C2476 a_21371_50959# a_17682_50095# 1.13fF
C2477 a_18151_52263# a_4191_33449# 0.34fF
C2478 a_25398_57174# a_25398_56170# 1.00fF
C2479 a_43362_28879# a_47486_61190# 0.38fF
C2480 a_19720_55394# a_19374_60186# 0.38fF
C2481 a_12907_56399# a_12981_59343# 0.34fF
C2482 vcm_commonmode a_49494_66210# 0.90fF
C2483 a_34251_52263# a_35438_67214# 0.38fF
C2484 a_5963_36585# a_7381_35407# 0.41fF
C2485 a_6831_63303# a_27509_47695# 0.47fF
C2486 a_21290_21906# a_21382_21540# 0.32fF
C2487 a_40458_62194# VDD 0.51fF
C2488 a_6372_38279# a_1761_32143# 0.90fF
C2489 a_4555_55233# VDD 0.49fF
C2490 vcm_commonmode a_26402_12504# 0.87fF
C2491 ctopn a_27406_9492# 3.58fF
C2492 a_12341_3311# a_22386_24552# 0.50fF
C2493 a_11710_58487# VDD 3.06fF
C2494 a_4811_34855# VDD 14.19fF
C2495 ctopn a_43470_16520# 3.59fF
C2496 a_21012_30761# a_22562_28023# 0.54fF
C2497 a_2021_17973# a_13835_43177# 2.01fF
C2498 vcm_commonmode a_47394_62194# 0.31fF
C2499 a_12907_56399# a_8123_56399# 1.48fF
C2500 a_17507_52047# a_21382_56170# 0.38fF
C2501 ctopn a_12546_22351# 3.23fF
C2502 a_21187_29415# a_26523_28111# 0.44fF
C2503 a_48490_15516# VDD 0.54fF
C2504 a_4563_32900# VDD 1.74fF
C2505 vcm_commonmode a_18278_68218# 0.31fF
C2506 a_28318_59182# a_28410_59182# 0.32fF
C2507 a_12869_2741# a_12341_3311# 0.70fF
C2508 a_7775_10625# a_7736_10499# 0.75fF
C2509 a_48490_63198# ctopp 3.49fF
C2510 a_46482_71230# VDD 0.58fF
C2511 a_43362_28879# a_12901_58799# 0.40fF
C2512 a_76180_38962# VDD 0.33fF
C2513 vcm_commonmode a_21382_21540# 0.87fF
C2514 a_11067_23759# a_12899_3855# 5.92fF
C2515 VDD config_2_in[0] 2.04fF
C2516 a_26310_17890# a_26402_17524# 0.32fF
C2517 a_36629_27791# a_36442_8488# 0.38fF
C2518 a_2011_34837# a_5079_35639# 0.34fF
C2519 a_42466_59182# ctopp 3.59fF
C2520 a_32951_27247# a_33430_22544# 0.38fF
C2521 a_32772_7638# a_32426_21540# 0.38fF
C2522 a_32426_64202# a_32426_63198# 1.23fF
C2523 a_45386_12870# a_45478_12504# 0.32fF
C2524 vcm_commonmode a_26402_17524# 0.87fF
C2525 a_18151_52263# a_12981_59343# 0.40fF
C2526 a_25398_13508# VDD 0.51fF
C2527 a_1950_59887# a_9513_65301# 0.52fF
C2528 a_3339_43023# a_1761_41935# 0.69fF
C2529 VDD config_2_in[10] 1.05fF
C2530 a_1770_14441# a_1803_19087# 1.82fF
C2531 a_24394_22544# a_24394_21540# 1.00fF
C2532 vcm_commonmode a_32334_13874# 0.31fF
C2533 a_11053_69135# VDD 0.88fF
C2534 a_31422_13508# a_32426_13508# 0.97fF
C2535 a_1761_22895# a_4701_43567# 0.59fF
C2536 a_1761_25071# a_12357_37999# 0.79fF
C2537 a_1761_44111# a_12549_44212# 0.63fF
C2538 a_3339_32463# a_2411_26133# 0.40fF
C2539 a_36442_68218# a_37446_68218# 0.97fF
C2540 vcm_commonmode a_18278_56170# 0.31fF
C2541 a_38557_32143# a_12516_7093# 0.40fF
C2542 a_39223_32463# a_39454_9492# 0.38fF
C2543 a_11067_47695# a_2872_44111# 1.27fF
C2544 a_12340_29967# VDD 0.34fF
C2545 a_17366_56170# a_18370_56170# 0.97fF
C2546 a_44474_57174# a_44474_56170# 1.00fF
C2547 a_47394_72234# VDD 0.61fF
C2548 vcm_commonmode a_47486_59182# 0.87fF
C2549 a_4119_70741# a_5190_59575# 1.23fF
C2550 ctopn a_17366_19532# 3.43fF
C2551 a_27752_7638# a_27406_7484# 0.34fF
C2552 a_1761_30511# a_12641_36596# 1.51fF
C2553 a_1761_37039# a_13669_35253# 1.24fF
C2554 a_13445_50639# VDD 1.01fF
C2555 a_13183_52047# a_17507_52047# 0.83fF
C2556 a_40366_21906# a_40458_21540# 0.32fF
C2557 a_10975_60975# VDD 0.37fF
C2558 a_13643_28327# a_17712_7638# 0.43fF
C2559 a_46482_60186# ctopp 3.59fF
C2560 a_6559_59663# a_7749_55535# 0.61fF
C2561 a_21382_58178# a_21382_57174# 1.00fF
C2562 a_49494_68218# VDD 1.14fF
C2563 vcm_commonmode a_27406_18528# 0.87fF
C2564 a_49402_7850# VDD 0.73fF
C2565 vcm_commonmode a_17274_61190# 0.33fF
C2566 a_28410_16520# a_28410_15516# 1.00fF
C2567 ctopn a_45478_22544# 3.58fF
C2568 a_2689_65103# a_3143_66972# 0.33fF
C2569 a_23736_7638# a_23390_8488# 0.38fF
C2570 a_47394_59182# a_47486_59182# 0.32fF
C2571 a_24413_39087# a_25133_37571# 0.33fF
C2572 a_6831_63303# a_28959_49783# 0.34fF
C2573 a_5363_30503# a_5915_35943# 0.31fF
C2574 a_3295_62083# a_3938_61493# 0.31fF
C2575 a_1952_60431# a_2959_47113# 2.14fF
C2576 a_17274_10862# a_17366_10496# 0.32fF
C2577 a_18370_62194# ctopp 3.58fF
C2578 a_22448_38341# VDD 1.78fF
C2579 vcm_commonmode a_18370_55166# 0.84fF
C2580 a_75199_40594# VDD 0.48fF
C2581 a_11067_67279# a_11999_67477# 0.37fF
C2582 a_45386_17890# a_45478_17524# 0.32fF
C2583 a_13669_35253# a_1761_32143# 4.53fF
C2584 a_20156_49667# VDD 0.31fF
C2585 vcm_commonmode a_21290_70226# 0.31fF
C2586 a_5671_21495# a_2411_18517# 0.48fF
C2587 a_38358_58178# vcm_commonmode 0.31fF
C2588 a_32334_60186# a_32426_60186# 0.32fF
C2589 vcm_commonmode a_36442_10496# 0.87fF
C2590 a_12161_31849# VDD 0.97fF
C2591 ctopn a_41462_14512# 3.59fF
C2592 a_23195_29967# a_17712_7638# 0.43fF
C2593 a_12725_44527# a_13909_39747# 2.29fF
C2594 a_2322_72631# VDD 0.62fF
C2595 a_24394_71230# ctopp 3.40fF
C2596 ctopn a_20378_20536# 3.59fF
C2597 a_25398_7484# m3_25300_7346# 2.80fF
C2598 a_27314_18894# a_27406_18528# 0.32fF
C2599 a_2411_18517# a_2292_17179# 1.04fF
C2600 a_43470_22544# a_43470_21540# 1.00fF
C2601 a_16362_62194# VDD 2.48fF
C2602 a_20635_29415# a_37699_27221# 0.62fF
C2603 a_49494_56170# VDD 1.14fF
C2604 a_5079_35639# VDD 0.47fF
C2605 a_36613_48169# a_37446_55166# 0.46fF
C2606 a_6649_25615# a_5087_29423# 0.41fF
C2607 a_32426_8488# VDD 0.58fF
C2608 vcm_commonmode a_23390_62194# 0.87fF
C2609 a_22386_68218# a_22386_67214# 1.00fF
C2610 a_21371_52263# a_26402_63198# 0.42fF
C2611 ctopn a_46482_23548# 3.40fF
C2612 a_2163_57853# VDD 0.49fF
C2613 a_3339_43023# a_1761_25071# 0.40fF
C2614 a_12901_58799# a_16362_59182# 19.89fF
C2615 vcm_commonmode a_39362_8854# 0.31fF
C2616 m3_29316_7346# VDD 0.40fF
C2617 a_24740_7638# a_12895_13967# 0.41fF
C2618 vcm_commonmode a_31422_15516# 0.87fF
C2619 ctopn a_20378_12504# 3.59fF
C2620 a_3143_22364# a_4571_26677# 0.42fF
C2621 a_41967_31375# a_42466_23548# 0.38fF
C2622 a_42466_57174# ctopp 3.58fF
C2623 a_36442_56170# a_37446_56170# 0.97fF
C2624 a_39299_48783# a_10515_22671# 0.40fF
C2625 a_18811_39141# VDD 0.86fF
C2626 a_20715_41245# VDD 1.38fF
C2627 a_2689_65103# a_3668_56311# 0.36fF
C2628 ctopn a_32951_27247# 2.67fF
C2629 a_28410_72234# a_29414_72234# 0.97fF
C2630 vcm_commonmode a_29414_71230# 0.86fF
C2631 a_40675_27791# a_12727_15529# 0.41fF
C2632 a_48490_61190# VDD 0.54fF
C2633 a_18278_55166# a_18370_55166# 0.33fF
C2634 a_19374_8488# a_20378_8488# 0.97fF
C2635 vcm_commonmode a_41462_11500# 0.87fF
C2636 a_36797_27497# a_12546_22351# 0.41fF
C2637 a_3325_18543# a_5535_18012# 0.31fF
C2638 a_20378_67214# VDD 0.51fF
C2639 a_47486_16520# a_47486_15516# 1.00fF
C2640 vcm_commonmode a_45478_24552# 0.84fF
C2641 a_2292_43291# a_1591_45205# 0.34fF
C2642 a_20378_70226# a_21382_70226# 0.97fF
C2643 vcm_commonmode a_27314_67214# 0.31fF
C2644 a_19720_7638# a_19374_11500# 0.38fF
C2645 a_32426_19532# a_32426_18528# 1.00fF
C2646 a_3987_19623# a_7059_24135# 0.83fF
C2647 a_37446_58178# a_38450_58178# 0.97fF
C2648 a_37919_28111# a_38450_18528# 0.38fF
C2649 a_36350_10862# a_36442_10496# 0.32fF
C2650 a_11902_27497# VDD 3.41fF
C2651 a_24740_7638# a_24394_24552# 0.46fF
C2652 a_3972_25615# a_4333_22895# 0.41fF
C2653 a_34639_37737# VDD 0.60fF
C2654 a_27406_68218# ctopp 3.59fF
C2655 ctopn a_20378_17524# 3.59fF
C2656 a_34759_31029# a_38436_29941# 0.33fF
C2657 a_17366_9492# VDD 0.58fF
C2658 vcm_commonmode a_47486_57174# 0.87fF
C2659 a_33430_16520# VDD 0.51fF
C2660 a_13183_52047# a_17366_70226# 0.38fF
C2661 a_18370_60186# a_18370_59182# 1.00fF
C2662 vcm_commonmode a_24302_9858# 0.31fF
C2663 m2_15446_6268# VDD 0.59fF
C2664 a_43175_28335# a_46482_20536# 0.38fF
C2665 a_8295_47388# a_11619_3303# 0.56fF
C2666 a_22294_11866# a_22386_11500# 0.32fF
C2667 a_29926_30511# VDD 1.09fF
C2668 vcm_commonmode a_40366_16886# 0.31fF
C2669 a_15459_41781# a_12713_41923# 0.38fF
C2670 a_29414_72234# VDD 1.60fF
C2671 a_28547_51175# a_12727_58255# 0.40fF
C2672 a_27406_15516# a_27406_14512# 1.00fF
C2673 a_46390_18894# a_46482_18528# 0.32fF
C2674 ctopn a_43175_28335# 2.63fF
C2675 a_3339_43023# a_4578_40455# 0.33fF
C2676 a_13669_37429# a_1761_31055# 1.26fF
C2677 a_2216_28309# a_1761_30511# 0.90fF
C2678 vcm_commonmode a_34434_72234# 0.69fF
C2679 a_35438_61190# a_36442_61190# 0.97fF
C2680 a_26748_7638# a_11067_21583# 0.41fF
C2681 a_26310_24918# a_26402_24552# 0.32fF
C2682 a_4191_33449# a_1761_34319# 0.48fF
C2683 a_12907_56399# a_11067_47695# 3.03fF
C2684 a_25398_7484# VDD 1.59fF
C2685 a_41462_68218# a_41462_67214# 1.00fF
C2686 a_12727_13353# a_16746_15514# 0.41fF
C2687 vcm_commonmode a_32426_68218# 0.87fF
C2688 a_12355_15055# a_5363_30503# 0.83fF
C2689 a_4379_18756# a_4241_18543# 0.56fF
C2690 a_43175_28335# a_46482_12504# 0.38fF
C2691 a_19374_64202# VDD 0.51fF
C2692 a_20359_29199# a_41597_29967# 0.66fF
C2693 a_23298_62194# a_23390_62194# 0.32fF
C2694 a_13239_29575# VDD 1.15fF
C2695 a_27406_56170# ctopp 3.40fF
C2696 ctopn a_21382_18528# 3.59fF
C2697 a_48490_72234# m3_48392_72146# 2.80fF
C2698 a_8375_40847# VDD 0.40fF
C2699 vcm_commonmode a_26310_64202# 0.31fF
C2700 a_26402_69222# a_26402_68218# 1.00fF
C2701 a_13005_35823# a_19594_35823# 1.29fF
C2702 a_12663_35431# a_13669_35253# 0.50fF
C2703 a_41872_29423# a_43470_72234# 0.34fF
C2704 a_38450_8488# a_39454_8488# 0.97fF
C2705 a_36350_55166# a_36442_55166# 0.32fF
C2706 a_8491_57487# a_8453_51727# 0.38fF
C2707 a_21187_29415# a_35815_31751# 1.40fF
C2708 a_6831_63303# a_7097_63151# 0.35fF
C2709 a_11067_63143# a_10515_63143# 1.90fF
C2710 a_42941_32143# VDD 0.44fF
C2711 a_28318_57174# a_28410_57174# 0.32fF
C2712 a_31330_15882# a_31422_15516# 0.32fF
C2713 a_36116_44765# VDD 1.25fF
C2714 a_39454_70226# a_40458_70226# 0.97fF
C2715 a_12516_7093# a_16746_69224# 2.28fF
C2716 a_14293_37455# a_20827_37737# 0.37fF
C2717 a_5135_19061# VDD 0.50fF
C2718 a_43175_28335# a_46482_17524# 0.38fF
C2719 a_40491_27247# a_43470_18528# 0.38fF
C2720 a_7295_44647# a_30565_30199# 2.25fF
C2721 vcm_commonmode a_46482_13508# 0.87fF
C2722 a_26402_61190# ctopp 3.59fF
C2723 ctopn a_30418_10496# 3.59fF
C2724 a_28410_69222# VDD 0.51fF
C2725 a_12889_35537# VDD 0.96fF
C2726 a_18611_52047# a_12869_2741# 0.44fF
C2727 a_18151_52263# a_11067_47695# 0.69fF
C2728 a_11067_23759# a_9503_26151# 11.31fF
C2729 a_20378_16520# a_21382_16520# 0.97fF
C2730 vcm_commonmode a_32426_56170# 0.87fF
C2731 a_2606_41079# a_17280_48695# 0.30fF
C2732 vcm_commonmode a_35346_69222# 0.31fF
C2733 a_29322_71230# a_29414_71230# 0.32fF
C2734 a_3339_43023# a_2787_32679# 0.44fF
C2735 a_37446_60186# a_37446_59182# 1.00fF
C2736 a_35438_22544# VDD 0.51fF
C2737 a_10975_66407# a_17488_48731# 1.48fF
C2738 a_1952_60431# a_1823_53885# 0.35fF
C2739 a_26402_65206# VDD 0.51fF
C2740 a_26402_63198# a_26402_62194# 1.00fF
C2741 a_41370_11866# a_41462_11500# 0.32fF
C2742 a_8531_70543# a_17039_51157# 1.24fF
C2743 a_46482_15516# a_46482_14512# 1.00fF
C2744 vcm_commonmode a_42374_22910# 0.31fF
C2745 a_30418_70226# ctopp 3.58fF
C2746 a_19743_42359# VDD 0.61fF
C2747 vcm_commonmode a_33338_65206# 0.31fF
C2748 ctopn a_43270_27791# 2.63fF
C2749 a_37423_51335# VDD 0.36fF
C2750 a_31422_9492# a_31422_8488# 1.00fF
C2751 a_45386_24918# a_45478_24552# 0.32fF
C2752 ctopn a_25398_15516# 3.59fF
C2753 a_23395_52047# a_2872_44111# 0.55fF
C2754 a_26402_67214# a_27406_67214# 0.97fF
C2755 vcm_commonmode a_31422_61190# 0.87fF
C2756 a_17711_32385# a_17672_32259# 0.46fF
C2757 a_31422_14512# VDD 0.51fF
C2758 a_12516_7093# a_16746_70228# 0.41fF
C2759 a_26310_55166# VDD 0.35fF
C2760 a_6816_19355# a_5535_18012# 0.85fF
C2761 a_5963_20149# a_4792_20443# 1.06fF
C2762 a_11067_46823# a_28841_29575# 0.53fF
C2763 a_42374_62194# a_42466_62194# 0.32fF
C2764 vcm_commonmode a_38358_14878# 0.31fF
C2765 ctopn a_35438_11500# 3.59fF
C2766 a_12473_37429# VDD 7.11fF
C2767 vcm_commonmode a_17274_20902# 0.33fF
C2768 vcm_commonmode a_32426_55166# 0.84fF
C2769 a_20713_40193# VDD 1.75fF
C2770 a_45478_69222# a_45478_68218# 1.00fF
C2771 a_1761_32143# a_23567_35507# 0.47fF
C2772 a_4495_35925# a_4903_31849# 1.17fF
C2773 a_20635_29415# VDD 12.62fF
C2774 a_39299_48783# a_12901_66665# 0.40fF
C2775 vcm_commonmode a_35438_70226# 0.87fF
C2776 a_28547_51175# a_32426_71230# 0.38fF
C2777 a_35438_8488# a_35438_7484# 1.00fF
C2778 a_36442_23548# VDD 0.52fF
C2779 a_19374_58178# ctopp 3.59fF
C2780 a_28756_7638# a_28410_20536# 0.38fF
C2781 a_33430_66210# VDD 0.51fF
C2782 vcm_commonmode a_16746_16518# 5.36fF
C2783 a_1952_60431# a_2589_55535# 0.35fF
C2784 a_47394_57174# a_47486_57174# 0.32fF
C2785 a_41872_29423# a_43470_61190# 0.38fF
C2786 vcm_commonmode a_43378_23914# 0.31fF
C2787 vcm_commonmode a_40366_66210# 0.31fF
C2788 a_31768_55394# a_31422_67214# 0.38fF
C2789 a_28410_58178# a_29414_58178# 0.97fF
C2790 a_1761_37039# a_12473_36341# 1.64fF
C2791 a_45478_19532# VDD 0.51fF
C2792 a_16746_21538# a_12985_7663# 2.28fF
C2793 a_23390_9492# a_24394_9492# 0.97fF
C2794 a_33430_55166# m3_33332_55078# 1.39fF
C2795 vcm_commonmode a_17274_12870# 0.33fF
C2796 a_4647_63937# a_4608_63811# 0.75fF
C2797 a_24394_13508# a_24394_12504# 1.00fF
C2798 a_36442_67214# ctopp 3.59fF
C2799 a_5831_39189# a_4314_40821# 0.57fF
C2800 a_2021_17973# a_1803_19087# 1.38fF
C2801 a_39454_16520# a_40458_16520# 0.97fF
C2802 a_11067_67279# a_39223_32463# 0.41fF
C2803 a_48398_71230# a_48490_71230# 0.32fF
C2804 a_29760_7638# a_29414_13508# 0.38fF
C2805 a_28756_7638# a_28410_12504# 0.38fF
C2806 a_27752_7638# a_27406_11500# 0.38fF
C2807 a_11067_46823# a_30565_30199# 0.79fF
C2808 a_45478_63198# a_45478_62194# 1.00fF
C2809 a_19807_28111# a_7841_12167# 3.70fF
C2810 a_39222_48169# a_12901_58799# 0.40fF
C2811 vcm_commonmode a_24394_58178# 0.87fF
C2812 a_49402_11866# VDD 0.31fF
C2813 a_13835_41001# VDD 0.48fF
C2814 a_35196_35425# a_1761_35407# 0.32fF
C2815 a_17039_51157# a_16587_49007# 0.33fF
C2816 a_34342_72234# a_34434_72234# 0.32fF
C2817 a_4187_60673# VDD 0.45fF
C2818 a_1867_23983# VDD 0.35fF
C2819 a_16510_8760# a_12727_15529# 1.08fF
C2820 a_49494_62194# m3_49396_62106# 2.78fF
C2821 a_12158_32143# VDD 0.38fF
C2822 vcm_commonmode a_17274_17890# 0.33fF
C2823 a_13390_29575# a_18307_27791# 0.62fF
C2824 a_12631_28585# a_10873_27497# 0.34fF
C2825 a_45478_67214# a_46482_67214# 0.97fF
C2826 a_11067_66191# a_9307_30663# 1.09fF
C2827 a_41261_28335# a_3339_43023# 0.98fF
C2828 a_12725_44527# VDD 7.52fF
C2829 vcm_commonmode a_41462_67214# 0.87fF
C2830 a_48490_20536# VDD 0.54fF
C2831 a_37459_51183# a_35568_49525# 0.81fF
C2832 a_4036_54421# VDD 0.35fF
C2833 a_7755_74581# a_6224_73095# 0.63fF
C2834 a_28756_7638# a_28410_17524# 0.38fF
C2835 a_37446_63198# VDD 0.57fF
C2836 a_25787_28327# a_18979_30287# 0.46fF
C2837 a_43269_29967# a_11067_21583# 0.41fF
C2838 a_27314_13874# a_27406_13508# 0.32fF
C2839 a_7841_12167# a_7377_18012# 0.35fF
C2840 a_1591_29973# a_1757_29973# 0.58fF
C2841 vcm_commonmode a_44382_63198# 0.31fF
C2842 a_41872_29423# a_12355_15055# 0.40fF
C2843 a_32334_68218# a_32426_68218# 0.32fF
C2844 a_4287_48634# VDD 0.58fF
C2845 a_31768_55394# a_12516_7093# 0.40fF
C2846 a_48490_72234# a_48490_71230# 1.00fF
C2847 a_31422_59182# VDD 0.51fF
C2848 a_2021_22325# a_3143_22364# 0.59fF
C2849 a_31422_7484# a_32426_7484# 0.97fF
C2850 vcm_commonmode a_38450_9492# 0.87fF
C2851 a_45478_24552# m3_45380_24414# 2.81fF
C2852 a_35438_64202# ctopp 3.59fF
C2853 ctopn a_40458_13508# 3.59fF
C2854 a_6835_46823# a_3339_43023# 0.60fF
C2855 a_40366_72234# VDD 0.62fF
C2856 vcm_commonmode a_38358_59182# 0.31fF
C2857 a_13183_52047# a_10515_22671# 0.41fF
C2858 vcm_commonmode a_18370_22544# 0.88fF
C2859 a_48490_12504# VDD 0.54fF
C2860 a_30415_43177# VDD 0.63fF
C2861 a_11803_55311# a_12983_63151# 1.06fF
C2862 a_28881_52271# a_36464_49783# 0.52fF
C2863 a_8539_18231# VDD 0.33fF
C2864 a_5909_51433# VDD 0.47fF
C2865 a_5877_70197# a_11049_71855# 0.59fF
C2866 a_11067_63143# a_7571_26151# 1.56fF
C2867 a_5363_30503# a_7939_30503# 1.01fF
C2868 a_42466_9492# a_43470_9492# 0.97fF
C2869 a_16863_29415# a_16510_8760# 1.02fF
C2870 a_25398_64202# a_26402_64202# 0.97fF
C2871 a_43470_13508# a_43470_12504# 1.00fF
C2872 a_24515_34789# VDD 1.03fF
C2873 vcm_commonmode a_18278_18894# 0.31fF
C2874 a_6243_30662# a_5993_32687# 0.47fF
C2875 a_10515_22671# a_7571_29199# 0.43fF
C2876 a_43470_21540# VDD 0.51fF
C2877 vcm_commonmode a_46482_7484# 0.69fF
C2878 a_22386_22544# a_23390_22544# 0.97fF
C2879 a_24959_30503# a_34759_31029# 0.45fF
C2880 a_10680_52245# a_10687_52553# 0.86fF
C2881 a_44474_69222# ctopp 3.59fF
C2882 a_2004_42453# config_2_in[7] 1.02fF
C2883 a_20946_30669# a_21057_30669# 0.47fF
C2884 a_20378_10496# VDD 0.51fF
C2885 a_22132_40865# VDD 1.70fF
C2886 vcm_commonmode a_40458_64202# 0.87fF
C2887 a_1959_68053# a_2125_68053# 0.72fF
C2888 ctopn a_12341_3311# 2.62fF
C2889 a_38115_52263# a_37557_32463# 9.74fF
C2890 a_48490_17524# VDD 0.54fF
C2891 a_9301_49557# VDD 0.33fF
C2892 a_35438_60186# VDD 0.51fF
C2893 a_3339_43023# a_6559_22671# 0.66fF
C2894 vcm_commonmode a_27314_10862# 0.31fF
C2895 a_27535_30503# a_33798_31145# 0.41fF
C2896 a_18328_31573# VDD 0.34fF
C2897 a_42466_65206# ctopp 3.59fF
C2898 a_15661_29199# a_20685_28335# 0.35fF
C2899 a_2163_73085# VDD 0.53fF
C2900 vcm_commonmode a_42374_60186# 0.31fF
C2901 a_33430_67214# a_33430_66210# 1.00fF
C2902 vcm_commonmode a_19374_23548# 0.87fF
C2903 a_18370_7484# m3_18272_7346# 2.80fF
C2904 a_14646_29423# a_19626_31751# 1.27fF
C2905 a_6863_42692# a_5831_39189# 0.38fF
C2906 vcm_commonmode a_16746_66212# 5.36fF
C2907 a_2012_33927# a_2011_34837# 0.52fF
C2908 a_16219_51183# a_17039_51157# 0.34fF
C2909 a_2971_73493# a_3137_73493# 0.75fF
C2910 a_8003_72917# a_9353_72399# 0.70fF
C2911 a_6831_63303# a_28524_47919# 0.37fF
C2912 a_29414_65206# a_29414_64202# 1.00fF
C2913 a_46390_13874# a_46482_13508# 0.32fF
C2914 a_35463_36415# VDD 0.86fF
C2915 vcm_commonmode a_28410_19532# 0.87fF
C2916 ctopn a_12985_16367# 3.23fF
C2917 a_1761_22895# a_1803_19087# 0.72fF
C2918 a_17599_52263# a_22386_63198# 0.42fF
C2919 a_41261_28335# a_12257_56623# 0.40fF
C2920 a_1761_34319# a_11067_23759# 0.33fF
C2921 a_20635_29415# a_34482_29941# 0.42fF
C2922 a_16863_29415# a_18703_29199# 6.00fF
C2923 a_1761_52815# a_2021_17973# 1.16fF
C2924 vcm_commonmode a_49494_69222# 0.91fF
C2925 a_11080_58229# VDD 0.51fF
C2926 a_7050_53333# a_7217_53047# 0.66fF
C2927 a_2473_34293# start_conversion_in 0.36fF
C2928 a_10515_22671# a_12546_22351# 0.67fF
C2929 a_23390_23548# a_23390_22544# 1.00fF
C2930 a_37527_29397# VDD 1.05fF
C2931 vcm_commonmode a_22294_15882# 0.31fF
C2932 a_8583_33551# a_42709_29199# 0.39fF
C2933 a_32334_56170# a_32426_56170# 0.32fF
C2934 a_36613_48169# a_10515_22671# 0.40fF
C2935 a_17366_66210# a_17366_65206# 1.00fF
C2936 a_18370_14512# a_19374_14512# 0.97fF
C2937 a_14926_31849# a_17554_30663# 0.47fF
C2938 a_2787_30503# a_13390_29575# 0.33fF
C2939 a_25398_11500# VDD 0.51fF
C2940 a_5880_41641# VDD 0.47fF
C2941 a_34434_69222# a_35438_69222# 0.97fF
C2942 vcm_commonmode a_47486_65206# 0.87fF
C2943 a_12473_36341# a_12663_35431# 4.04fF
C2944 a_49494_18528# VDD 1.12fF
C2945 a_5147_50943# VDD 0.41fF
C2946 vcm_commonmode a_20286_71230# 0.31fF
C2947 a_29414_61190# a_29414_60186# 1.00fF
C2948 a_29414_24552# VDD 0.60fF
C2949 vcm_commonmode a_32334_11866# 0.31fF
C2950 ctopn a_47486_8488# 3.39fF
C2951 a_44474_64202# a_45478_64202# 0.97fF
C2952 a_12671_43222# a_12473_42869# 0.30fF
C2953 vcm_commonmode a_36350_24918# 0.31fF
C2954 a_1761_50639# a_2021_17973# 0.88fF
C2955 a_39454_55166# VDD 0.60fF
C2956 a_2959_47113# a_28881_52271# 0.81fF
C2957 a_41462_22544# a_42466_22544# 0.97fF
C2958 a_31422_57174# VDD 0.51fF
C2959 a_9503_26151# a_8491_27023# 3.73fF
C2960 a_29927_29199# a_7841_12167# 2.57fF
C2961 a_32426_65206# a_33430_65206# 0.97fF
C2962 a_7387_64239# a_4339_64521# 0.34fF
C2963 vcm_commonmode a_31422_20536# 0.87fF
C2964 vcm_commonmode a_46390_55166# 0.30fF
C2965 a_6927_39215# VDD 0.32fF
C2966 vcm_commonmode a_20378_63198# 0.92fF
C2967 a_29760_7638# a_29414_7484# 0.34fF
C2968 a_28410_17524# a_28410_16520# 1.00fF
C2969 vcm_commonmode a_38358_57174# 0.31fF
C2970 a_4119_70741# a_3143_66972# 0.84fF
C2971 a_1689_10396# a_3325_18543# 0.91fF
C2972 a_2411_19605# a_1591_21807# 0.52fF
C2973 a_23390_23548# a_24394_23548# 0.97fF
C2974 a_9643_63125# a_7523_62581# 0.34fF
C2975 ctopn a_16746_13506# 1.68fF
C2976 a_22386_72234# VDD 1.40fF
C2977 a_20378_66210# a_21382_66210# 0.97fF
C2978 a_21371_50959# a_12727_58255# 0.40fF
C2979 a_1768_16367# config_1_in[14] 0.47fF
C2980 a_23395_32463# a_34759_31029# 1.51fF
C2981 a_4674_40277# a_3339_32463# 0.71fF
C2982 a_4119_70741# a_1823_65853# 0.38fF
C2983 a_9319_69141# a_9485_69141# 0.72fF
C2984 a_13123_38231# a_13669_35253# 2.04fF
C2985 a_2872_44111# a_2606_41079# 0.72fF
C2986 a_14985_51701# VDD 1.66fF
C2987 vcm_commonmode a_27406_72234# 0.69fF
C2988 a_45478_62194# VDD 0.51fF
C2989 a_31330_61190# a_31422_61190# 0.32fF
C2990 a_6138_54599# VDD 0.50fF
C2991 vcm_commonmode a_31422_12504# 0.87fF
C2992 ctopn a_32426_9492# 3.58fF
C2993 a_26748_7638# a_12546_22351# 0.41fF
C2994 a_12727_67753# VDD 7.19fF
C2995 a_48490_65206# a_48490_64202# 1.00fF
C2996 ctopn a_48490_16520# 3.43fF
C2997 a_16270_7850# VDD 0.73fF
C2998 vcm_commonmode a_23298_68218# 0.31fF
C2999 a_20378_71230# a_20378_70226# 1.00fF
C3000 a_32426_19532# a_33430_19532# 0.97fF
C3001 a_42466_23548# a_42466_22544# 1.00fF
C3002 a_8531_70543# a_30928_49007# 0.41fF
C3003 a_36442_66210# a_36442_65206# 1.00fF
C3004 a_37446_14512# a_38450_14512# 0.97fF
C3005 a_2012_33927# VDD 11.58fF
C3006 vcm_commonmode a_26402_21540# 0.87fF
C3007 a_4503_10687# VDD 0.44fF
C3008 vcm_commonmode a_16362_64202# 4.48fF
C3009 vcm_commonmode a_44474_58178# 0.87fF
C3010 a_12549_35836# a_15968_36061# 1.90fF
C3011 a_19885_50095# VDD 0.46fF
C3012 a_13183_52047# a_12901_66665# 0.40fF
C3013 a_25744_7638# a_12727_15529# 0.41fF
C3014 a_48490_61190# a_48490_60186# 1.00fF
C3015 a_34342_8854# a_34434_8488# 0.32fF
C3016 a_32334_55166# a_32426_55166# 0.33fF
C3017 a_47486_59182# ctopp 3.58fF
C3018 a_23736_7638# a_12899_10927# 0.41fF
C3019 a_11067_23759# a_12727_13353# 0.36fF
C3020 a_49402_67214# VDD 0.31fF
C3021 vcm_commonmode a_31422_17524# 0.87fF
C3022 a_6224_73095# VDD 3.56fF
C3023 vcm_commonmode a_18370_60186# 0.88fF
C3024 a_30418_13508# VDD 0.51fF
C3025 a_35346_70226# a_35438_70226# 0.32fF
C3026 a_4119_70741# a_3668_56311# 1.08fF
C3027 a_2419_48783# a_9779_47919# 0.71fF
C3028 a_8491_27023# a_9642_10357# 0.43fF
C3029 a_13123_38231# a_13835_36649# 0.34fF
C3030 a_2847_19605# VDD 0.47fF
C3031 a_18127_35797# a_1761_35407# 1.34fF
C3032 a_34434_62194# a_34434_61190# 1.00fF
C3033 a_25398_10496# a_25398_9492# 1.00fF
C3034 a_16746_56172# VDD 33.41fF
C3035 vcm_commonmode a_37354_13874# 0.31fF
C3036 a_41289_36893# VDD 0.99fF
C3037 a_47486_17524# a_47486_16520# 1.00fF
C3038 a_16362_16520# a_16746_16518# 2.28fF
C3039 vcm_commonmode a_23298_56170# 0.31fF
C3040 a_2926_15253# VDD 0.38fF
C3041 a_34434_20536# a_34434_19532# 1.00fF
C3042 a_11067_63143# a_2872_44111# 0.79fF
C3043 a_42466_23548# a_43470_23548# 0.97fF
C3044 a_8933_22583# a_9955_21807# 0.82fF
C3045 a_3339_32463# a_7862_34025# 0.36fF
C3046 ctopp a_18370_55166# 0.57fF
C3047 a_39454_66210# a_40458_66210# 0.97fF
C3048 a_1923_59583# a_6515_62037# 0.43fF
C3049 a_4351_67279# a_2959_47113# 0.30fF
C3050 ctopn a_22386_19532# 3.59fF
C3051 a_4811_34855# a_23051_28023# 0.72fF
C3052 a_1761_47919# a_1761_22895# 1.12fF
C3053 a_5601_11471# VDD 0.49fF
C3054 a_41261_28335# a_10975_66407# 0.40fF
C3055 a_11067_21583# a_12985_19087# 0.40fF
C3056 a_36797_27497# a_12985_16367# 0.41fF
C3057 a_2840_66103# a_5135_50069# 0.47fF
C3058 a_7444_34025# VDD 0.46fF
C3059 vcm_commonmode a_32426_18528# 0.87fF
C3060 ctopn a_16362_15516# 1.35fF
C3061 a_16955_52047# a_2872_44111# 0.57fF
C3062 a_11067_23759# a_10515_23975# 0.39fF
C3063 a_22294_67214# a_22386_67214# 0.32fF
C3064 vcm_commonmode a_22294_61190# 0.31fF
C3065 a_2411_18517# a_11455_12157# 0.34fF
C3066 a_13183_52047# a_10680_52245# 0.32fF
C3067 a_39454_71230# a_39454_70226# 1.00fF
C3068 a_12899_2767# VDD 6.08fF
C3069 a_23390_62194# ctopp 3.59fF
C3070 a_4571_26677# a_4351_26703# 0.37fF
C3071 a_3339_43023# a_4571_26677# 1.52fF
C3072 a_19374_70226# VDD 0.51fF
C3073 a_32795_38053# VDD 0.87fF
C3074 a_11067_67279# a_42718_27497# 0.41fF
C3075 a_10975_66407# a_6835_46823# 0.89fF
C3076 vcm_commonmode a_23390_55166# 0.84fF
C3077 a_2052_38377# VDD 0.52fF
C3078 a_12899_11471# a_16746_16518# 0.41fF
C3079 a_3983_16617# VDD 0.59fF
C3080 a_36613_48169# a_12901_66665# 0.40fF
C3081 a_28756_55394# a_28410_71230# 0.38fF
C3082 vcm_commonmode a_26310_70226# 0.31fF
C3083 a_35438_20536# a_36442_20536# 0.97fF
C3084 a_43378_58178# vcm_commonmode 0.31fF
C3085 a_8273_42479# a_8739_28879# 0.47fF
C3086 vcm_commonmode a_41462_10496# 0.87fF
C3087 a_24394_63198# a_25398_63198# 0.97fF
C3088 a_20773_31849# VDD 0.61fF
C3089 a_11067_13095# a_12341_3311# 1.50fF
C3090 ctopn a_46482_14512# 3.59fF
C3091 a_1761_43567# a_32121_40741# 0.41fF
C3092 a_39389_52271# a_39454_61190# 0.38fF
C3093 a_29414_71230# ctopp 3.40fF
C3094 ctopn a_25398_20536# 3.59fF
C3095 a_2787_30503# a_10531_31055# 1.40fF
C3096 a_23395_52047# a_27406_67214# 0.38fF
C3097 a_19720_7638# a_19374_10496# 0.38fF
C3098 a_24302_58178# a_24394_58178# 0.32fF
C3099 a_1591_64239# a_1591_63151# 4.20fF
C3100 a_41967_31375# a_42466_14512# 0.38fF
C3101 a_17712_7638# a_12877_16911# 0.40fF
C3102 a_22291_29415# a_28963_28853# 0.42fF
C3103 a_44474_10496# a_44474_9492# 1.00fF
C3104 a_19282_9858# a_19374_9492# 0.32fF
C3105 a_10964_25615# VDD 0.95fF
C3106 a_22843_29415# a_4811_34855# 0.48fF
C3107 a_15069_35805# VDD 0.95fF
C3108 a_37446_8488# VDD 0.58fF
C3109 a_1761_22895# a_32695_43455# 0.76fF
C3110 vcm_commonmode a_28410_62194# 0.87fF
C3111 a_35346_16886# a_35438_16520# 0.32fF
C3112 a_22351_47893# VDD 0.65fF
C3113 a_12907_56399# a_12516_7093# 0.78fF
C3114 a_18370_59182# a_19374_59182# 0.97fF
C3115 a_4839_21495# VDD 0.59fF
C3116 vcm_commonmode a_44382_8854# 0.31fF
C3117 a_10975_66407# a_6559_22671# 0.37fF
C3118 vcm_commonmode a_36442_15516# 0.87fF
C3119 ctopn a_25398_12504# 3.59fF
C3120 a_47486_57174# ctopp 3.57fF
C3121 a_25787_28327# a_12901_58799# 0.40fF
C3122 a_26447_39141# VDD 1.05fF
C3123 a_28943_42089# VDD 0.61fF
C3124 vcm_commonmode a_34434_71230# 0.86fF
C3125 a_33430_21540# a_33430_20536# 1.00fF
C3126 a_1761_27791# a_15011_34717# 0.88fF
C3127 vcm_commonmode a_46482_11500# 0.87fF
C3128 a_20378_24552# a_20378_23548# 1.00fF
C3129 a_3339_43023# a_5963_20149# 0.42fF
C3130 a_25398_67214# VDD 0.51fF
C3131 a_35438_12504# a_36442_12504# 0.97fF
C3132 a_12412_32143# VDD 0.56fF
C3133 a_41370_67214# a_41462_67214# 0.32fF
C3134 a_34251_52263# a_3339_43023# 5.37fF
C3135 ctopn a_20378_21540# 3.59fF
C3136 vcm_commonmode a_32334_67214# 0.31fF
C3137 a_2451_72373# a_8575_74853# 0.97fF
C3138 a_6559_59879# a_4215_51157# 1.13fF
C3139 a_27752_7638# a_12727_13353# 0.41fF
C3140 a_39673_28111# a_40458_18528# 0.38fF
C3141 a_43269_29967# a_12546_22351# 0.41fF
C3142 a_36717_47375# a_36442_58178# 0.38fF
C3143 a_1761_35951# VDD 0.54fF
C3144 a_32426_68218# ctopp 3.59fF
C3145 ctopn a_25398_17524# 3.59fF
C3146 a_22386_9492# VDD 0.51fF
C3147 a_1689_10396# a_1761_43567# 1.14fF
C3148 a_1761_25071# a_1803_20719# 1.02fF
C3149 a_36717_47375# a_12355_15055# 0.40fF
C3150 a_11067_67279# a_7862_34025# 1.20fF
C3151 a_38450_16520# VDD 0.51fF
C3152 a_18151_52263# a_12516_7093# 0.47fF
C3153 a_44474_72234# a_44474_71230# 1.00fF
C3154 a_27314_7850# a_27406_7484# 0.32fF
C3155 vcm_commonmode a_29322_9858# 0.31fF
C3156 m3_29316_72146# VDD 0.40fF
C3157 a_3983_65327# VDD 0.44fF
C3158 a_38450_24552# m3_38352_24414# 2.81fF
C3159 a_43470_63198# a_44474_63198# 0.97fF
C3160 vcm_commonmode a_45386_16886# 0.31fF
C3161 a_4960_40847# a_5098_41641# 0.77fF
C3162 a_15193_41781# a_15189_39889# 1.01fF
C3163 a_33338_72234# VDD 0.63fF
C3164 a_16928_42919# VDD 1.45fF
C3165 a_17366_18528# a_17366_17524# 1.00fF
C3166 a_10883_18543# VDD 0.40fF
C3167 a_30418_21540# a_31422_21540# 0.97fF
C3168 a_38358_9858# a_38450_9492# 0.32fF
C3169 a_4528_26159# VDD 2.17fF
C3170 a_21290_64202# a_21382_64202# 0.32fF
C3171 a_30418_7484# VDD 1.37fF
C3172 a_48490_58178# a_49494_58178# 0.97fF
C3173 a_1586_66567# a_5428_63669# 0.33fF
C3174 a_1950_59887# a_3024_67191# 0.55fF
C3175 vcm_commonmode a_37446_68218# 0.87fF
C3176 a_37446_59182# a_38450_59182# 0.97fF
C3177 a_18278_22910# a_18370_22544# 0.32fF
C3178 a_24394_64202# VDD 0.51fF
C3179 a_8123_56399# a_22989_48437# 0.30fF
C3180 a_1591_9839# a_1757_9839# 0.69fF
C3181 a_27752_7638# a_10515_23975# 0.41fF
C3182 a_32426_56170# ctopp 3.46fF
C3183 a_11521_66567# a_10515_63143# 0.36fF
C3184 a_18370_14512# a_18370_13508# 1.00fF
C3185 a_29035_38825# VDD 0.62fF
C3186 ctopn a_26402_18528# 3.59fF
C3187 a_5449_25071# a_4248_29967# 0.70fF
C3188 vcm_commonmode a_31330_64202# 0.31fF
C3189 a_35438_17524# a_36442_17524# 0.97fF
C3190 a_5915_35943# a_14646_29423# 0.31fF
C3191 a_22386_60186# a_23390_60186# 0.97fF
C3192 a_43175_28335# a_46482_21540# 0.38fF
C3193 a_39454_24552# a_39454_23548# 1.00fF
C3194 a_24394_12504# a_24394_11500# 1.00fF
C3195 a_41842_27221# VDD 1.65fF
C3196 a_1586_9991# a_1757_9839# 0.60fF
C3197 a_29760_7638# a_29414_11500# 0.38fF
C3198 a_17366_18528# a_18370_18528# 0.97fF
C3199 a_13123_38231# a_12473_36341# 0.35fF
C3200 a_2451_72373# a_1823_72381# 0.35fF
C3201 a_10575_62911# VDD 0.35fF
C3202 a_16863_29415# a_29175_28335# 0.77fF
C3203 a_31422_61190# ctopp 3.59fF
C3204 ctopn a_35438_10496# 3.59fF
C3205 a_33430_69222# VDD 0.51fF
C3206 a_20957_36604# VDD 0.88fF
C3207 vcm_commonmode a_19282_19898# 0.31fF
C3208 a_37527_29397# a_38436_29941# 0.30fF
C3209 a_2021_22325# a_12357_37999# 0.36fF
C3210 a_21371_50959# a_6831_63303# 1.19fF
C3211 a_14287_51175# a_18370_63198# 0.42fF
C3212 vcm_commonmode a_37446_56170# 0.87fF
C3213 a_34251_52263# a_12257_56623# 0.40fF
C3214 a_8289_14741# VDD 0.64fF
C3215 a_1761_8751# config_1_in[1] 0.31fF
C3216 a_34221_47695# VDD 0.34fF
C3217 vcm_commonmode a_40366_69222# 0.31fF
C3218 a_6559_59663# a_8199_58229# 0.72fF
C3219 a_46390_7850# a_46482_7484# 0.32fF
C3220 a_40458_22544# VDD 0.51fF
C3221 vcm_commonmode a_20378_8488# 0.86fF
C3222 a_31422_65206# VDD 0.51fF
C3223 ctopp a_32426_55166# 1.02fF
C3224 a_3339_43023# a_12869_2741# 0.86fF
C3225 a_7210_55081# a_8123_56399# 0.35fF
C3226 a_20027_27221# a_19889_27497# 0.42fF
C3227 a_21371_52263# a_6559_59663# 2.56fF
C3228 a_25971_52263# a_10515_22671# 0.40fF
C3229 a_7841_12167# VDD 9.25fF
C3230 vcm_commonmode a_47394_22910# 0.31fF
C3231 a_35438_70226# ctopp 3.58fF
C3232 a_35647_42405# VDD 0.85fF
C3233 vcm_commonmode a_38358_65206# 0.31fF
C3234 a_30326_69222# a_30418_69222# 0.32fF
C3235 a_36442_18528# a_36442_17524# 1.00fF
C3236 a_3339_43023# a_24029_39355# 0.39fF
C3237 a_19720_55394# a_21371_50959# 0.49fF
C3238 a_21382_72234# a_22386_72234# 0.97fF
C3239 a_14287_51175# a_21371_52263# 0.55fF
C3240 a_16955_52047# a_18151_52263# 0.89fF
C3241 a_8491_27023# a_12727_13353# 0.41fF
C3242 a_20286_24918# VDD 0.36fF
C3243 a_12355_15055# a_8295_47388# 0.41fF
C3244 a_40366_64202# a_40458_64202# 0.32fF
C3245 a_39331_34191# VDD 0.35fF
C3246 ctopn a_30418_15516# 3.59fF
C3247 a_29760_55394# a_28881_52271# 0.37fF
C3248 vcm_commonmode a_36442_61190# 0.87fF
C3249 a_5039_42167# a_3339_32463# 0.41fF
C3250 a_36442_14512# VDD 0.51fF
C3251 a_27752_7638# a_27406_10496# 0.38fF
C3252 a_10311_20175# VDD 0.33fF
C3253 a_31330_55166# VDD 0.35fF
C3254 a_39673_28111# a_12899_10927# 0.41fF
C3255 a_37354_22910# a_37446_22544# 0.32fF
C3256 a_2163_63293# VDD 0.49fF
C3257 a_26402_10496# a_27406_10496# 0.97fF
C3258 a_22562_28023# VDD 0.79fF
C3259 vcm_commonmode a_43378_14878# 0.31fF
C3260 ctopn a_40458_11500# 3.59fF
C3261 a_28318_65206# a_28410_65206# 0.32fF
C3262 a_37446_14512# a_37446_13508# 1.00fF
C3263 vcm_commonmode a_22294_20902# 0.31fF
C3264 a_28115_40183# VDD 0.62fF
C3265 a_16510_8760# a_2235_30503# 0.75fF
C3266 a_21187_29415# a_16863_29415# 0.37fF
C3267 a_14421_49007# VDD 0.54fF
C3268 vcm_commonmode a_40458_70226# 0.87fF
C3269 a_1586_51335# a_4891_47388# 2.22fF
C3270 a_41462_60186# a_42466_60186# 0.97fF
C3271 a_41462_23548# VDD 0.52fF
C3272 a_24394_58178# ctopp 3.59fF
C3273 a_19282_23914# a_19374_23548# 0.32fF
C3274 a_38450_66210# VDD 0.51fF
C3275 VDD dummypin[10] 0.94fF
C3276 a_43470_12504# a_43470_11500# 1.00fF
C3277 vcm_commonmode a_21382_16520# 0.87fF
C3278 a_14287_51175# a_12727_58255# 0.40fF
C3279 vcm_commonmode a_48398_23914# 0.31fF
C3280 a_1761_52815# a_3305_38671# 0.39fF
C3281 a_22671_43439# VDD 2.07fF
C3282 a_43267_31055# a_12983_63151# 0.40fF
C3283 a_30418_70226# a_30418_69222# 1.00fF
C3284 vcm_commonmode a_45386_66210# 0.31fF
C3285 a_36442_18528# a_37446_18528# 0.97fF
C3286 vcm_commonmode a_20378_72234# 0.69fF
C3287 a_32772_7638# a_32426_16520# 0.38fF
C3288 a_1803_19087# a_1849_31599# 0.35fF
C3289 vcm_commonmode a_22294_12870# 0.31fF
C3290 a_8491_27023# a_10515_23975# 0.41fF
C3291 a_16362_24552# a_17366_24552# 0.97fF
C3292 a_36579_35831# VDD 0.66fF
C3293 a_41462_67214# ctopp 3.59fF
C3294 a_30052_32117# a_9503_26151# 4.95fF
C3295 a_42985_46831# a_12981_62313# 0.40fF
C3296 a_11067_13095# a_1761_39215# 0.33fF
C3297 a_28318_19898# a_28410_19532# 0.32fF
C3298 a_32951_27247# a_33430_13508# 0.38fF
C3299 a_2021_22325# a_4351_26703# 0.81fF
C3300 a_3339_43023# a_2021_22325# 0.41fF
C3301 a_9135_27239# a_12985_19087# 0.41fF
C3302 a_21187_29415# a_23685_29111# 0.33fF
C3303 a_29414_11500# a_29414_10496# 1.00fF
C3304 vcm_commonmode a_29414_58178# 0.87fF
C3305 a_33338_14878# a_33430_14512# 0.32fF
C3306 vcm_commonmode a_17274_21906# 0.33fF
C3307 a_2787_30503# a_13143_29575# 0.51fF
C3308 a_49402_69222# a_49494_69222# 0.32fF
C3309 a_42718_27497# a_44474_9492# 0.38fF
C3310 a_14831_50095# a_17682_50095# 3.49fF
C3311 a_36717_47375# a_36442_72234# 0.35fF
C3312 a_27406_55166# a_28410_55166# 0.97fF
C3313 a_5531_22895# a_5839_22351# 0.62fF
C3314 a_28756_7638# a_28410_21540# 0.38fF
C3315 a_24716_31757# VDD 0.69fF
C3316 vcm_commonmode a_22294_17890# 0.31fF
C3317 a_11067_13095# a_8453_51727# 0.48fF
C3318 a_43269_29967# a_43175_28335# 3.06fF
C3319 a_13067_38517# a_19967_41781# 0.57fF
C3320 a_18370_57174# a_19374_57174# 0.97fF
C3321 a_21382_15516# a_22386_15516# 0.97fF
C3322 vcm_commonmode a_46482_67214# 0.87fF
C3323 a_25744_7638# a_25398_18528# 0.38fF
C3324 a_8491_27023# a_18370_18528# 0.38fF
C3325 a_42466_63198# VDD 0.57fF
C3326 a_12447_29199# a_16101_31029# 0.67fF
C3327 a_45478_10496# a_46482_10496# 0.97fF
C3328 a_47394_65206# a_47486_65206# 0.32fF
C3329 vcm_commonmode a_49402_63198# 0.30fF
C3330 a_19374_71230# a_20378_71230# 0.97fF
C3331 vcm_commonmode a_12901_66959# 6.23fF
C3332 a_36442_59182# VDD 0.51fF
C3333 a_11067_21583# VDD 9.09fF
C3334 vcm_commonmode a_43470_9492# 0.87fF
C3335 a_38358_23914# a_38450_23548# 0.32fF
C3336 a_31422_11500# a_32426_11500# 0.97fF
C3337 a_40458_64202# ctopp 3.59fF
C3338 ctopn a_45478_13508# 3.59fF
C3339 a_12899_3311# a_25744_7638# 1.78fF
C3340 a_1761_43567# a_1761_27791# 0.72fF
C3341 a_39299_48783# VDD 7.00fF
C3342 a_35346_66210# a_35438_66210# 0.32fF
C3343 vcm_commonmode a_43378_59182# 0.31fF
C3344 vcm_commonmode a_23390_22544# 0.87fF
C3345 a_40585_42369# VDD 1.87fF
C3346 a_34251_52263# a_10975_66407# 0.40fF
C3347 a_49494_70226# a_49494_69222# 1.00fF
C3348 a_16746_18526# VDD 33.20fF
C3349 a_17274_72234# a_17366_72234# 0.32fF
C3350 a_12546_22351# a_12985_19087# 24.16fF
C3351 a_13669_39605# a_1761_35407# 1.50fF
C3352 a_11067_67279# a_5039_42167# 0.81fF
C3353 a_35438_24552# a_36442_24552# 0.97fF
C3354 vcm_commonmode a_23298_18894# 0.31fF
C3355 a_16746_66212# ctopp 1.68fF
C3356 a_16863_29415# a_26523_28111# 1.91fF
C3357 a_20359_29199# a_8491_41383# 0.70fF
C3358 a_47394_19898# a_47486_19532# 0.32fF
C3359 a_11067_47695# a_22989_48437# 1.25fF
C3360 a_48490_21540# VDD 0.55fF
C3361 a_32426_62194# a_33430_62194# 0.97fF
C3362 a_48490_11500# a_48490_10496# 1.00fF
C3363 vcm_commonmode a_19374_14512# 0.87fF
C3364 ctopn a_16746_11498# 1.68fF
C3365 a_2191_68565# VDD 5.30fF
C3366 a_12355_65103# a_16362_64202# 1.15fF
C3367 a_42985_46831# a_48490_59182# 0.38fF
C3368 a_13909_37571# VDD 0.55fF
C3369 a_25398_10496# VDD 0.51fF
C3370 a_30035_40767# VDD 0.82fF
C3371 vcm_commonmode a_45478_64202# 0.87fF
C3372 a_7580_61751# a_7155_55509# 0.34fF
C3373 a_22843_29415# a_20635_29415# 1.05fF
C3374 a_18151_52263# a_24394_71230# 0.38fF
C3375 a_25971_52263# a_12901_66665# 0.40fF
C3376 vcm_commonmode a_16362_70226# 4.47fF
C3377 a_31330_20902# a_31422_20536# 0.32fF
C3378 a_40458_60186# VDD 0.51fF
C3379 a_45478_55166# a_46482_55166# 0.97fF
C3380 vcm_commonmode a_32334_10862# 0.31fF
C3381 vcm_commonmode a_76971_38925# 673.41fF
C3382 a_10501_65871# VDD 0.50fF
C3383 a_20635_29415# a_23395_32463# 0.40fF
C3384 a_20286_63198# a_20378_63198# 0.32fF
C3385 a_47486_65206# ctopp 3.58fF
C3386 a_37446_57174# a_38450_57174# 0.97fF
C3387 vcm_commonmode a_47394_60186# 0.31fF
C3388 a_34251_52263# a_35438_61190# 0.38fF
C3389 a_40458_15516# a_41462_15516# 0.97fF
C3390 vcm_commonmode a_24394_23548# 0.87fF
C3391 a_24800_44129# VDD 1.37fF
C3392 a_18611_52047# a_23390_67214# 0.38fF
C3393 vcm_commonmode a_21382_66210# 0.87fF
C3394 a_10687_52553# VDD 6.42fF
C3395 a_26748_7638# a_12985_16367# 0.41fF
C3396 a_13743_35836# VDD 1.14fF
C3397 vcm_commonmode a_33430_19532# 0.87fF
C3398 a_40458_58178# a_40458_59182# 1.00fF
C3399 a_12549_44212# a_13005_43983# 0.31fF
C3400 vcm_commonmode a_19282_62194# 0.31fF
C3401 a_20378_15516# VDD 0.51fF
C3402 a_1586_40455# a_1761_47919# 0.32fF
C3403 a_38450_71230# a_39454_71230# 0.97fF
C3404 a_16362_19532# a_12895_13967# 1.27fF
C3405 m3_16264_7346# VDD 0.38fF
C3406 a_2411_19605# a_3983_20719# 0.52fF
C3407 vcm_commonmode a_27314_15882# 0.31fF
C3408 a_20378_63198# ctopp 3.64fF
C3409 a_3143_22364# a_3972_25615# 0.53fF
C3410 a_18370_71230# VDD 0.58fF
C3411 a_21371_52263# a_12901_58799# 0.40fF
C3412 a_30418_11500# VDD 0.51fF
C3413 vcm_commonmode a_25306_71230# 0.31fF
C3414 a_27314_72234# a_27406_72234# 0.32fF
C3415 a_36629_27791# a_12727_15529# 0.41fF
C3416 a_34434_24552# VDD 0.60fF
C3417 vcm_commonmode a_37354_11866# 0.31fF
C3418 a_16746_67216# VDD 33.19fF
C3419 a_18370_64202# a_18370_63198# 1.23fF
C3420 a_31330_12870# a_31422_12504# 0.32fF
C3421 a_5993_32687# VDD 1.74fF
C3422 a_2099_59861# a_17711_32385# 0.34fF
C3423 a_8531_70543# a_12869_2741# 0.57fF
C3424 vcm_commonmode a_41370_24918# 0.31fF
C3425 a_19788_48981# a_20853_47375# 0.38fF
C3426 a_26402_59182# a_26402_58178# 1.00fF
C3427 a_44474_55166# VDD 0.60fF
C3428 a_20635_29415# a_41334_29575# 0.33fF
C3429 a_12447_29199# a_14926_31849# 0.44fF
C3430 a_1823_54973# a_1757_51183# 0.32fF
C3431 a_6066_28309# VDD 0.47fF
C3432 a_36442_57174# VDD 0.51fF
C3433 a_8491_27023# a_9669_26703# 0.50fF
C3434 a_28547_51175# a_32426_58178# 0.38fF
C3435 a_17366_13508# a_18370_13508# 0.97fF
C3436 vcm_commonmode a_36442_20536# 0.87fF
C3437 ctopn a_16362_17524# 1.35fF
C3438 a_4427_30511# a_4248_29967# 0.42fF
C3439 a_2927_39733# a_2021_17973# 0.70fF
C3440 a_13097_39631# VDD 1.26fF
C3441 a_22386_68218# a_23390_68218# 0.97fF
C3442 a_29760_55394# a_12355_15055# 0.40fF
C3443 vcm_commonmode a_25398_63198# 0.92fF
C3444 a_32951_27247# a_33430_7484# 0.34fF
C3445 vcm_commonmode a_43378_57174# 0.31fF
C3446 a_22259_48981# VDD 0.67fF
C3447 a_40458_72234# a_40458_71230# 1.00fF
C3448 a_7871_59049# VDD 0.58fF
C3449 a_12727_58255# a_12901_58799# 23.51fF
C3450 a_17488_48731# a_17711_32385# 0.63fF
C3451 a_34434_56170# a_34434_55166# 1.00fF
C3452 a_31422_24552# m3_31324_24414# 2.81fF
C3453 a_39362_63198# a_39454_63198# 0.32fF
C3454 a_16362_64202# ctopp 1.35fF
C3455 a_17507_52047# a_20359_29199# 0.68fF
C3456 a_44474_58178# ctopp 3.59fF
C3457 a_30418_57174# a_30418_56170# 1.00fF
C3458 a_26310_72234# VDD 0.62fF
C3459 vcm_commonmode a_19374_59182# 0.87fF
C3460 VDD result_out[7] 0.66fF
C3461 a_3339_43023# m2_48260_24282# 0.37fF
C3462 a_12641_43124# VDD 2.59fF
C3463 a_5924_69135# a_4307_67477# 0.79fF
C3464 a_6271_72943# a_5023_72068# 0.34fF
C3465 a_26310_21906# a_26402_21540# 0.32fF
C3466 a_22291_29415# a_31768_7638# 0.75fF
C3467 vcm_commonmode a_36442_12504# 0.87fF
C3468 a_18370_60186# ctopp 3.58fF
C3469 ctopn a_37446_9492# 3.58fF
C3470 a_21382_68218# VDD 0.51fF
C3471 a_16746_64204# a_16362_64202# 2.28fF
C3472 a_24800_35425# VDD 1.71fF
C3473 a_2840_53511# a_6835_46823# 0.91fF
C3474 a_1591_43029# a_1757_43029# 0.44fF
C3475 a_21290_7850# VDD 0.63fF
C3476 a_44382_58178# a_44474_58178# 0.32fF
C3477 a_42985_46831# a_48490_57174# 0.38fF
C3478 ctopn a_17366_22544# 3.24fF
C3479 a_7939_30503# a_14646_29423# 1.68fF
C3480 a_1761_49007# a_1761_47919# 1.32fF
C3481 a_5831_39189# VDD 10.85fF
C3482 vcm_commonmode a_28318_68218# 0.31fF
C3483 a_33338_59182# a_33430_59182# 0.32fF
C3484 a_32951_27247# a_12985_19087# 0.41fF
C3485 a_17712_7638# a_12895_13967# 0.40fF
C3486 a_22843_29415# a_26694_29473# 0.40fF
C3487 a_15305_38543# VDD 2.02fF
C3488 vcm_commonmode a_31422_21540# 0.87fF
C3489 a_3983_45743# a_4149_45743# 0.72fF
C3490 a_30875_41271# VDD 0.63fF
C3491 a_31330_17890# a_31422_17524# 0.32fF
C3492 vcm_commonmode a_49494_58178# 0.91fF
C3493 a_12473_36341# a_31131_35281# 0.31fF
C3494 a_1761_50639# a_1761_49007# 3.61fF
C3495 a_16362_60186# VDD 2.48fF
C3496 a_18278_60186# a_18370_60186# 0.32fF
C3497 a_37446_64202# a_37446_63198# 1.23fF
C3498 vcm_commonmode a_36442_17524# 0.87fF
C3499 a_12725_44527# a_27263_40871# 0.64fF
C3500 a_6435_74005# VDD 0.36fF
C3501 vcm_commonmode a_23390_60186# 0.87fF
C3502 a_35438_13508# VDD 0.51fF
C3503 a_12907_27023# a_20267_30503# 0.97fF
C3504 a_40458_58178# a_40458_57174# 1.00fF
C3505 a_7794_53903# VDD 0.34fF
C3506 a_29414_22544# a_29414_21540# 1.00fF
C3507 a_8935_27791# VDD 1.25fF
C3508 a_21382_56170# VDD 0.52fF
C3509 a_1768_16367# config_2_in[10] 0.63fF
C3510 vcm_commonmode a_42374_13874# 0.31fF
C3511 a_8491_27023# a_9263_24501# 1.72fF
C3512 a_36442_13508# a_37446_13508# 0.97fF
C3513 a_32121_44545# a_13716_43047# 0.53fF
C3514 a_4211_67655# a_3668_56311# 0.48fF
C3515 a_41462_68218# a_42466_68218# 0.97fF
C3516 vcm_commonmode a_28318_56170# 0.31fF
C3517 a_28756_55394# a_12257_56623# 0.40fF
C3518 ctopn a_18370_23548# 3.28fF
C3519 a_43175_28335# a_12985_19087# 0.41fF
C3520 a_6607_42167# a_6372_38279# 0.88fF
C3521 a_22386_56170# a_23390_56170# 0.97fF
C3522 a_49494_57174# a_49494_56170# 1.00fF
C3523 a_18611_52047# a_10515_22671# 0.45fF
C3524 a_7917_13885# a_3327_9308# 0.40fF
C3525 ctopn a_27406_19532# 3.59fF
C3526 a_3983_10927# VDD 0.39fF
C3527 a_15775_42405# VDD 0.96fF
C3528 a_42709_29199# a_48490_8488# 0.38fF
C3529 a_25939_51157# VDD 0.53fF
C3530 a_8575_74853# a_9063_71553# 0.34fF
C3531 a_45386_21906# a_45478_21540# 0.32fF
C3532 a_20378_61190# VDD 0.51fF
C3533 a_4333_22895# VDD 0.91fF
C3534 a_26402_58178# a_26402_57174# 1.00fF
C3535 a_24740_7638# a_11067_21583# 0.41fF
C3536 a_11943_63125# a_11067_63143# 1.03fF
C3537 a_27560_34337# VDD 1.14fF
C3538 vcm_commonmode a_37446_18528# 0.87fF
C3539 a_22671_43439# a_12663_40871# 0.42fF
C3540 a_1761_43567# a_1761_41935# 1.23fF
C3541 vcm_commonmode a_27314_61190# 0.31fF
C3542 a_33430_16520# a_33430_15516# 1.00fF
C3543 vcm_commonmode a_17366_24552# 0.84fF
C3544 a_1689_10396# a_2283_15797# 0.84fF
C3545 a_18370_19532# a_18370_18528# 1.00fF
C3546 a_1867_20175# VDD 0.42fF
C3547 a_43269_29967# a_12985_16367# 0.41fF
C3548 a_22294_10862# a_22386_10496# 0.32fF
C3549 a_28410_62194# ctopp 3.59fF
C3550 a_24394_70226# VDD 0.51fF
C3551 a_41351_38053# VDD 1.19fF
C3552 a_41462_58178# VDD 0.51fF
C3553 vcm_commonmode a_28410_55166# 0.84fF
C3554 a_32367_28309# a_12899_3855# 0.54fF
C3555 vcm_commonmode a_19374_57174# 0.87fF
C3556 a_10239_16367# VDD 0.46fF
C3557 vcm_commonmode a_31330_70226# 0.31fF
C3558 a_2843_71829# a_5213_70223# 0.46fF
C3559 a_37354_60186# a_37446_60186# 0.32fF
C3560 vcm_commonmode a_46482_10496# 0.87fF
C3561 a_16863_29415# a_35815_31751# 0.62fF
C3562 a_13183_52047# VDD 11.11fF
C3563 a_34434_71230# ctopp 3.40fF
C3564 a_2004_42453# a_2283_15797# 1.03fF
C3565 ctopn a_30418_20536# 3.59fF
C3566 a_11416_12283# VDD 0.51fF
C3567 a_39389_52271# a_12983_63151# 0.40fF
C3568 a_43269_29967# a_47486_8488# 0.38fF
C3569 a_32334_18894# a_32426_18528# 0.32fF
C3570 a_1761_37039# a_1761_30511# 0.35fF
C3571 a_48490_22544# a_48490_21540# 1.00fF
C3572 a_11067_46823# a_27250_27791# 0.50fF
C3573 a_21382_61190# a_22386_61190# 0.97fF
C3574 a_9135_27239# VDD 10.58fF
C3575 a_1586_18695# config_1_in[12] 0.39fF
C3576 a_39223_32463# a_39454_19532# 0.38fF
C3577 a_2927_68565# VDD 1.77fF
C3578 a_19594_35823# VDD 1.25fF
C3579 a_42466_8488# VDD 0.58fF
C3580 a_41427_52263# a_12981_62313# 0.40fF
C3581 a_27406_68218# a_27406_67214# 1.00fF
C3582 vcm_commonmode a_33430_62194# 0.87fF
C3583 a_7571_29199# VDD 10.39fF
C3584 a_2099_59861# a_7295_44647# 2.40fF
C3585 a_12263_20969# VDD 0.56fF
C3586 vcm_commonmode a_49402_8854# 0.30fF
C3587 a_43270_27791# a_12985_19087# 0.41fF
C3588 vcm_commonmode a_41462_15516# 0.87fF
C3589 ctopn a_30418_12504# 3.59fF
C3590 a_11866_27791# a_9135_27239# 0.43fF
C3591 a_41462_56170# a_42466_56170# 0.97fF
C3592 vcm_commonmode a_20286_58178# 0.31fF
C3593 a_35647_39141# VDD 0.87fF
C3594 a_36797_27497# a_37446_9492# 0.38fF
C3595 a_3339_43023# ctopn 0.43fF
C3596 a_1761_30511# a_1761_32143# 1.02fF
C3597 vcm_commonmode a_39454_71230# 0.86fF
C3598 a_19720_7638# a_19374_15516# 0.38fF
C3599 a_23298_55166# a_23390_55166# 0.32fF
C3600 a_24394_8488# a_25398_8488# 0.97fF
C3601 a_30418_67214# VDD 0.51fF
C3602 a_12631_28585# a_15661_29199# 0.34fF
C3603 a_11803_55311# a_4758_45369# 0.32fF
C3604 a_4351_67279# a_11145_60431# 0.43fF
C3605 a_17274_15882# a_17366_15516# 0.32fF
C3606 ctopn a_25398_21540# 3.59fF
C3607 a_7695_31573# a_11143_31599# 0.35fF
C3608 a_1895_12730# VDD 0.51fF
C3609 a_41872_29423# a_12727_67753# 0.40fF
C3610 vcm_commonmode a_37354_67214# 0.31fF
C3611 a_25398_70226# a_26402_70226# 0.97fF
C3612 a_37446_19532# a_37446_18528# 1.00fF
C3613 a_41370_10862# a_41462_10496# 0.32fF
C3614 vcm_commonmode a_18370_13508# 0.88fF
C3615 a_1757_69141# VDD 0.66fF
C3616 a_37446_68218# ctopp 3.59fF
C3617 ctopn a_30418_17524# 3.59fF
C3618 a_1761_25071# a_1761_43567# 1.10fF
C3619 a_27406_9492# VDD 0.51fF
C3620 a_36671_39913# VDD 0.63fF
C3621 a_43470_16520# VDD 0.51fF
C3622 a_23390_60186# a_23390_59182# 1.00fF
C3623 a_1591_38677# a_1757_38677# 0.47fF
C3624 a_12546_22351# VDD 11.16fF
C3625 vcm_commonmode a_34342_9858# 0.31fF
C3626 a_27314_11866# a_27406_11500# 0.32fF
C3627 a_32823_29397# VDD 4.21fF
C3628 a_25787_28327# a_21187_29415# 0.50fF
C3629 a_12473_41781# a_19967_41781# 2.66fF
C3630 a_36613_48169# VDD 7.05fF
C3631 a_32426_15516# a_32426_14512# 1.00fF
C3632 vcm_commonmode m3_16264_64114# 3.25fF
C3633 a_28756_55394# a_10975_66407# 0.40fF
C3634 a_29760_7638# a_29414_10496# 0.38fF
C3635 a_16152_37601# a_1761_35407# 3.47fF
C3636 a_1757_51183# VDD 0.44fF
C3637 vcm_commonmode a_41261_28335# 10.07fF
C3638 a_2497_61519# VDD 0.48fF
C3639 a_7571_29199# a_18053_28879# 0.55fF
C3640 a_40458_61190# a_41462_61190# 0.97fF
C3641 a_17366_9492# a_17366_8488# 1.00fF
C3642 a_31330_24918# a_31422_24552# 0.32fF
C3643 a_21187_29415# a_2235_30503# 0.58fF
C3644 a_15345_34717# VDD 0.97fF
C3645 a_32038_29575# a_33008_28853# 0.35fF
C3646 a_35438_7484# VDD 1.23fF
C3647 a_11521_66567# a_11659_66567# 0.65fF
C3648 a_46482_68218# a_46482_67214# 1.00fF
C3649 a_1591_59343# result_out[5] 0.51fF
C3650 a_4681_13621# VDD 0.57fF
C3651 vcm_commonmode a_42466_68218# 0.87fF
C3652 a_40050_48463# a_12901_66959# 0.40fF
C3653 a_26748_7638# a_26402_18528# 0.38fF
C3654 a_29414_64202# VDD 0.51fF
C3655 a_28318_62194# a_28410_62194# 0.32fF
C3656 a_37446_56170# ctopp 3.40fF
C3657 a_39299_48783# a_44474_59182# 0.38fF
C3658 ctopn a_31422_18528# 3.59fF
C3659 vcm_commonmode a_36350_64202# 0.31fF
C3660 a_31422_69222# a_31422_68218# 1.00fF
C3661 a_18611_52047# a_12901_66665# 0.40fF
C3662 a_46482_72234# a_47486_72234# 0.97fF
C3663 a_16955_52047# a_20378_71230# 0.38fF
C3664 a_43267_31055# a_42985_46831# 0.40fF
C3665 a_41370_55166# a_41462_55166# 0.32fF
C3666 a_11130_22869# VDD 0.97fF
C3667 a_43470_8488# a_44474_8488# 0.97fF
C3668 a_21382_8488# a_21382_7484# 1.00fF
C3669 a_4339_64521# a_10472_52423# 0.31fF
C3670 a_12357_37999# a_13837_38772# 0.30fF
C3671 a_5767_31573# VDD 0.41fF
C3672 a_33338_57174# a_33430_57174# 0.32fF
C3673 a_1950_59887# a_6737_60431# 0.41fF
C3674 a_31768_55394# a_31422_61190# 0.38fF
C3675 a_36350_15882# a_36442_15516# 0.32fF
C3676 a_19720_55394# a_19374_67214# 0.38fF
C3677 a_44474_70226# a_45478_70226# 0.97fF
C3678 a_32951_27247# a_33430_11500# 0.38fF
C3679 a_17366_19532# VDD 0.57fF
C3680 a_36442_61190# ctopp 3.59fF
C3681 ctopn a_40458_10496# 3.59fF
C3682 a_38450_69222# VDD 0.51fF
C3683 vcm_commonmode a_24302_19898# 0.31fF
C3684 a_40050_48463# a_45478_64202# 0.38fF
C3685 a_25398_16520# a_26402_16520# 0.97fF
C3686 vcm_commonmode a_42466_56170# 0.87fF
C3687 a_2873_13879# VDD 1.02fF
C3688 a_4427_25071# start_conversion_in 0.45fF
C3689 a_34342_71230# a_34434_71230# 0.32fF
C3690 vcm_commonmode a_45386_69222# 0.31fF
C3691 a_1923_54591# VDD 5.01fF
C3692 a_40458_58178# a_39222_48169# 0.38fF
C3693 a_1823_58773# a_2695_58951# 0.43fF
C3694 a_42466_60186# a_42466_59182# 1.00fF
C3695 a_38315_39141# a_38101_38565# 0.32fF
C3696 a_45478_22544# VDD 0.51fF
C3697 vcm_commonmode a_25398_8488# 0.86fF
C3698 m3_16264_21402# VDD 0.34fF
C3699 a_36442_65206# VDD 0.51fF
C3700 a_31422_63198# a_31422_62194# 1.00fF
C3701 a_46390_11866# a_46482_11500# 0.32fF
C3702 a_28670_30663# VDD 0.91fF
C3703 a_19720_55394# a_12901_58799# 0.40fF
C3704 a_40458_70226# ctopp 3.58fF
C3705 vcm_commonmode m3_16264_11362# 3.21fF
C3706 a_17366_72234# m3_17268_72146# 2.80fF
C3707 a_1761_49007# a_12889_40977# 0.32fF
C3708 a_7295_44647# a_1761_25071# 0.57fF
C3709 a_15459_41781# VDD 2.94fF
C3710 vcm_commonmode a_43378_65206# 0.31fF
C3711 a_40675_27791# a_41462_9492# 0.38fF
C3712 a_17712_7638# a_17366_9492# 0.38fF
C3713 a_17039_51157# a_11067_46823# 1.59fF
C3714 vcm_commonmode a_16746_71232# 5.34fF
C3715 a_12447_29199# a_31117_28879# 0.30fF
C3716 a_36442_9492# a_36442_8488# 1.00fF
C3717 a_25306_24918# VDD 0.36fF
C3718 a_1823_66941# VDD 3.26fF
C3719 ctopn a_35438_15516# 3.59fF
C3720 a_28547_51175# a_38115_52263# 0.67fF
C3721 vcm_commonmode a_41462_61190# 0.87fF
C3722 a_31422_67214# a_32426_67214# 0.97fF
C3723 a_2292_43291# a_7407_46529# 0.34fF
C3724 a_41462_14512# VDD 0.51fF
C3725 a_1895_18756# a_1757_18543# 0.70fF
C3726 a_10687_52553# a_19502_51157# 0.32fF
C3727 a_20378_20536# VDD 0.51fF
C3728 a_35346_55166# VDD 0.35fF
C3729 a_6831_63303# a_26662_48981# 0.56fF
C3730 a_12341_3311# a_12985_19087# 0.41fF
C3731 a_3305_38671# a_5691_36727# 0.36fF
C3732 a_6372_38279# a_6883_37019# 0.64fF
C3733 a_47394_62194# a_47486_62194# 0.32fF
C3734 vcm_commonmode a_48398_14878# 0.31fF
C3735 ctopn a_45478_11500# 3.59fF
C3736 a_28756_55394# a_28410_58178# 0.38fF
C3737 a_14859_37737# VDD 0.56fF
C3738 vcm_commonmode a_27314_20902# 0.31fF
C3739 a_49876_37608# VDD 0.97fF
C3740 vcm_commonmode a_15439_49525# 4.81fF
C3741 a_18278_68218# a_18370_68218# 0.32fF
C3742 a_17599_52263# a_12355_15055# 0.40fF
C3743 a_42985_46831# a_48490_65206# 0.38fF
C3744 a_11067_13095# a_5631_38127# 0.32fF
C3745 a_11297_49257# VDD 0.66fF
C3746 vcm_commonmode a_45478_70226# 0.87fF
C3747 a_36442_72234# a_36442_71230# 1.00fF
C3748 a_46482_23548# VDD 0.52fF
C3749 a_17366_7484# a_18370_7484# 0.97fF
C3750 a_40458_8488# a_40458_7484# 1.00fF
C3751 a_29414_58178# ctopp 3.59fF
C3752 a_43470_66210# VDD 0.51fF
C3753 VDD dummypin[14] 0.95fF
C3754 a_24394_24552# m3_24296_24414# 2.81fF
C3755 a_5254_67503# a_8491_57487# 0.52fF
C3756 a_14679_31288# VDD 0.52fF
C3757 vcm_commonmode a_26402_16520# 0.87fF
C3758 a_34251_52263# a_27535_30503# 5.66fF
C3759 a_19282_72234# VDD 0.61fF
C3760 a_11803_55311# a_12981_59343# 1.07fF
C3761 a_20378_12504# VDD 0.51fF
C3762 a_3339_43023# a_12801_38517# 1.40fF
C3763 a_33430_58178# a_34434_58178# 0.97fF
C3764 a_27752_7638# a_27406_15516# 0.38fF
C3765 a_28410_9492# a_29414_9492# 0.97fF
C3766 a_32951_27247# VDD 6.31fF
C3767 vcm_commonmode a_27314_12870# 0.31fF
C3768 a_29414_13508# a_29414_12504# 1.00fF
C3769 a_46482_67214# ctopp 3.59fF
C3770 a_1689_10396# a_4446_40553# 0.57fF
C3771 a_44474_16520# a_45478_16520# 0.97fF
C3772 a_39299_48783# a_44474_57174# 0.38fF
C3773 a_2235_30503# a_2787_30503# 1.08fF
C3774 a_20635_29415# a_38067_47349# 0.50fF
C3775 a_3247_20495# a_4528_26159# 0.70fF
C3776 vcm_commonmode a_18370_7484# 0.69fF
C3777 a_1823_63677# VDD 2.02fF
C3778 a_2315_24540# a_2899_27023# 0.35fF
C3779 a_30023_41959# a_26550_40871# 0.50fF
C3780 vcm_commonmode a_34434_58178# 0.87fF
C3781 a_76346_38962# VDD 0.72fF
C3782 vcm_commonmode a_22294_21906# 0.31fF
C3783 a_12901_66959# ctopp 3.23fF
C3784 a_16707_41271# VDD 0.62fF
C3785 a_20378_17524# VDD 0.51fF
C3786 a_26155_50095# a_26321_50095# 0.69fF
C3787 a_19531_49007# VDD 0.59fF
C3788 a_29760_7638# a_12727_15529# 0.41fF
C3789 vcm_commonmode a_27314_17890# 0.31fF
C3790 a_11067_13095# a_4351_26703# 0.40fF
C3791 a_19374_67214# a_19374_66210# 1.00fF
C3792 a_23395_32463# a_41842_27221# 2.31fF
C3793 a_21479_44581# VDD 0.83fF
C3794 a_3228_54171# VDD 0.69fF
C3795 a_47486_63198# VDD 0.57fF
C3796 a_13669_39605# a_27652_38237# 0.59fF
C3797 a_43175_28335# VDD 6.32fF
C3798 ctopn a_16746_10494# 1.68fF
C3799 a_9955_20969# a_9751_25071# 0.94fF
C3800 a_32334_13874# a_32426_13508# 0.32fF
C3801 a_29943_36965# VDD 0.96fF
C3802 a_2021_22325# a_1803_20719# 5.14fF
C3803 a_1768_13103# rst_n 0.41fF
C3804 a_7580_61751# a_7833_66415# 0.31fF
C3805 a_1586_66567# a_7000_65595# 0.60fF
C3806 a_37354_68218# a_37446_68218# 0.32fF
C3807 a_17507_52047# a_12257_56623# 0.40fF
C3808 vcm_commonmode a_21382_69222# 0.87fF
C3809 a_41462_59182# VDD 0.51fF
C3810 a_36442_7484# a_37446_7484# 0.97fF
C3811 vcm_commonmode a_48490_9492# 0.87fF
C3812 VDD dummypin[5] 0.94fF
C3813 a_12786_30761# VDD 0.55fF
C3814 a_45478_64202# ctopp 3.59fF
C3815 a_18278_56170# a_18370_56170# 0.32fF
C3816 vcm_commonmode a_48398_59182# 0.31fF
C3817 vcm_commonmode a_28410_22544# 0.87fF
C3818 a_11067_67279# a_31768_7638# 0.41fF
C3819 a_16362_70226# ctopp 1.35fF
C3820 a_7295_44647# a_2787_32679# 0.76fF
C3821 vcm_commonmode a_19374_65206# 0.87fF
C3822 a_20378_69222# a_21382_69222# 0.97fF
C3823 a_21382_18528# VDD 0.51fF
C3824 a_47486_9492# a_48490_9492# 0.97fF
C3825 a_7519_59575# a_7749_55535# 0.82fF
C3826 ctopn a_19374_8488# 3.40fF
C3827 a_24740_7638# a_12546_22351# 0.41fF
C3828 a_4443_46607# a_13097_36367# 0.39fF
C3829 a_30418_64202# a_31422_64202# 0.97fF
C3830 a_48490_13508# a_48490_12504# 1.00fF
C3831 a_8570_34319# VDD 0.40fF
C3832 vcm_commonmode a_28318_18894# 0.31fF
C3833 a_21382_66210# ctopp 3.59fF
C3834 a_7695_31573# a_9367_29397# 0.81fF
C3835 a_11067_46823# a_20853_47375# 0.41fF
C3836 a_6831_63303# a_27869_50095# 1.60fF
C3837 a_27406_22544# a_28410_22544# 0.97fF
C3838 a_12447_29199# a_30788_28487# 0.32fF
C3839 a_3016_60949# a_2775_46025# 0.40fF
C3840 a_4771_56597# VDD 0.36fF
C3841 vcm_commonmode a_24394_14512# 0.87fF
C3842 a_18370_65206# a_19374_65206# 0.97fF
C3843 a_11067_67279# a_30764_7638# 0.41fF
C3844 vcm_commonmode a_19282_55166# 0.30fF
C3845 a_41842_27221# a_41334_29575# 0.48fF
C3846 a_4191_33449# a_4685_37583# 0.45fF
C3847 a_30418_10496# VDD 0.51fF
C3848 a_75475_40594# VDD 0.82fF
C3849 a_2689_65103# a_2840_66103# 0.48fF
C3850 a_6559_49557# a_6725_49557# 0.61fF
C3851 a_45478_60186# VDD 0.51fF
C3852 vcm_commonmode a_37354_10862# 0.31fF
C3853 a_18370_56170# a_18370_55166# 1.00fF
C3854 a_19004_40413# a_12473_41781# 1.93fF
C3855 a_7803_55509# a_2840_66103# 0.45fF
C3856 a_38450_67214# a_38450_66210# 1.00fF
C3857 a_12727_15529# a_16746_14510# 2.28fF
C3858 vcm_commonmode a_29414_23548# 0.87fF
C3859 a_4811_34855# a_23195_29967# 0.62fF
C3860 vcm_commonmode a_26402_66210# 0.87fF
C3861 a_28547_51175# a_12983_63151# 0.40fF
C3862 a_2143_15271# a_3983_16617# 0.68fF
C3863 a_1586_18695# a_10405_16367# 0.60fF
C3864 a_4831_52413# VDD 0.43fF
C3865 a_4758_45369# a_2292_43291# 1.11fF
C3866 a_17366_62194# VDD 0.57fF
C3867 a_12641_37684# a_25517_37455# 0.43fF
C3868 a_17274_61190# a_17366_61190# 0.32fF
C3869 a_43270_27791# VDD 6.68fF
C3870 a_34434_65206# a_34434_64202# 1.00fF
C3871 vcm_commonmode a_38450_19532# 0.87fF
C3872 ctopn a_20378_16520# 3.59fF
C3873 a_32823_29397# a_36904_28879# 0.62fF
C3874 vcm_commonmode a_24302_62194# 0.31fF
C3875 a_34780_56398# a_12981_62313# 0.40fF
C3876 a_25398_15516# VDD 0.51fF
C3877 a_18370_19532# a_19374_19532# 0.97fF
C3878 a_28410_23548# a_28410_22544# 1.00fF
C3879 a_6649_25615# VDD 1.91fF
C3880 vcm_commonmode a_32334_15882# 0.31fF
C3881 a_25398_63198# ctopp 3.64fF
C3882 a_37354_56170# a_37446_56170# 0.32fF
C3883 a_23390_71230# VDD 0.58fF
C3884 a_22386_66210# a_22386_65206# 1.00fF
C3885 a_23390_14512# a_24394_14512# 0.97fF
C3886 a_16615_39095# VDD 0.65fF
C3887 a_35438_11500# VDD 0.51fF
C3888 a_22595_42089# VDD 0.62fF
C3889 a_39454_69222# a_40458_69222# 0.97fF
C3890 a_22989_48437# a_23631_50069# 0.66fF
C3891 a_29760_55394# a_29414_72234# 0.34fF
C3892 vcm_commonmode a_30326_71230# 0.31fF
C3893 a_49402_61190# VDD 0.31fF
C3894 a_34434_61190# a_34434_60186# 1.00fF
C3895 a_20286_8854# a_20378_8488# 0.32fF
C3896 a_39454_24552# VDD 0.60fF
C3897 vcm_commonmode a_42374_11866# 0.31fF
C3898 a_19374_59182# ctopp 3.59fF
C3899 a_7571_26151# a_7598_36103# 0.36fF
C3900 a_4702_32143# VDD 0.52fF
C3901 a_2099_59861# a_9765_32143# 1.15fF
C3902 vcm_commonmode a_46390_24918# 0.31fF
C3903 ctopn a_16362_21540# 1.35fF
C3904 a_22015_28111# a_12447_29199# 0.81fF
C3905 a_21290_70226# a_21382_70226# 0.32fF
C3906 a_36717_47375# a_12727_67753# 0.40fF
C3907 a_5915_35943# a_5915_30287# 2.02fF
C3908 a_38358_58178# a_38450_58178# 0.32fF
C3909 a_46482_22544# a_47486_22544# 0.97fF
C3910 a_28756_7638# a_12877_16911# 0.41fF
C3911 a_20378_62194# a_20378_61190# 1.00fF
C3912 a_41462_57174# VDD 0.51fF
C3913 a_37446_65206# a_38450_65206# 0.97fF
C3914 a_7580_61751# a_6559_59879# 1.22fF
C3915 a_38499_37503# VDD 0.99fF
C3916 vcm_commonmode a_41462_20536# 0.87fF
C3917 a_32823_29397# a_38436_29941# 0.30fF
C3918 vcm_commonmode a_30418_63198# 0.92fF
C3919 a_10055_58791# ctopn 3.23fF
C3920 a_33430_17524# a_33430_16520# 1.00fF
C3921 a_18611_52047# a_9529_28335# 0.36fF
C3922 vcm_commonmode a_48398_57174# 0.31fF
C3923 a_23487_49007# VDD 0.50fF
C3924 a_20378_20536# a_20378_19532# 1.00fF
C3925 m3_16264_72146# VDD 0.38fF
C3926 a_19720_7638# a_19374_20536# 0.38fF
C3927 a_28410_23548# a_29414_23548# 0.97fF
C3928 a_4351_67279# a_28881_52271# 0.35fF
C3929 a_22671_43439# a_27263_40871# 0.40fF
C3930 a_25971_52263# VDD 17.35fF
C3931 vcm_commonmode a_24394_59182# 0.87fF
C3932 a_25398_66210# a_26402_66210# 0.97fF
C3933 a_17507_52047# a_10975_66407# 0.40fF
C3934 a_4495_35925# a_1761_30511# 0.52fF
C3935 vcm_commonmode a_34251_52263# 10.02fF
C3936 a_43175_28335# a_46482_16520# 0.38fF
C3937 a_36350_61190# a_36442_61190# 0.32fF
C3938 a_4758_45369# a_5190_59575# 1.04fF
C3939 a_1757_26159# VDD 0.31fF
C3940 vcm_commonmode a_41462_12504# 0.87fF
C3941 a_23390_60186# ctopp 3.59fF
C3942 ctopn a_42466_9492# 3.58fF
C3943 a_26402_68218# VDD 0.51fF
C3944 a_32143_35281# VDD 1.59fF
C3945 a_26310_7850# VDD 0.62fF
C3946 a_19410_43439# a_22671_43439# 1.17fF
C3947 ctopn a_22386_22544# 3.58fF
C3948 a_49494_10496# m3_49396_10358# 2.78fF
C3949 a_7862_34025# a_13357_32143# 0.31fF
C3950 a_25398_71230# a_25398_70226# 1.00fF
C3951 vcm_commonmode a_33338_68218# 0.31fF
C3952 a_38557_32143# a_12901_66959# 0.40fF
C3953 a_19720_7638# a_19374_12504# 0.38fF
C3954 a_37446_19532# a_38450_19532# 0.97fF
C3955 a_47486_23548# a_47486_22544# 1.00fF
C3956 a_9955_21807# a_11067_21583# 0.50fF
C3957 a_49876_37608# a_50198_39208# 0.73fF
C3958 a_14273_27791# a_12341_3311# 0.81fF
C3959 a_5682_69367# VDD 7.15fF
C3960 a_41462_66210# a_41462_65206# 1.00fF
C3961 a_39222_48169# a_40458_59182# 0.38fF
C3962 a_42466_14512# a_43470_14512# 0.97fF
C3963 a_24331_38591# VDD 1.01fF
C3964 vcm_commonmode a_36442_21540# 0.87fF
C3965 a_33641_29967# a_31084_30485# 0.72fF
C3966 a_2952_46805# a_1761_22895# 0.32fF
C3967 a_1757_40303# VDD 0.66fF
C3968 a_43270_27791# a_45478_8488# 0.38fF
C3969 a_6863_49722# a_6559_49557# 0.30fF
C3970 a_41872_29423# a_39299_48783# 1.67fF
C3971 a_21382_20536# a_22386_20536# 0.97fF
C3972 a_39362_8854# a_39454_8488# 0.32fF
C3973 a_1689_10396# a_4123_37013# 0.44fF
C3974 vcm_commonmode a_41462_17524# 0.87fF
C3975 ctopn a_18370_14512# 3.58fF
C3976 a_15661_29199# a_20027_27221# 0.83fF
C3977 a_11311_74005# VDD 0.47fF
C3978 a_23395_52047# a_27406_61190# 0.38fF
C3979 vcm_commonmode a_28410_60186# 0.87fF
C3980 a_40458_13508# VDD 0.51fF
C3981 a_39742_44527# VDD 0.47fF
C3982 a_40366_70226# a_40458_70226# 0.32fF
C3983 a_12516_7093# a_16362_69222# 1.15fF
C3984 a_13123_38231# a_1761_30511# 0.84fF
C3985 a_3063_19087# VDD 0.60fF
C3986 a_19720_7638# a_19374_17524# 0.38fF
C3987 a_4792_20443# a_7377_18012# 1.72fF
C3988 a_39454_62194# a_39454_61190# 1.00fF
C3989 a_30418_10496# a_30418_9492# 1.00fF
C3990 a_26402_56170# VDD 0.52fF
C3991 vcm_commonmode a_47394_13874# 0.31fF
C3992 a_1586_66567# a_6095_44807# 0.39fF
C3993 a_41427_52263# a_41462_64202# 0.38fF
C3994 a_21290_16886# a_21382_16520# 0.32fF
C3995 vcm_commonmode a_33338_56170# 0.31fF
C3996 ctopn a_23390_23548# 3.40fF
C3997 a_39454_20536# a_39454_19532# 1.00fF
C3998 a_11067_47695# a_2411_18517# 0.64fF
C3999 a_47486_23548# a_48490_23548# 0.97fF
C4000 a_20635_29415# a_29667_31055# 0.38fF
C4001 a_18979_30287# a_7862_34025# 0.76fF
C4002 a_7571_29199# a_9307_30663# 0.44fF
C4003 a_19374_57174# ctopp 3.58fF
C4004 a_11521_66567# a_11943_63125# 0.74fF
C4005 a_2840_66103# a_9735_63669# 0.30fF
C4006 a_44474_66210# a_45478_66210# 0.97fF
C4007 ctopn a_32426_19532# 3.59fF
C4008 a_41261_28335# a_12355_65103# 0.40fF
C4009 a_36629_27791# a_36442_9492# 0.38fF
C4010 a_1923_73087# a_1591_71317# 0.34fF
C4011 a_20286_72234# a_20378_72234# 0.32fF
C4012 a_19374_21540# a_19374_20536# 1.00fF
C4013 a_25398_61190# VDD 0.51fF
C4014 a_3987_19623# a_1586_21959# 0.76fF
C4015 a_12341_3311# VDD 12.87fF
C4016 vcm_commonmode a_18370_11500# 0.88fF
C4017 a_21382_12504# a_22386_12504# 0.97fF
C4018 a_35602_34191# VDD 0.37fF
C4019 vcm_commonmode a_42466_18528# 0.87fF
C4020 a_1761_2767# VDD 1.02fF
C4021 a_27314_67214# a_27406_67214# 0.32fF
C4022 vcm_commonmode a_32334_61190# 0.31fF
C4023 vcm_commonmode a_22386_24552# 0.84fF
C4024 a_7939_30503# a_19626_31751# 0.42fF
C4025 a_44474_71230# a_44474_70226# 1.00fF
C4026 a_2872_44111# a_27627_51733# 0.35fF
C4027 a_6831_63303# a_14831_50095# 1.43fF
C4028 a_8123_28879# VDD 0.35fF
C4029 a_33430_62194# ctopp 3.59fF
C4030 a_14287_51175# a_4674_40277# 0.35fF
C4031 a_8531_70543# a_23830_49525# 0.42fF
C4032 a_29414_70226# VDD 0.51fF
C4033 a_18151_52263# a_24394_58178# 0.38fF
C4034 a_12343_36893# VDD 0.50fF
C4035 a_39299_48783# a_44474_65206# 0.38fF
C4036 vcm_commonmode a_24394_57174# 0.87fF
C4037 a_20359_29199# a_19807_28111# 1.65fF
C4038 a_12985_16367# VDD 6.95fF
C4039 vcm_commonmode a_36350_70226# 0.31fF
C4040 a_32426_72234# a_32426_71230# 1.00fF
C4041 a_1768_16367# a_2052_38377# 0.65fF
C4042 a_40458_20536# a_41462_20536# 0.97fF
C4043 a_7571_26151# a_9751_25071# 0.68fF
C4044 a_17366_24552# m3_17268_24414# 2.81fF
C4045 a_29414_63198# a_30418_63198# 0.97fF
C4046 vcm_commonmode a_17274_16886# 0.33fF
C4047 a_2004_42453# a_1761_40847# 0.98fF
C4048 a_3668_56311# a_5595_63125# 0.64fF
C4049 a_39454_71230# ctopp 3.40fF
C4050 ctopn a_35438_20536# 3.59fF
C4051 a_2235_30503# a_13390_29575# 0.41fF
C4052 a_22291_29415# a_12447_29199# 0.62fF
C4053 a_29322_58178# a_29414_58178# 0.32fF
C4054 a_4215_51157# VDD 13.53fF
C4055 a_10515_63143# a_17488_48731# 0.33fF
C4056 a_28756_7638# a_28410_16520# 0.38fF
C4057 a_49494_10496# a_49494_9492# 1.00fF
C4058 a_24302_9858# a_24394_9492# 0.32fF
C4059 a_10055_58791# a_36797_27497# 0.41fF
C4060 a_3215_68351# VDD 0.44fF
C4061 a_47486_8488# VDD 0.58fF
C4062 a_7571_29199# a_5363_30503# 0.34fF
C4063 vcm_commonmode a_38450_62194# 0.87fF
C4064 a_3023_16341# a_2873_13879# 0.38fF
C4065 a_40366_16886# a_40458_16520# 0.32fF
C4066 a_39222_48169# a_40458_57174# 0.38fF
C4067 a_40050_48463# a_45478_70226# 0.38fF
C4068 a_4482_57863# a_2606_41079# 0.42fF
C4069 a_23736_7638# a_23390_9492# 0.38fF
C4070 a_18370_58178# VDD 0.52fF
C4071 a_23390_59182# a_24394_59182# 0.97fF
C4072 a_13867_38870# a_13669_38517# 0.31fF
C4073 a_7295_44647# a_33694_30761# 0.54fF
C4074 a_25493_29967# VDD 0.48fF
C4075 vcm_commonmode a_46482_15516# 0.87fF
C4076 ctopn a_35438_12504# 3.59fF
C4077 vcm_commonmode a_25306_58178# 0.31fF
C4078 a_43362_28879# a_47486_66210# 0.38fF
C4079 a_21382_17524# a_22386_17524# 0.97fF
C4080 a_12549_35836# a_13743_35836# 2.01fF
C4081 a_12641_36596# a_1761_32143# 0.96fF
C4082 a_32370_50871# VDD 0.34fF
C4083 vcm_commonmode a_44474_71230# 0.86fF
C4084 a_38450_21540# a_38450_20536# 1.00fF
C4085 a_4903_23983# VDD 0.43fF
C4086 a_25398_24552# a_25398_23548# 1.00fF
C4087 a_27752_7638# a_27406_20536# 0.38fF
C4088 a_35438_67214# VDD 0.51fF
C4089 a_40458_12504# a_41462_12504# 0.97fF
C4090 a_46390_67214# a_46482_67214# 0.32fF
C4091 a_23395_52047# a_2775_46025# 0.82fF
C4092 a_43267_31055# a_46482_62194# 0.38fF
C4093 a_41261_28335# ctopp 2.63fF
C4094 ctopn a_30418_21540# 3.59fF
C4095 a_16746_13506# VDD 33.20fF
C4096 vcm_commonmode a_42374_67214# 0.31fF
C4097 a_14287_51175# a_7862_34025# 1.19fF
C4098 a_13925_51727# a_14859_51183# 0.33fF
C4099 a_15607_46805# a_33839_28309# 0.61fF
C4100 vcm_commonmode a_23390_13508# 0.87fF
C4101 a_10515_22671# a_12257_56623# 23.52fF
C4102 a_10575_69439# VDD 0.37fF
C4103 a_12355_65103# a_15439_49525# 1.36fF
C4104 a_11619_56615# a_12341_3311# 1.52fF
C4105 a_42466_68218# ctopp 3.59fF
C4106 ctopn a_35438_17524# 3.59fF
C4107 a_32426_9492# VDD 0.51fF
C4108 a_48490_16520# VDD 0.55fF
C4109 a_27752_7638# a_27406_12504# 0.38fF
C4110 a_32334_7850# a_32426_7484# 0.32fF
C4111 vcm_commonmode a_39362_9858# 0.31fF
C4112 a_11067_13095# a_10055_58791# 1.57fF
C4113 a_48490_63198# a_49494_63198# 0.97fF
C4114 vcm_commonmode a_19282_22910# 0.31fF
C4115 a_32121_42369# VDD 1.79fF
C4116 a_16746_69224# a_12901_66959# 0.41fF
C4117 a_32951_27247# a_33430_10496# 0.38fF
C4118 a_22386_18528# a_22386_17524# 1.00fF
C4119 a_3339_43023# a_26550_40871# 0.65fF
C4120 a_6671_51183# VDD 0.37fF
C4121 a_35438_21540# a_36442_21540# 0.97fF
C4122 a_8273_42479# a_9405_31599# 0.53fF
C4123 a_43378_9858# a_43470_9492# 0.32fF
C4124 a_26310_64202# a_26402_64202# 0.32fF
C4125 a_27183_34789# VDD 0.92fF
C4126 a_40458_7484# VDD 1.25fF
C4127 vcm_commonmode a_47486_68218# 0.87fF
C4128 a_42466_59182# a_43470_59182# 0.97fF
C4129 a_6467_55527# a_27793_51733# 0.79fF
C4130 a_23298_22910# a_23390_22544# 0.32fF
C4131 a_27752_7638# a_27406_17524# 0.38fF
C4132 a_34434_64202# VDD 0.51fF
C4133 a_2411_26133# a_1761_30511# 0.64fF
C4134 a_24959_30503# a_32823_29397# 0.39fF
C4135 a_27422_29789# VDD 0.30fF
C4136 a_42466_56170# ctopp 3.40fF
C4137 a_1586_66567# VDD 6.15fF
C4138 a_23390_14512# a_23390_13508# 1.00fF
C4139 ctopn a_36442_18528# 3.59fF
C4140 vcm_commonmode a_41370_64202# 0.31fF
C4141 a_2689_65103# a_1923_59583# 0.31fF
C4142 a_40458_17524# a_41462_17524# 0.97fF
C4143 a_48490_72234# a_49494_72234# 0.97fF
C4144 a_1923_73087# a_4351_67279# 0.51fF
C4145 a_29760_7638# a_29414_15516# 0.38fF
C4146 m2_48260_24282# inn_analog 0.73fF
C4147 a_27406_60186# a_28410_60186# 0.97fF
C4148 a_44474_24552# a_44474_23548# 1.00fF
C4149 a_11067_46823# a_33694_30761# 0.30fF
C4150 a_29414_12504# a_29414_11500# 1.00fF
C4151 a_15548_30761# VDD 5.36fF
C4152 a_1803_19087# a_2339_38129# 2.23fF
C4153 a_43267_31055# a_12981_59343# 0.40fF
C4154 vcm_commonmode a_20286_23914# 0.31fF
C4155 a_16746_71232# ctopp 1.36fF
C4156 a_18197_44220# VDD 0.87fF
C4157 vcm_commonmode a_17274_66210# 0.33fF
C4158 a_21371_50959# a_12983_63151# 0.40fF
C4159 a_22386_18528# a_23390_18528# 0.97fF
C4160 a_2012_33927# a_1915_35015# 0.89fF
C4161 a_22386_19532# VDD 0.51fF
C4162 a_41462_61190# ctopp 3.59fF
C4163 ctopn a_45478_10496# 3.59fF
C4164 a_43470_69222# VDD 0.51fF
C4165 a_1761_31055# VDD 9.05fF
C4166 vcm_commonmode a_29322_19898# 0.31fF
C4167 a_4535_43567# a_4701_43567# 0.69fF
C4168 a_23395_52047# a_12981_62313# 0.40fF
C4169 vcm_commonmode a_47486_56170# 0.87fF
C4170 a_16362_15516# VDD 2.47fF
C4171 a_20359_29199# a_29927_29199# 9.26fF
C4172 a_10515_63143# a_8273_42479# 1.34fF
C4173 vcm_commonmode a_30418_8488# 0.86fF
C4174 a_41462_65206# VDD 0.51fF
C4175 a_15439_49525# ctopp 1.54fF
C4176 a_22632_41831# a_23415_41263# 0.32fF
C4177 a_19282_14878# a_19374_14512# 0.32fF
C4178 a_12251_39069# VDD 1.86fF
C4179 a_45478_70226# ctopp 3.58fF
C4180 a_20378_72234# m3_20280_72146# 2.80fF
C4181 a_13909_41923# VDD 8.15fF
C4182 a_35346_69222# a_35438_69222# 0.32fF
C4183 vcm_commonmode a_48398_65206# 0.31fF
C4184 a_41462_18528# a_41462_17524# 1.00fF
C4185 a_12641_36596# a_12663_35431# 3.03fF
C4186 a_19720_7638# a_12727_15529# 0.41fF
C4187 a_30326_24918# VDD 0.36fF
C4188 a_12947_8725# a_16362_8488# 1.25fF
C4189 a_45386_64202# a_45478_64202# 0.32fF
C4190 a_4259_32687# VDD 0.36fF
C4191 ctopn a_40458_15516# 3.59fF
C4192 vcm_commonmode a_46482_61190# 0.87fF
C4193 a_46482_14512# VDD 0.51fF
C4194 a_1757_45205# VDD 0.61fF
C4195 a_16746_70228# a_16362_70226# 2.28fF
C4196 a_29760_55394# a_12727_67753# 0.40fF
C4197 vcm_commonmode a_18370_67214# 0.88fF
C4198 a_1683_27399# config_2_in[1] 0.40fF
C4199 a_25398_20536# VDD 0.51fF
C4200 a_40366_55166# VDD 0.35fF
C4201 a_42374_22910# a_42466_22544# 0.32fF
C4202 a_20359_29199# a_28817_29111# 0.38fF
C4203 a_31422_10496# a_32426_10496# 0.97fF
C4204 a_77451_38925# a_76971_38925# 1285.84fF
C4205 a_12516_7093# a_11251_59879# 0.60fF
C4206 a_33338_65206# a_33430_65206# 0.32fF
C4207 a_42466_14512# a_42466_13508# 1.00fF
C4208 vcm_commonmode a_32334_20902# 0.31fF
C4209 a_1761_39215# VDD 5.63fF
C4210 vcm_commonmode a_21290_63198# 0.31fF
C4211 a_38115_52263# a_18979_30287# 5.65fF
C4212 a_46482_60186# a_47486_60186# 0.97fF
C4213 a_34434_58178# ctopp 3.59fF
C4214 a_24302_23914# a_24394_23548# 0.32fF
C4215 a_48490_66210# VDD 0.54fF
C4216 a_10975_66407# a_10515_22671# 8.12fF
C4217 a_17366_11500# a_18370_11500# 0.97fF
C4218 a_48490_12504# a_48490_11500# 1.00fF
C4219 vcm_commonmode a_31422_16520# 0.87fF
C4220 ctopn a_17366_13508# 3.43fF
C4221 a_36613_48169# a_22843_29415# 0.39fF
C4222 a_1761_43567# a_24029_39355# 4.48fF
C4223 a_18611_52047# VDD 15.05fF
C4224 a_21290_66210# a_21382_66210# 0.32fF
C4225 a_47486_7484# m3_47388_7346# 2.80fF
C4226 a_2011_34837# a_2317_28892# 0.68fF
C4227 a_25398_12504# VDD 0.51fF
C4228 a_36392_43677# VDD 1.68fF
C4229 a_35438_70226# a_35438_69222# 1.00fF
C4230 a_4119_70741# a_2840_66103# 0.38fF
C4231 a_2952_66139# a_5024_67885# 0.65fF
C4232 a_41462_18528# a_42466_18528# 0.97fF
C4233 vcm_commonmode a_28756_55394# 10.02fF
C4234 a_6921_72943# a_5877_70197# 0.79fF
C4235 a_6559_59879# a_18335_50645# 0.70fF
C4236 a_24740_7638# a_12985_16367# 0.41fF
C4237 a_15607_46805# a_26350_28585# 0.32fF
C4238 a_8453_51727# VDD 1.69fF
C4239 a_44474_55166# m3_44376_55078# 2.81fF
C4240 vcm_commonmode a_32334_12870# 0.31fF
C4241 a_21382_24552# a_22386_24552# 0.97fF
C4242 a_16891_35561# VDD 0.66fF
C4243 a_27535_30503# a_8491_41383# 1.45fF
C4244 a_31768_55394# a_12901_66959# 0.40fF
C4245 a_33338_19898# a_33430_19532# 0.32fF
C4246 a_18151_52263# a_7598_36103# 0.74fF
C4247 a_20378_21540# VDD 0.51fF
C4248 vcm_commonmode a_23390_7484# 0.69fF
C4249 a_6467_55527# a_19478_51959# 1.90fF
C4250 a_12202_54599# a_12818_52521# 0.52fF
C4251 a_18370_62194# a_19374_62194# 0.97fF
C4252 a_34434_11500# a_34434_10496# 1.00fF
C4253 a_41427_52263# a_12907_27023# 0.64fF
C4254 a_3339_43023# a_5085_23047# 1.92fF
C4255 a_36717_47375# a_36442_59182# 0.38fF
C4256 a_1929_12131# a_3983_12879# 0.56fF
C4257 a_38358_14878# a_38450_14512# 0.32fF
C4258 vcm_commonmode a_27314_21906# 0.31fF
C4259 a_21382_69222# ctopp 3.59fF
C4260 a_7255_10357# VDD 0.42fF
C4261 a_25221_41281# VDD 1.61fF
C4262 vcm_commonmode a_17366_64202# 1.83fF
C4263 vcm_commonmode a_45386_58178# 0.31fF
C4264 a_25398_17524# VDD 0.51fF
C4265 vcm_commonmode m2_48260_24282# 0.46fF
C4266 a_39454_72234# a_40458_72234# 0.97fF
C4267 a_17274_20902# a_17366_20536# 0.32fF
C4268 a_40491_27247# a_12727_15529# 0.41fF
C4269 a_1689_10396# a_2223_28617# 0.86fF
C4270 a_1761_39215# a_33486_34191# 0.71fF
C4271 a_28757_27247# VDD 4.42fF
C4272 vcm_commonmode a_32334_17890# 0.31fF
C4273 a_12355_15055# a_7461_27247# 0.46fF
C4274 a_19374_65206# ctopp 3.59fF
C4275 a_23390_57174# a_24394_57174# 0.97fF
C4276 a_18611_52047# a_23390_61190# 0.38fF
C4277 vcm_commonmode a_19282_60186# 0.31fF
C4278 a_26402_15516# a_27406_15516# 0.97fF
C4279 a_30035_44581# VDD 0.78fF
C4280 a_5147_19605# VDD 0.47fF
C4281 a_11067_63143# a_11251_59879# 1.61fF
C4282 a_3143_22364# VDD 2.81fF
C4283 a_37039_36919# VDD 0.65fF
C4284 a_1689_10396# a_1887_12342# 0.31fF
C4285 a_36613_48169# a_37446_64202# 0.38fF
C4286 a_13183_52047# a_17366_63198# 0.42fF
C4287 a_16746_16518# a_12727_13353# 2.28fF
C4288 vcm_commonmode a_26402_69222# 0.87fF
C4289 a_24394_71230# a_25398_71230# 0.97fF
C4290 a_46482_59182# VDD 0.51fF
C4291 a_28756_7638# a_12895_13967# 0.41fF
C4292 a_43378_23914# a_43470_23548# 0.32fF
C4293 a_2787_32679# a_3607_34639# 0.63fF
C4294 ctopn inn_analog 1.63fF
C4295 a_33515_30511# VDD 0.51fF
C4296 a_36442_11500# a_37446_11500# 0.97fF
C4297 a_34251_52263# a_11067_46823# 1.58fF
C4298 a_6162_28487# a_4351_26703# 0.85fF
C4299 a_40366_66210# a_40458_66210# 0.32fF
C4300 a_1929_10651# a_1929_12131# 2.12fF
C4301 vcm_commonmode a_33430_22544# 0.87fF
C4302 a_3339_32463# a_12447_29199# 0.38fF
C4303 a_18979_30287# a_20267_30503# 1.85fF
C4304 a_6579_42255# VDD 0.36fF
C4305 a_34251_52263# a_12355_65103# 0.40fF
C4306 vcm_commonmode a_24394_65206# 0.87fF
C4307 a_32971_35281# a_13097_36367# 0.31fF
C4308 a_26402_18528# VDD 0.51fF
C4309 a_16746_61192# VDD 33.19fF
C4310 a_1799_29556# a_2011_34837# 0.63fF
C4311 ctopn a_24394_8488# 3.40fF
C4312 a_40458_24552# a_41462_24552# 0.97fF
C4313 a_7580_61751# a_4298_58951# 0.39fF
C4314 a_17274_12870# a_17366_12504# 0.32fF
C4315 a_16707_34473# VDD 0.61fF
C4316 vcm_commonmode a_33338_18894# 0.31fF
C4317 a_26402_66210# ctopp 3.59fF
C4318 ctopn a_12877_14441# 3.23fF
C4319 a_26221_29423# a_27234_29789# 0.35fF
C4320 a_2959_47113# a_10687_52553# 0.66fF
C4321 a_42718_27497# a_44474_19532# 0.38fF
C4322 a_6467_55527# a_7210_55081# 0.65fF
C4323 a_37446_62194# a_38450_62194# 0.97fF
C4324 a_2317_28892# VDD 5.98fF
C4325 a_8082_56775# VDD 0.32fF
C4326 vcm_commonmode a_29414_14512# 0.87fF
C4327 a_16955_52047# a_20378_58178# 0.38fF
C4328 a_31059_38007# VDD 0.63fF
C4329 a_1768_13103# a_1586_21959# 0.32fF
C4330 vcm_commonmode a_24302_55166# 0.30fF
C4331 a_35438_10496# VDD 0.51fF
C4332 a_3759_39991# VDD 0.66fF
C4333 a_39222_48169# a_40458_65206# 0.38fF
C4334 a_9135_49557# a_9301_49557# 0.42fF
C4335 a_5363_16367# VDD 0.50fF
C4336 a_28410_72234# a_28410_71230# 1.00fF
C4337 a_36350_20902# a_36442_20536# 0.32fF
C4338 vcm_commonmode a_42374_10862# 0.31fF
C4339 a_25306_63198# a_25398_63198# 0.32fF
C4340 a_12947_56817# a_16362_56170# 19.83fF
C4341 a_42466_57174# a_43470_57174# 0.97fF
C4342 a_7925_72399# VDD 1.12fF
C4343 a_45478_15516# a_46482_15516# 0.97fF
C4344 vcm_commonmode a_34434_23548# 0.87fF
C4345 a_2787_30503# a_12935_31287# 0.39fF
C4346 vcm_commonmode a_31422_66210# 0.87fF
C4347 a_15557_52245# VDD 0.39fF
C4348 a_3751_72373# a_2686_70223# 1.27fF
C4349 a_22386_62194# VDD 0.51fF
C4350 a_8273_42479# a_9135_29423# 0.65fF
C4351 a_27406_55166# m3_27308_55078# 2.81fF
C4352 vcm_commonmode a_43470_19532# 0.87fF
C4353 ctopn a_25398_16520# 3.59fF
C4354 vcm_commonmode a_29322_62194# 0.31fF
C4355 a_36717_47375# a_36442_57174# 0.38fF
C4356 a_30418_15516# VDD 0.51fF
C4357 a_25879_48169# VDD 0.30fF
C4358 a_41427_52263# a_41462_70226# 0.38fF
C4359 a_43470_71230# a_44474_71230# 0.97fF
C4360 a_11803_55311# a_12516_7093# 1.15fF
C4361 a_19282_59182# a_19374_59182# 0.32fF
C4362 a_4792_20443# VDD 5.86fF
C4363 m3_46384_7346# VDD 0.33fF
C4364 a_29927_29199# a_28446_31375# 1.96fF
C4365 a_8485_29673# VDD 1.43fF
C4366 vcm_commonmode a_37354_15882# 0.31fF
C4367 a_30418_63198# ctopp 3.64fF
C4368 a_13183_52047# a_24209_48463# 0.43fF
C4369 a_28410_71230# VDD 0.58fF
C4370 a_40458_11500# VDD 0.51fF
C4371 a_30023_41959# VDD 2.22fF
C4372 a_41872_29423# a_43470_66210# 0.38fF
C4373 a_17274_17890# a_17366_17524# 0.32fF
C4374 a_5533_17455# VDD 0.59fF
C4375 vcm_commonmode a_35346_71230# 0.31fF
C4376 a_44474_24552# VDD 0.60fF
C4377 vcm_commonmode a_47394_11866# 0.31fF
C4378 a_24394_59182# ctopp 3.59fF
C4379 a_17712_7638# a_11067_21583# 0.40fF
C4380 a_4443_46607# a_1761_32143# 0.80fF
C4381 a_23390_64202# a_23390_63198# 1.23fF
C4382 a_36350_12870# a_36442_12504# 0.32fF
C4383 a_17191_32117# VDD 0.31fF
C4384 a_10515_63143# a_6835_46823# 1.14fF
C4385 a_41261_28335# a_42466_62194# 0.38fF
C4386 a_34251_52263# ctopp 2.62fF
C4387 a_25321_29673# a_26505_31599# 0.31fF
C4388 a_1586_45431# a_1591_45205# 0.80fF
C4389 a_5715_44343# VDD 0.63fF
C4390 a_31422_59182# a_31422_58178# 1.00fF
C4391 a_12869_2741# a_11067_46823# 0.52fF
C4392 a_5441_72399# a_5599_74549# 0.40fF
C4393 a_2411_19605# a_1586_18695# 0.37fF
C4394 a_13643_28327# a_12899_2767# 0.60fF
C4395 a_46482_57174# VDD 0.51fF
C4396 a_10055_58791# a_26748_7638# 0.41fF
C4397 a_12355_65103# a_12869_2741# 0.57fF
C4398 a_3668_56311# a_4758_45369# 2.60fF
C4399 a_22386_13508# a_23390_13508# 0.97fF
C4400 vcm_commonmode a_46482_20536# 0.87fF
C4401 a_39223_32463# a_29175_28335# 0.43fF
C4402 a_1799_29556# VDD 6.60fF
C4403 vcm_commonmode a_35438_63198# 0.92fF
C4404 a_27406_68218# a_28410_68218# 0.97fF
C4405 a_12381_35836# a_5595_33205# 0.52fF
C4406 a_32856_48463# VDD 1.04fF
C4407 a_1923_73087# a_1591_69141# 0.34fF
C4408 vcm_commonmode ctopn 97.04fF
C4409 a_4149_65327# VDD 0.66fF
C4410 a_39454_56170# a_39454_55166# 1.00fF
C4411 a_44382_63198# a_44474_63198# 0.32fF
C4412 a_1761_41935# a_1761_40847# 1.30fF
C4413 a_35438_57174# a_35438_56170# 1.00fF
C4414 vcm_commonmode a_29414_59182# 0.87fF
C4415 a_10956_14459# a_10995_14333# 0.65fF
C4416 a_2787_30503# a_12999_29423# 0.45fF
C4417 a_4351_67279# a_11710_58487# 1.38fF
C4418 a_35039_51335# VDD 0.68fF
C4419 a_31330_21906# a_31422_21540# 0.32fF
C4420 a_12546_22351# a_2143_15271# 0.98fF
C4421 a_7571_26151# a_10873_27497# 0.42fF
C4422 a_10286_26311# VDD 1.11fF
C4423 vcm_commonmode a_46482_12504# 0.87fF
C4424 a_28410_60186# ctopp 3.59fF
C4425 ctopn a_47486_9492# 3.57fF
C4426 a_2840_66103# a_15261_51433# 0.34fF
C4427 a_31422_68218# VDD 0.51fF
C4428 a_9491_12297# a_9484_11989# 0.31fF
C4429 a_2503_34319# VDD 0.36fF
C4430 a_31330_7850# VDD 0.61fF
C4431 a_49402_58178# a_49494_58178# 0.32fF
C4432 a_11803_55311# a_11067_63143# 0.67fF
C4433 a_19374_16520# a_19374_15516# 1.00fF
C4434 ctopn a_27406_22544# 3.58fF
C4435 a_3339_30503# a_8461_32937# 0.31fF
C4436 a_1586_45431# a_4674_40277# 0.44fF
C4437 vcm_commonmode a_38358_68218# 0.31fF
C4438 a_38358_59182# a_38450_59182# 0.32fF
C4439 a_14289_29687# VDD 0.30fF
C4440 a_10515_22671# a_8739_28879# 0.31fF
C4441 a_11067_66191# a_12355_15055# 2.32fF
C4442 vcm_commonmode a_41462_21540# 0.87fF
C4443 a_9503_26151# a_20378_8488# 0.38fF
C4444 a_36350_17890# a_36442_17524# 0.32fF
C4445 a_27869_50095# a_29561_49667# 0.30fF
C4446 a_20359_29199# VDD 11.11fF
C4447 a_45386_72234# a_45478_72234# 0.32fF
C4448 a_16955_52047# a_11803_55311# 1.18fF
C4449 a_36797_27497# a_12877_14441# 0.41fF
C4450 a_8583_33551# a_22291_29415# 0.94fF
C4451 a_23298_60186# a_23390_60186# 0.32fF
C4452 vcm_commonmode a_18370_10496# 0.88fF
C4453 a_19720_7638# a_19374_21540# 0.38fF
C4454 a_18703_29199# a_7862_34025# 0.32fF
C4455 a_7773_63927# a_3295_62083# 0.46fF
C4456 a_42466_64202# a_42466_63198# 1.23fF
C4457 a_1683_31599# VDD 0.43fF
C4458 vcm_commonmode a_46482_17524# 0.87fF
C4459 ctopn a_23390_14512# 3.59fF
C4460 a_39389_52271# a_12981_59343# 0.40fF
C4461 vcm_commonmode a_33430_60186# 0.87fF
C4462 a_45478_13508# VDD 0.51fF
C4463 a_14287_51175# a_12983_63151# 0.40fF
C4464 a_18278_18894# a_18370_18528# 0.32fF
C4465 a_1761_27791# a_2223_28617# 0.46fF
C4466 a_16152_37601# a_25133_37571# 0.55fF
C4467 a_8162_53609# VDD 0.34fF
C4468 a_2451_72373# a_2843_71829# 0.44fF
C4469 a_34434_22544# a_34434_21540# 1.00fF
C4470 a_11763_62581# VDD 0.40fF
C4471 a_12641_37684# a_12473_37429# 1.68fF
C4472 a_31422_56170# VDD 0.52fF
C4473 a_1923_59583# a_1823_62589# 0.39fF
C4474 a_41462_13508# a_42466_13508# 0.97fF
C4475 a_19096_36513# VDD 1.63fF
C4476 a_16955_52047# a_12981_62313# 0.40fF
C4477 a_46482_68218# a_47486_68218# 0.97fF
C4478 vcm_commonmode a_38358_56170# 0.31fF
C4479 ctopn a_28410_23548# 3.40fF
C4480 a_2872_44111# a_1761_25071# 0.35fF
C4481 a_7519_59575# a_8199_58229# 1.74fF
C4482 vcm_commonmode a_21290_8854# 0.31fF
C4483 a_29760_7638# a_29414_20536# 0.38fF
C4484 a_25787_28327# a_16863_29415# 1.89fF
C4485 a_39223_32463# a_39454_22544# 0.38fF
C4486 a_24394_57174# ctopp 3.58fF
C4487 a_27406_56170# a_28410_56170# 0.97fF
C4488 a_2847_71615# VDD 0.46fF
C4489 ctopn a_37446_19532# 3.59fF
C4490 a_30788_28487# a_30891_28309# 0.80fF
C4491 a_16746_11498# VDD 33.20fF
C4492 a_17599_52263# a_22386_72234# 0.34fF
C4493 a_4298_58951# a_7933_51433# 0.42fF
C4494 a_30418_61190# VDD 0.51fF
C4495 vcm_commonmode a_23390_11500# 0.87fF
C4496 a_31422_58178# a_31422_57174# 1.00fF
C4497 a_16863_29415# a_2235_30503# 0.37fF
C4498 vcm_commonmode a_47486_18528# 0.87fF
C4499 a_9529_28335# a_12631_28585# 1.26fF
C4500 a_1954_61677# a_1923_59583# 1.50fF
C4501 vcm_commonmode a_37354_61190# 0.31fF
C4502 a_38450_16520# a_38450_15516# 1.00fF
C4503 vcm_commonmode a_27406_24552# 0.84fF
C4504 a_17599_52263# a_12727_67753# 0.40fF
C4505 a_12907_56399# a_12901_66959# 0.41fF
C4506 a_43362_28879# a_47486_69222# 0.38fF
C4507 a_23390_19532# a_23390_18528# 1.00fF
C4508 a_29760_7638# a_29414_12504# 0.38fF
C4509 a_40675_27791# a_12899_10927# 0.41fF
C4510 a_6417_62215# a_6559_59879# 0.47fF
C4511 a_27314_10862# a_27406_10496# 0.32fF
C4512 a_38450_62194# ctopp 3.59fF
C4513 a_3668_56311# a_4240_53083# 1.48fF
C4514 a_34434_70226# VDD 0.51fF
C4515 vcm_commonmode a_37446_55166# 0.84fF
C4516 a_1761_47919# a_6473_40277# 0.43fF
C4517 vcm_commonmode a_29414_57174# 0.87fF
C4518 a_15660_49257# VDD 0.35fF
C4519 vcm_commonmode a_41370_70226# 0.31fF
C4520 a_42374_60186# a_42466_60186# 0.32fF
C4521 a_10055_58791# a_4298_58951# 0.32fF
C4522 VDD config_1_in[11] 1.00fF
C4523 vcm_commonmode a_22294_16886# 0.31fF
C4524 a_25971_52263# a_22843_29415# 2.71fF
C4525 a_28099_42895# a_30023_41959# 0.69fF
C4526 a_10969_71631# VDD 0.50fF
C4527 a_16746_66212# a_16362_66210# 2.28fF
C4528 a_18370_15516# a_18370_14512# 1.00fF
C4529 a_44474_71230# ctopp 3.40fF
C4530 ctopn a_40458_20536# 3.59fF
C4531 a_40458_7484# m3_40360_7346# 2.80fF
C4532 a_21675_43447# VDD 0.63fF
C4533 a_37354_18894# a_37446_18528# 0.32fF
C4534 a_1761_37039# a_13097_36367# 0.79fF
C4535 vcm_commonmode a_17507_52047# 10.02fF
C4536 a_29760_7638# a_29414_17524# 0.38fF
C4537 a_1823_76181# a_2952_66139# 0.58fF
C4538 a_26402_61190# a_27406_61190# 0.97fF
C4539 a_37446_55166# m3_37348_55078# 2.81fF
C4540 a_17274_24918# a_17366_24552# 0.32fF
C4541 a_13716_43047# a_16152_43677# 0.84fF
C4542 a_32426_68218# a_32426_67214# 1.00fF
C4543 vcm_commonmode a_43470_62194# 0.87fF
C4544 vcm_commonmode a_36797_27497# 10.35fF
C4545 a_18151_52263# a_12901_66959# 0.40fF
C4546 a_23390_58178# VDD 0.51fF
C4547 a_10055_58791# a_43269_29967# 0.41fF
C4548 a_10975_66407# a_7377_18012# 0.93fF
C4549 ctopn a_40458_12504# 3.59fF
C4550 a_46482_56170# a_47486_56170# 0.97fF
C4551 vcm_commonmode a_30326_58178# 0.31fF
C4552 a_28547_51175# a_32426_59182# 0.38fF
C4553 a_7987_40821# VDD 0.62fF
C4554 a_17366_69222# a_17366_68218# 1.00fF
C4555 a_13097_36367# a_1761_32143# 1.61fF
C4556 a_16362_17524# VDD 2.47fF
C4557 vcm_commonmode a_49494_71230# 0.89fF
C4558 a_25971_52263# a_41872_29423# 9.36fF
C4559 a_28547_51175# a_41427_52263# 0.46fF
C4560 a_36717_47375# a_36613_48169# 0.39fF
C4561 a_9411_60437# VDD 0.43fF
C4562 a_1761_27791# a_1761_34319# 3.16fF
C4563 a_4758_45369# a_4891_47388# 0.50fF
C4564 a_29414_8488# a_30418_8488# 0.97fF
C4565 a_28318_55166# a_28410_55166# 0.32fF
C4566 a_40458_67214# VDD 0.51fF
C4567 a_19282_57174# a_19374_57174# 0.32fF
C4568 a_8059_74746# VDD 0.47fF
C4569 a_19720_55394# a_19374_61190# 0.38fF
C4570 a_22294_15882# a_22386_15516# 0.32fF
C4571 ctopn a_35438_21540# 3.59fF
C4572 a_30052_32117# a_30788_28487# 0.40fF
C4573 vcm_commonmode a_47394_67214# 0.31fF
C4574 a_30418_70226# a_31422_70226# 0.97fF
C4575 a_42466_19532# a_42466_18528# 1.00fF
C4576 a_46390_10862# a_46482_10496# 0.32fF
C4577 vcm_commonmode a_28410_13508# 0.87fF
C4578 a_37919_28111# a_38450_24552# 0.47fF
C4579 a_4307_67477# VDD 2.18fF
C4580 a_21479_36965# VDD 1.05fF
C4581 a_47486_68218# ctopp 3.58fF
C4582 ctopn a_40458_17524# 3.59fF
C4583 a_1761_47919# a_30855_41809# 0.73fF
C4584 a_1761_44111# a_2021_17973# 0.37fF
C4585 a_37446_9492# VDD 0.51fF
C4586 a_25787_28327# a_33430_64202# 0.38fF
C4587 a_11067_67279# a_11067_23759# 0.58fF
C4588 a_20359_29199# a_34482_29941# 0.47fF
C4589 vcm_commonmode a_17274_69222# 0.33fF
C4590 a_20286_71230# a_20378_71230# 0.32fF
C4591 a_28410_60186# a_28410_59182# 1.00fF
C4592 a_17366_22544# VDD 0.58fF
C4593 vcm_commonmode a_44382_9858# 0.31fF
C4594 m3_16264_59094# VDD 0.34fF
C4595 a_15607_46805# a_30788_28487# 0.64fF
C4596 a_17366_63198# a_17366_62194# 1.00fF
C4597 a_1770_14441# a_2419_48783# 2.32fF
C4598 a_32334_11866# a_32426_11500# 0.32fF
C4599 a_11067_67279# a_16362_20536# 1.27fF
C4600 a_12899_3311# a_40491_27247# 0.52fF
C4601 a_44474_72234# VDD 1.25fF
C4602 a_43362_28879# a_12727_58255# 0.40fF
C4603 a_37446_15516# a_37446_14512# 1.00fF
C4604 vcm_commonmode a_24302_22910# 0.31fF
C4605 vcm_commonmode a_11067_13095# 1.41fF
C4606 a_28756_55394# a_12355_65103# 0.40fF
C4607 a_32772_7638# a_12727_15529# 0.41fF
C4608 a_45478_61190# a_46482_61190# 0.97fF
C4609 a_22386_9492# a_22386_8488# 1.00fF
C4610 a_27752_7638# a_27406_21540# 0.38fF
C4611 a_36350_24918# a_36442_24552# 0.32fF
C4612 a_30764_7638# a_30418_23548# 0.38fF
C4613 a_1923_59583# a_1586_51335# 0.31fF
C4614 a_4248_29967# a_6066_28309# 0.31fF
C4615 a_45478_7484# VDD 1.65fF
C4616 a_17366_67214# a_18370_67214# 0.97fF
C4617 a_6467_55527# a_32582_51701# 0.66fF
C4618 a_36797_27497# a_37446_19532# 0.38fF
C4619 a_39454_64202# VDD 0.51fF
C4620 a_33338_62194# a_33430_62194# 0.32fF
C4621 vcm_commonmode a_20286_14878# 0.31fF
C4622 ctopn a_17366_11500# 3.43fF
C4623 a_47486_56170# ctopp 3.39fF
C4624 a_10699_69679# VDD 0.42fF
C4625 ctopn a_41462_18528# 3.59fF
C4626 vcm_commonmode a_16362_55166# 1.87fF
C4627 a_30967_41001# VDD 0.61fF
C4628 a_3024_67191# a_7155_55509# 0.70fF
C4629 a_36717_47375# a_36442_65206# 0.38fF
C4630 a_36442_69222# a_36442_68218# 1.00fF
C4631 vcm_commonmode a_46390_64202# 0.31fF
C4632 a_24394_72234# a_24394_71230# 1.00fF
C4633 vcm_commonmode a_17366_70226# 1.83fF
C4634 a_32951_27247# a_33430_15516# 0.38fF
C4635 a_5363_30503# a_15548_30761# 0.62fF
C4636 a_2959_47113# a_1923_54591# 0.33fF
C4637 a_48490_8488# a_49494_8488# 0.97fF
C4638 a_26402_8488# a_26402_7484# 1.00fF
C4639 a_46390_55166# a_46482_55166# 0.32fF
C4640 a_18370_23548# VDD 0.52fF
C4641 a_12355_15055# a_16362_62194# 19.89fF
C4642 a_28446_31375# VDD 4.88fF
C4643 a_1761_43567# a_15397_39631# 0.53fF
C4644 a_38358_57174# a_38450_57174# 0.32fF
C4645 a_6835_73193# VDD 0.67fF
C4646 a_1586_66567# a_9319_62613# 0.71fF
C4647 a_41370_15882# a_41462_15516# 0.32fF
C4648 vcm_commonmode a_25306_23914# 0.31fF
C4649 ctopn a_16746_20534# 1.68fF
C4650 a_8583_33551# a_13484_39325# 0.45fF
C4651 a_12357_37999# VDD 9.98fF
C4652 vcm_commonmode a_22294_66210# 0.31fF
C4653 a_19374_58178# a_20378_58178# 0.97fF
C4654 a_27406_19532# VDD 0.51fF
C4655 a_20635_29415# a_28756_7638# 0.52fF
C4656 a_20378_55166# m3_20280_55078# 2.81fF
C4657 a_10515_63143# a_5963_20149# 0.30fF
C4658 a_46482_61190# ctopp 3.59fF
C4659 a_40491_27247# a_43470_24552# 0.52fF
C4660 a_48490_69222# VDD 0.55fF
C4661 a_1823_66941# a_2959_47113# 0.34fF
C4662 a_1823_65853# a_3016_60949# 1.25fF
C4663 vcm_commonmode a_34342_19898# 0.31fF
C4664 a_18370_67214# ctopp 3.58fF
C4665 ctopn a_16362_16520# 1.35fF
C4666 a_30418_16520# a_31422_16520# 0.97fF
C4667 a_28547_51175# a_32426_57174# 0.38fF
C4668 a_22015_28111# a_15607_46805# 2.35fF
C4669 a_36613_48169# a_37446_70226# 0.38fF
C4670 a_39362_71230# a_39454_71230# 0.32fF
C4671 a_47486_60186# a_47486_59182# 1.00fF
C4672 vcm_commonmode a_35438_8488# 0.86fF
C4673 m3_18272_7346# VDD 0.34fF
C4674 a_46482_65206# VDD 0.51fF
C4675 a_22843_29415# a_25493_29967# 0.64fF
C4676 a_3339_32463# a_7695_31573# 0.39fF
C4677 a_36442_63198# a_36442_62194# 1.00fF
C4678 ctopn a_16746_12502# 1.68fF
C4679 a_3325_18543# a_3972_25615# 0.79fF
C4680 a_1761_40847# a_1895_40516# 0.34fF
C4681 a_5631_38127# VDD 2.76fF
C4682 a_23390_72234# m3_23292_72146# 2.80fF
C4683 a_17983_41855# VDD 0.85fF
C4684 a_39389_52271# a_39454_66210# 0.38fF
C4685 a_12967_50943# VDD 0.41fF
C4686 a_37919_28111# a_12727_15529# 0.41fF
C4687 a_35346_24918# VDD 0.36fF
C4688 a_41462_9492# a_41462_8488# 1.00fF
C4689 a_17712_7638# a_12546_22351# 0.40fF
C4690 a_16362_67214# VDD 2.48fF
C4691 ctopn a_45478_15516# 3.59fF
C4692 a_38557_32143# a_38450_62194# 0.38fF
C4693 a_36442_67214# a_37446_67214# 0.97fF
C4694 a_28756_55394# ctopp 2.62fF
C4695 a_15607_46805# a_37557_32463# 0.55fF
C4696 vcm_commonmode a_23390_67214# 0.87fF
C4697 a_30418_20536# VDD 0.51fF
C4698 a_27627_51733# a_27793_51733# 0.42fF
C4699 a_45386_55166# VDD 0.35fF
C4700 a_19374_63198# VDD 0.57fF
C4701 a_16510_8760# a_12899_10927# 1.09fF
C4702 a_3668_56311# a_3016_60949# 0.47fF
C4703 a_30591_37455# VDD 0.41fF
C4704 a_18278_13874# a_18370_13508# 0.32fF
C4705 vcm_commonmode a_37354_20902# 0.31fF
C4706 a_12355_65103# a_7479_54439# 0.60fF
C4707 ctopn a_12899_11471# 3.23fF
C4708 a_1761_22895# a_1761_44111# 1.77fF
C4709 vcm_commonmode a_26310_63198# 0.31fF
C4710 a_23298_68218# a_23390_68218# 0.32fF
C4711 a_4811_34855# a_7939_30503# 1.38fF
C4712 a_3618_58487# VDD 0.35fF
C4713 a_12727_58255# a_16362_59182# 1.15fF
C4714 a_45478_8488# a_45478_7484# 1.00fF
C4715 a_22386_7484# a_23390_7484# 0.97fF
C4716 vcm_commonmode a_20378_9492# 0.87fF
C4717 a_1823_63677# a_2959_47113# 0.82fF
C4718 a_20911_31055# VDD 0.38fF
C4719 vcm_commonmode a_36442_16520# 0.87fF
C4720 a_17366_64202# ctopp 3.43fF
C4721 ctopn a_22386_13508# 3.59fF
C4722 a_23192_27791# a_24768_27247# 0.37fF
C4723 vcm_commonmode a_20286_59182# 0.31fF
C4724 VDD result_out[5] 0.66fF
C4725 a_11067_67279# a_27752_7638# 0.41fF
C4726 a_30052_32117# a_23736_7638# 0.60fF
C4727 a_30418_12504# VDD 0.51fF
C4728 a_7295_44647# a_8491_41383# 1.93fF
C4729 a_7571_68047# a_4307_67477# 0.31fF
C4730 a_4075_18543# VDD 0.43fF
C4731 a_4351_26703# VDD 2.37fF
C4732 a_33430_9492# a_34434_9492# 0.97fF
C4733 a_3339_43023# VDD 48.50fF
C4734 vcm_commonmode a_37354_12870# 0.31fF
C4735 a_4891_47388# a_8123_56399# 0.44fF
C4736 a_9135_27239# a_21382_23548# 0.38fF
C4737 a_4443_46607# a_4495_35925# 0.44fF
C4738 a_34434_13508# a_34434_12504# 1.00fF
C4739 a_26523_29199# a_26350_28585# 0.48fF
C4740 a_1586_66567# a_4339_64521# 0.76fF
C4741 VDD result_out[14] 0.87fF
C4742 a_25398_21540# VDD 0.51fF
C4743 vcm_commonmode a_28410_7484# 0.68fF
C4744 a_17712_7638# a_17366_19532# 0.38fF
C4745 a_40675_27791# a_41462_19532# 0.38fF
C4746 a_2411_26133# a_2216_28309# 0.72fF
C4747 a_11430_26159# a_10964_25615# 1.09fF
C4748 a_1768_16367# a_1823_63677# 1.12fF
C4749 vcm_commonmode a_32334_21906# 0.31fF
C4750 a_26402_69222# ctopp 3.59fF
C4751 a_35647_41317# VDD 0.94fF
C4752 vcm_commonmode a_22386_64202# 0.87fF
C4753 a_30418_17524# VDD 0.51fF
C4754 a_17366_60186# VDD 0.57fF
C4755 a_1761_25071# a_2223_28617# 0.81fF
C4756 a_1591_23445# VDD 0.36fF
C4757 vcm_commonmode a_37354_17890# 0.31fF
C4758 a_24394_65206# ctopp 3.59fF
C4759 a_28756_55394# a_30762_49641# 0.37fF
C4760 a_6098_73095# VDD 1.32fF
C4761 a_28547_51175# a_12981_59343# 0.40fF
C4762 vcm_commonmode a_24302_60186# 0.31fF
C4763 a_24394_67214# a_24394_66210# 1.00fF
C4764 a_35815_31751# a_39223_32463# 0.75fF
C4765 a_18703_29199# a_20267_30503# 0.50fF
C4766 a_1586_45431# a_3987_19623# 0.58fF
C4767 a_12473_37429# a_25517_37455# 0.79fF
C4768 a_9668_51451# a_9707_51325# 0.46fF
C4769 a_10055_58791# a_12985_19087# 1.02fF
C4770 a_3016_60949# a_3141_59887# 0.56fF
C4771 a_11602_25071# VDD 1.25fF
C4772 a_4443_46607# a_13123_38231# 0.40fF
C4773 a_20378_65206# a_20378_64202# 1.00fF
C4774 a_37354_13874# a_37446_13508# 0.32fF
C4775 a_1689_10396# a_1803_19087# 0.73fF
C4776 a_42374_68218# a_42466_68218# 0.32fF
C4777 a_43267_31055# a_12516_7093# 0.40fF
C4778 vcm_commonmode a_31422_69222# 0.87fF
C4779 a_41462_7484# a_42466_7484# 0.97fF
C4780 a_15439_49525# a_2872_44111# 0.42fF
C4781 a_34482_29941# a_28446_31375# 0.51fF
C4782 a_24959_30503# a_28757_27247# 0.59fF
C4783 a_1586_21959# a_2411_19605# 0.57fF
C4784 a_11602_25071# a_11866_27791# 0.76fF
C4785 a_6473_40277# a_6671_40630# 0.31fF
C4786 a_23298_56170# a_23390_56170# 0.32fF
C4787 a_7803_55509# a_6515_62037# 1.10fF
C4788 vcm_commonmode a_38450_22544# 0.87fF
C4789 a_4811_34855# a_28305_28879# 0.60fF
C4790 a_3417_10927# VDD 0.47fF
C4791 a_18811_42405# VDD 0.84fF
C4792 vcm_commonmode a_29414_65206# 0.87fF
C4793 a_25398_69222# a_26402_69222# 0.97fF
C4794 a_31422_18528# VDD 0.51fF
C4795 a_30375_51335# VDD 0.51fF
C4796 a_8491_57487# a_6775_53877# 0.39fF
C4797 a_26748_7638# a_12877_14441# 0.41fF
C4798 a_20378_61190# a_20378_60186# 1.00fF
C4799 a_7111_22351# VDD 0.41fF
C4800 ctopn a_29414_8488# 3.40fF
C4801 a_35438_64202# a_36442_64202# 0.97fF
C4802 vcm_commonmode a_38358_18894# 0.31fF
C4803 a_31422_66210# ctopp 3.59fF
C4804 a_13067_38517# a_27271_37455# 0.61fF
C4805 vcm_commonmode a_18278_24918# 0.31fF
C4806 a_11067_46823# a_8491_41383# 2.11fF
C4807 a_15607_46805# a_22291_29415# 2.38fF
C4808 a_41872_29423# a_43470_69222# 0.38fF
C4809 a_22386_55166# VDD 0.60fF
C4810 a_32426_22544# a_33430_22544# 0.97fF
C4811 a_10680_52245# a_27333_52271# 0.58fF
C4812 a_6467_55527# a_2775_46025# 1.19fF
C4813 a_12631_28585# VDD 1.17fF
C4814 a_12257_56623# VDD 7.40fF
C4815 vcm_commonmode a_34434_14512# 0.87fF
C4816 a_23390_65206# a_24394_65206# 0.97fF
C4817 a_39247_38007# VDD 0.62fF
C4818 a_11067_67279# a_8491_27023# 0.42fF
C4819 vcm_commonmode a_29322_55166# 0.30fF
C4820 a_40458_10496# VDD 0.51fF
C4821 a_11947_68279# a_11999_67477# 0.38fF
C4822 a_19374_17524# a_19374_16520# 1.00fF
C4823 vcm_commonmode a_20286_57174# 0.31fF
C4824 a_11067_47695# a_1586_18695# 0.79fF
C4825 vcm_commonmode a_47394_10862# 0.31fF
C4826 a_23390_56170# a_23390_55166# 1.00fF
C4827 a_43470_67214# a_43470_66210# 1.00fF
C4828 vcm_commonmode a_10515_22671# 6.27fF
C4829 vcm_commonmode a_39454_23548# 0.87fF
C4830 a_33430_7484# m3_33332_7346# 2.80fF
C4831 a_35815_31751# a_32970_31145# 0.44fF
C4832 a_7295_43031# VDD 0.32fF
C4833 vcm_commonmode a_36442_66210# 0.87fF
C4834 a_36797_27497# a_12899_11471# 0.41fF
C4835 a_27406_62194# VDD 0.51fF
C4836 a_22294_61190# a_22386_61190# 0.32fF
C4837 a_7580_61751# VDD 2.73fF
C4838 a_6515_62037# a_6831_63303# 0.40fF
C4839 a_39454_65206# a_39454_64202# 1.00fF
C4840 vcm_commonmode a_48490_19532# 0.87fF
C4841 ctopn a_30418_16520# 3.59fF
C4842 a_12725_44527# a_12473_42869# 1.24fF
C4843 vcm_commonmode a_34342_62194# 0.31fF
C4844 a_12546_22351# a_16746_9490# 0.41fF
C4845 a_35438_15516# VDD 0.51fF
C4846 a_23390_19532# a_24394_19532# 0.97fF
C4847 a_33430_23548# a_33430_22544# 1.00fF
C4848 a_2021_22325# a_3607_34639# 0.74fF
C4849 vcm_commonmode a_42374_15882# 0.31fF
C4850 a_35438_63198# ctopp 3.64fF
C4851 a_42374_56170# a_42466_56170# 0.32fF
C4852 a_33430_71230# VDD 0.58fF
C4853 a_27406_66210# a_27406_65206# 1.00fF
C4854 a_28756_55394# a_28410_59182# 0.38fF
C4855 a_28410_14512# a_29414_14512# 0.97fF
C4856 a_33543_39095# VDD 0.67fF
C4857 a_45478_11500# VDD 0.51fF
C4858 a_38011_42035# VDD 2.15fF
C4859 a_11053_69135# a_11710_58487# 0.52fF
C4860 a_44474_69222# a_45478_69222# 0.97fF
C4861 ctopp ctopn 1.94fF
C4862 vcm_commonmode a_40366_71230# 0.31fF
C4863 a_32426_72234# a_33430_72234# 0.97fF
C4864 a_8583_33551# a_12907_27023# 1.27fF
C4865 a_39454_61190# a_39454_60186# 1.00fF
C4866 a_25306_8854# a_25398_8488# 0.32fF
C4867 a_29414_59182# ctopp 3.59fF
C4868 a_28547_51175# a_37534_51701# 0.63fF
C4869 a_11803_55311# a_6467_55527# 0.52fF
C4870 a_7999_13083# VDD 1.05fF
C4871 a_1586_40455# a_1778_42631# 1.01fF
C4872 a_26310_70226# a_26402_70226# 0.32fF
C4873 a_4215_51157# a_24683_51183# 0.35fF
C4874 a_25744_7638# a_12899_10927# 0.41fF
C4875 a_25398_62194# a_25398_61190# 1.00fF
C4876 a_18126_28023# VDD 0.43fF
C4877 vcm_commonmode a_19282_13874# 0.31fF
C4878 a_42466_65206# a_43470_65206# 0.97fF
C4879 a_5963_36585# VDD 1.93fF
C4880 a_39055_39913# VDD 0.59fF
C4881 a_29760_55394# a_29414_64202# 0.38fF
C4882 vcm_commonmode a_40458_63198# 0.92fF
C4883 a_38450_17524# a_38450_16520# 1.00fF
C4884 vcm_commonmode a_26748_7638# 10.35fF
C4885 a_25398_20536# a_25398_19532# 1.00fF
C4886 m3_46384_72146# VDD 0.33fF
C4887 a_33430_23548# a_34434_23548# 0.97fF
C4888 a_12641_42036# a_19967_41781# 0.45fF
C4889 a_37446_72234# VDD 1.63fF
C4890 a_30418_66210# a_31422_66210# 0.97fF
C4891 a_39222_48169# a_12727_58255# 0.40fF
C4892 vcm_commonmode a_34434_59182# 0.87fF
C4893 a_11619_56615# a_12257_56623# 0.74fF
C4894 a_8197_31599# a_10506_29967# 1.17fF
C4895 vcm_commonmode m3_16264_63110# 3.21fF
C4896 a_23507_43177# VDD 0.59fF
C4897 a_17507_52047# a_12355_65103# 0.40fF
C4898 a_31768_7638# a_31422_8488# 0.38fF
C4899 a_49494_14512# m3_49396_14374# 2.78fF
C4900 vcm_commonmode a_42466_72234# 0.69fF
C4901 a_7467_61751# VDD 0.50fF
C4902 a_41370_61190# a_41462_61190# 0.32fF
C4903 a_33430_60186# ctopp 3.59fF
C4904 a_36442_68218# VDD 0.51fF
C4905 a_14039_34743# VDD 0.61fF
C4906 a_1823_63677# a_2589_55535# 0.37fF
C4907 a_13005_43983# a_12713_43011# 0.40fF
C4908 a_36350_7850# VDD 0.62fF
C4909 a_12907_56399# a_15439_49525# 0.32fF
C4910 ctopn a_32426_22544# 3.58fF
C4911 a_7862_34025# a_2787_30503# 3.42fF
C4912 a_32856_48463# a_24959_30503# 0.50fF
C4913 a_4057_13647# VDD 0.39fF
C4914 a_38805_47081# VDD 0.38fF
C4915 vcm_commonmode a_43378_68218# 0.31fF
C4916 a_30418_71230# a_30418_70226# 1.00fF
C4917 a_4891_47388# a_1761_49007# 0.36fF
C4918 a_42466_19532# a_43470_19532# 0.97fF
C4919 a_42188_37149# a_41636_37601# 0.37fF
C4920 a_19576_51701# a_19478_51959# 2.55fF
C4921 a_12355_15055# a_9301_49557# 0.47fF
C4922 a_8531_70543# VDD 7.95fF
C4923 a_46482_66210# a_46482_65206# 1.00fF
C4924 a_47486_14512# a_48490_14512# 0.97fF
C4925 vcm_commonmode a_46482_21540# 0.87fF
C4926 a_30788_28487# a_28841_29575# 0.47fF
C4927 a_16746_10494# VDD 33.20fF
C4928 a_28547_51175# a_32426_65206# 0.38fF
C4929 a_27535_30503# a_19807_28111# 2.54fF
C4930 a_43362_28879# a_47486_72234# 0.34fF
C4931 a_20378_72234# a_20378_71230# 1.00fF
C4932 a_26402_20536# a_27406_20536# 0.97fF
C4933 a_44382_8854# a_44474_8488# 0.32fF
C4934 vcm_commonmode a_23390_10496# 0.87fF
C4935 a_10975_66407# VDD 12.74fF
C4936 a_16746_63200# a_15439_49525# 2.24fF
C4937 a_7571_31599# VDD 0.67fF
C4938 ctopn a_28410_14512# 3.59fF
C4939 a_13067_38517# a_12801_38517# 1.69fF
C4940 vcm_commonmode a_38450_60186# 0.87fF
C4941 a_48490_56170# m2_48260_54946# 0.98fF
C4942 a_42985_46831# a_48490_68218# 0.38fF
C4943 a_45386_70226# a_45478_70226# 0.32fF
C4944 a_13123_38231# a_13097_36367# 0.92fF
C4945 a_2559_52789# VDD 0.34fF
C4946 a_1923_73087# a_2163_73085# 0.64fF
C4947 a_43269_29967# a_12877_14441# 0.41fF
C4948 a_12907_27023# a_14471_28585# 0.40fF
C4949 a_44474_62194# a_44474_61190# 1.00fF
C4950 a_35438_10496# a_35438_9492# 1.00fF
C4951 a_36442_56170# VDD 0.52fF
C4952 a_2124_64507# a_2163_64381# 0.79fF
C4953 a_29545_35841# VDD 1.24fF
C4954 a_25971_52263# a_8295_47388# 3.35fF
C4955 a_19374_8488# VDD 0.58fF
C4956 a_26310_16886# a_26402_16520# 0.32fF
C4957 vcm_commonmode a_43378_56170# 0.31fF
C4958 a_28756_55394# a_28410_57174# 0.38fF
C4959 ctopn a_33430_23548# 3.51fF
C4960 a_20359_29199# a_24959_30503# 0.73fF
C4961 a_25787_28327# a_33430_70226# 0.38fF
C4962 a_44474_20536# a_44474_19532# 1.00fF
C4963 a_4792_58371# VDD 0.53fF
C4964 vcm_commonmode a_26310_8854# 0.31fF
C4965 a_3016_60949# a_5541_53609# 0.32fF
C4966 a_32951_27247# a_33430_20536# 0.38fF
C4967 a_13643_28327# a_32823_29397# 0.32fF
C4968 vcm_commonmode a_18370_15516# 0.88fF
C4969 a_36613_48169# a_13643_28327# 0.33fF
C4970 a_29414_57174# ctopp 3.58fF
C4971 a_1761_52815# a_7598_36103# 0.74fF
C4972 a_12355_65103# a_11067_13095# 23.58fF
C4973 a_43267_31055# a_46482_60186# 0.38fF
C4974 ctopn a_42466_19532# 3.59fF
C4975 a_32970_31145# a_33641_29967# 0.73fF
C4976 vcm_commonmode m3_16264_10358# 3.21fF
C4977 a_34251_52263# a_35438_66210# 0.38fF
C4978 a_7571_16917# a_7737_16917# 0.42fF
C4979 a_3247_20495# a_4792_20443# 0.69fF
C4980 a_26397_51183# a_20359_29199# 0.64fF
C4981 vcm_commonmode a_12901_66665# 6.22fF
C4982 a_24394_21540# a_24394_20536# 1.00fF
C4983 a_35438_61190# VDD 0.51fF
C4984 vcm_commonmode a_28410_11500# 0.87fF
C4985 a_26402_12504# a_27406_12504# 0.97fF
C4986 a_5449_25071# a_4528_26159# 0.31fF
C4987 a_5831_39189# a_4941_35727# 0.44fF
C4988 a_34780_56398# a_34434_62194# 0.38fF
C4989 vcm_commonmode a_42374_61190# 0.31fF
C4990 a_32334_67214# a_32426_67214# 0.32fF
C4991 vcm_commonmode a_32426_24552# 0.84fF
C4992 a_42985_46831# a_48490_56170# 0.42fF
C4993 a_17507_52047# ctopp 2.62fF
C4994 a_49494_71230# a_49494_70226# 1.00fF
C4995 a_32951_27247# a_33430_12504# 0.38fF
C4996 a_3339_43023# a_12663_40871# 0.47fF
C4997 a_2959_47113# a_4215_51157# 0.61fF
C4998 a_43470_62194# ctopp 3.59fF
C4999 a_39454_70226# VDD 0.51fF
C5000 vcm_commonmode a_42466_55166# 0.84fF
C5001 vcm_commonmode a_16362_63198# 4.47fF
C5002 vcm_commonmode a_34434_57174# 0.87fF
C5003 a_20378_16520# VDD 0.51fF
C5004 a_16587_49007# VDD 0.46fF
C5005 vcm_commonmode a_46390_70226# 0.31fF
C5006 a_45478_20536# a_46482_20536# 0.97fF
C5007 a_2124_54715# a_2163_54589# 0.79fF
C5008 a_18278_7850# a_18370_7484# 0.32fF
C5009 a_29760_7638# a_29414_21540# 0.38fF
C5010 VDD config_1_in[6] 0.95fF
C5011 a_34434_63198# a_35438_63198# 0.97fF
C5012 a_14361_29967# VDD 0.72fF
C5013 vcm_commonmode a_27314_16886# 0.31fF
C5014 ctopn a_45478_20536# 3.59fF
C5015 a_3607_34639# a_5087_29423# 1.04fF
C5016 a_42709_29199# a_48490_9492# 0.38fF
C5017 a_34342_58178# a_34434_58178# 0.32fF
C5018 a_7933_51433# VDD 0.61fF
C5019 a_2686_70223# a_5877_70197# 0.42fF
C5020 a_32951_27247# a_33430_17524# 0.38fF
C5021 a_21382_21540# a_22386_21540# 0.97fF
C5022 a_29322_9858# a_29414_9492# 0.32fF
C5023 a_5336_54965# VDD 0.77fF
C5024 a_5211_24759# a_5531_22895# 0.72fF
C5025 a_1761_46287# a_15459_41781# 2.62fF
C5026 vcm_commonmode a_48490_62194# 0.87fF
C5027 a_45386_16886# a_45478_16520# 0.32fF
C5028 vcm_commonmode a_19374_68218# 0.87fF
C5029 a_28410_58178# VDD 0.51fF
C5030 a_28410_59182# a_29414_59182# 0.97fF
C5031 a_16362_21540# VDD 2.47fF
C5032 a_36629_27791# a_36442_19532# 0.38fF
C5033 a_8295_47388# a_12341_3311# 0.52fF
C5034 ctopn a_45478_12504# 3.59fF
C5035 a_42985_46831# a_12901_58799# 0.40fF
C5036 vcm_commonmode a_35346_58178# 0.31fF
C5037 a_1761_50639# a_13576_40413# 0.95fF
C5038 a_21049_41245# VDD 0.88fF
C5039 a_26402_17524# a_27406_17524# 0.97fF
C5040 vcm_commonmode a_43269_29967# 10.42fF
C5041 a_12621_36091# a_14258_34191# 2.27fF
C5042 a_22843_29415# a_20359_29199# 0.38fF
C5043 a_23535_50247# VDD 0.40fF
C5044 a_38358_72234# a_38450_72234# 0.32fF
C5045 a_8491_57487# a_2872_44111# 0.98fF
C5046 a_43470_21540# a_43470_20536# 1.00fF
C5047 a_10055_58791# VDD 17.88fF
C5048 a_30418_24552# a_30418_23548# 1.00fF
C5049 a_45478_67214# VDD 0.51fF
C5050 a_20359_29199# a_23395_32463# 0.50fF
C5051 a_12869_2741# a_12899_3855# 2.92fF
C5052 a_45478_12504# a_46482_12504# 0.97fF
C5053 a_11067_13095# ctopp 1.70fF
C5054 a_12889_40977# a_12343_42333# 0.43fF
C5055 a_1591_72943# VDD 0.79fF
C5056 a_21371_50959# a_12981_59343# 0.40fF
C5057 ctopn a_40458_21540# 3.59fF
C5058 a_32367_28309# a_30788_28487# 2.39fF
C5059 a_7281_29423# a_8197_31599# 0.41fF
C5060 a_15607_46805# a_3339_32463# 0.45fF
C5061 a_19559_44535# VDD 0.58fF
C5062 a_43269_29967# a_47486_9492# 0.38fF
C5063 a_3325_49551# VDD 2.39fF
C5064 vcm_commonmode a_33430_13508# 0.87fF
C5065 ctopn a_17366_10496# 3.43fF
C5066 a_39673_28111# a_40458_24552# 0.46fF
C5067 a_11067_13095# a_16746_64204# 0.37fF
C5068 a_2099_59861# a_2473_34293# 0.65fF
C5069 ctopn a_45478_17524# 3.59fF
C5070 a_42466_9492# VDD 0.51fF
C5071 vcm_commonmode a_19374_56170# 0.87fF
C5072 a_43362_28879# a_47486_58178# 0.38fF
C5073 a_27535_30503# a_29927_29199# 1.27fF
C5074 vcm_commonmode a_22294_69222# 0.31fF
C5075 a_39389_52271# a_12516_7093# 0.40fF
C5076 a_30764_7638# a_30418_14512# 0.38fF
C5077 a_37354_7850# a_37446_7484# 0.32fF
C5078 a_22386_22544# VDD 0.51fF
C5079 vcm_commonmode a_49402_9858# 0.30fF
C5080 a_17651_30485# VDD 0.74fF
C5081 a_48398_72234# VDD 0.62fF
C5082 a_11067_67279# a_11067_63143# 0.39fF
C5083 vcm_commonmode a_29322_22910# 0.31fF
C5084 a_17366_70226# ctopp 3.42fF
C5085 a_30788_28487# a_26523_29199# 0.44fF
C5086 a_3316_42313# VDD 0.31fF
C5087 vcm_commonmode a_20286_65206# 0.31fF
C5088 a_21290_69222# a_21382_69222# 0.32fF
C5089 a_27406_18528# a_27406_17524# 1.00fF
C5090 a_1761_37039# a_1761_32143# 2.37fF
C5091 a_16219_51183# VDD 0.39fF
C5092 a_13183_52047# a_17599_52263# 0.50fF
C5093 a_17712_7638# a_12985_16367# 0.40fF
C5094 a_40458_21540# a_41462_21540# 0.97fF
C5095 a_12231_60949# VDD 0.37fF
C5096 a_48398_9858# a_48490_9492# 0.32fF
C5097 a_23736_7638# a_23390_19532# 0.38fF
C5098 a_20635_29415# a_4811_34855# 0.61fF
C5099 a_31330_64202# a_31422_64202# 0.32fF
C5100 a_1681_5175# VDD 0.85fF
C5101 vcm_commonmode a_18370_61190# 0.88fF
C5102 a_21187_29415# a_20267_30503# 1.07fF
C5103 a_18370_14512# VDD 0.52fF
C5104 a_39389_52271# a_39454_69222# 0.38fF
C5105 a_47486_59182# a_48490_59182# 0.97fF
C5106 a_28318_22910# a_28410_22544# 0.32fF
C5107 a_44474_64202# VDD 0.51fF
C5108 a_1761_40847# a_13669_37429# 3.03fF
C5109 a_20359_29199# a_41334_29575# 0.46fF
C5110 a_17366_10496# a_18370_10496# 0.97fF
C5111 vcm_commonmode a_25306_14878# 0.31fF
C5112 ctopn a_22386_11500# 3.59fF
C5113 a_49876_41198# a_51330_39932# 0.30fF
C5114 a_19282_65206# a_19374_65206# 0.32fF
C5115 a_28410_14512# a_28410_13508# 1.00fF
C5116 ctopn a_46482_18528# 3.59fF
C5117 a_4842_45467# a_5173_44655# 0.34fF
C5118 a_76346_40594# VDD 1.01fF
C5119 a_1586_66567# a_1768_16367# 0.83fF
C5120 a_45478_17524# a_46482_17524# 0.97fF
C5121 a_38115_52263# a_26523_28111# 0.84fF
C5122 vcm_commonmode a_22386_70226# 0.87fF
C5123 a_39454_58178# vcm_commonmode 0.87fF
C5124 a_6559_22671# a_5211_24759# 0.38fF
C5125 a_32426_60186# a_33430_60186# 0.97fF
C5126 a_23390_23548# VDD 0.52fF
C5127 a_41967_31375# a_42466_18528# 0.38fF
C5128 a_20378_66210# VDD 0.51fF
C5129 a_6559_22671# a_1761_34319# 0.91fF
C5130 a_34434_12504# a_34434_11500# 1.00fF
C5131 vcm_commonmode a_30326_23914# 0.31fF
C5132 a_26402_7484# m3_26304_7346# 2.80fF
C5133 a_1761_49007# a_1761_44111# 2.17fF
C5134 a_39503_43957# VDD 0.45fF
C5135 vcm_commonmode a_27314_66210# 0.31fF
C5136 a_21382_70226# a_21382_69222# 1.00fF
C5137 a_2099_59861# a_1803_19087# 1.34fF
C5138 a_27406_18528# a_28410_18528# 0.97fF
C5139 a_32426_19532# VDD 0.51fF
C5140 a_11619_56615# a_10055_58791# 0.96fF
C5141 vcm_commonmode a_39362_19898# 0.31fF
C5142 a_23390_67214# ctopp 3.59fF
C5143 a_19282_19898# a_19374_19532# 0.32fF
C5144 vcm_commonmode a_40458_8488# 0.86fF
C5145 m3_33332_7346# VDD 0.41fF
C5146 a_1586_36727# a_1761_30511# 1.78fF
C5147 a_20378_11500# a_20378_10496# 1.00fF
C5148 a_8739_28879# VDD 0.35fF
C5149 a_20685_28335# a_17712_7638# 0.41fF
C5150 a_12263_4391# a_10515_23975# 0.72fF
C5151 a_2339_38129# config_2_in[3] 0.85fF
C5152 a_18151_52263# a_24394_59182# 0.38fF
C5153 a_40050_48463# a_10515_22671# 0.40fF
C5154 a_24302_14878# a_24394_14512# 0.32fF
C5155 a_20713_39105# VDD 1.71fF
C5156 a_26402_72234# m3_26304_72146# 2.80fF
C5157 a_4119_70741# a_6515_62037# 0.31fF
C5158 a_40366_69222# a_40458_69222# 0.32fF
C5159 a_46482_18528# a_46482_17524# 1.00fF
C5160 ctopn a_35601_27497# 2.62fF
C5161 a_18335_50645# VDD 0.45fF
C5162 a_29760_55394# a_25971_52263# 0.30fF
C5163 a_10515_63143# a_8491_41383# 1.51fF
C5164 a_18370_55166# a_19374_55166# 0.97fF
C5165 a_40366_24918# VDD 0.36fF
C5166 a_23192_27791# a_28817_29111# 0.34fF
C5167 a_1803_19087# a_1761_41935# 1.14fF
C5168 a_2021_22325# a_1761_40847# 0.80fF
C5169 ctopn a_12985_7663# 3.23fF
C5170 a_2235_30503# a_16228_28335# 0.50fF
C5171 vcm_commonmode a_28410_67214# 0.87fF
C5172 a_35438_20536# VDD 0.51fF
C5173 a_2451_72373# a_5483_74244# 0.52fF
C5174 a_47394_22910# a_47486_22544# 0.32fF
C5175 a_26748_7638# a_12899_11471# 0.41fF
C5176 a_24394_63198# VDD 0.57fF
C5177 a_12907_27023# a_32038_29575# 0.67fF
C5178 a_49494_22544# m3_49396_22406# 2.78fF
C5179 a_36442_10496# a_37446_10496# 0.97fF
C5180 a_20027_27221# VDD 1.23fF
C5181 a_12907_56399# a_8491_57487# 0.44fF
C5182 a_38358_65206# a_38450_65206# 0.32fF
C5183 a_40737_37692# VDD 0.99fF
C5184 a_47486_14512# a_47486_13508# 1.00fF
C5185 vcm_commonmode a_42374_20902# 0.31fF
C5186 a_11719_28023# a_12631_28585# 0.77fF
C5187 a_21371_50959# a_25398_64202# 0.38fF
C5188 vcm_commonmode a_31330_63198# 0.31fF
C5189 a_2872_44111# a_2656_45895# 0.42fF
C5190 a_26610_49257# VDD 0.47fF
C5191 a_10515_22671# a_11067_46823# 0.41fF
C5192 a_11067_21583# a_12877_16911# 0.76fF
C5193 a_9135_27239# a_21382_14512# 0.38fF
C5194 a_18370_59182# VDD 0.52fF
C5195 vcm_commonmode a_25398_9492# 0.87fF
C5196 m3_18272_72146# VDD 0.34fF
C5197 a_29322_23914# a_29414_23548# 0.32fF
C5198 a_6559_22671# a_3339_30503# 0.64fF
C5199 a_12355_65103# a_10515_22671# 1.45fF
C5200 a_22386_11500# a_23390_11500# 0.97fF
C5201 vcm_commonmode a_41462_16520# 0.87fF
C5202 a_22386_64202# ctopp 3.59fF
C5203 ctopn a_27406_13508# 3.59fF
C5204 a_12473_41781# a_12713_41923# 0.94fF
C5205 a_30418_72234# VDD 1.37fF
C5206 vcm_commonmode a_25306_59182# 0.31fF
C5207 a_25787_28327# a_12727_58255# 0.40fF
C5208 a_26310_66210# a_26402_66210# 0.32fF
C5209 a_35438_12504# VDD 0.51fF
C5210 a_40458_70226# a_40458_69222# 1.00fF
C5211 a_46482_18528# a_47486_18528# 0.97fF
C5212 a_1761_37039# a_12663_35431# 0.92fF
C5213 a_13669_37429# a_32327_35839# 1.51fF
C5214 a_8111_18825# VDD 0.39fF
C5215 vcm_commonmode a_35438_72234# 0.69fF
C5216 a_6559_59663# a_10503_52828# 1.86fF
C5217 a_19720_7638# a_19374_16520# 0.38fF
C5218 a_6467_55527# a_5190_59575# 0.75fF
C5219 vcm_commonmode a_42374_12870# 0.31fF
C5220 a_26402_24552# a_27406_24552# 0.97fF
C5221 a_28756_7638# a_11067_21583# 0.41fF
C5222 a_2952_46805# a_2339_38129# 1.24fF
C5223 a_7000_43541# a_9945_47919# 0.60fF
C5224 a_12907_27023# a_15607_46805# 0.86fF
C5225 a_10475_14165# VDD 0.35fF
C5226 a_20543_46831# VDD 0.60fF
C5227 a_38358_19898# a_38450_19532# 0.32fF
C5228 a_30418_21540# VDD 0.51fF
C5229 vcm_commonmode a_33430_7484# 0.69fF
C5230 a_16362_22544# a_11067_21583# 1.27fF
C5231 a_12447_29199# a_13357_32143# 0.95fF
C5232 a_23390_62194# a_24394_62194# 0.97fF
C5233 a_39454_11500# a_39454_10496# 1.00fF
C5234 a_48490_58178# VDD 0.54fF
C5235 a_3301_26703# a_4571_26677# 1.05fF
C5236 a_1591_57711# VDD 2.78fF
C5237 a_43378_14878# a_43470_14512# 0.32fF
C5238 vcm_commonmode a_37354_21906# 0.31fF
C5239 a_31422_69222# ctopp 3.59fF
C5240 a_49494_72234# m3_49396_72146# 2.80fF
C5241 a_28756_55394# a_28410_65206# 0.38fF
C5242 vcm_commonmode a_27406_64202# 0.87fF
C5243 a_12663_35431# a_1761_32143# 0.30fF
C5244 a_13097_36367# a_31131_35281# 0.43fF
C5245 a_35438_17524# VDD 0.51fF
C5246 a_22294_20902# a_22386_20536# 0.32fF
C5247 a_22386_60186# VDD 0.51fF
C5248 a_7571_29199# a_11430_26159# 0.35fF
C5249 a_3339_43023# a_24959_30503# 0.88fF
C5250 a_36442_55166# a_37446_55166# 0.97fF
C5251 a_5839_22351# VDD 0.63fF
C5252 a_42718_27497# a_44474_22544# 0.38fF
C5253 a_22843_29415# a_28446_31375# 0.83fF
C5254 a_1823_63677# a_1952_60431# 2.52fF
C5255 a_6515_62037# a_1586_51335# 1.70fF
C5256 vcm_commonmode a_42374_17890# 0.31fF
C5257 a_29414_65206# ctopp 3.59fF
C5258 a_15661_29199# a_17869_28585# 0.81fF
C5259 a_49494_68218# m3_49396_68130# 2.78fF
C5260 a_28410_57174# a_29414_57174# 0.97fF
C5261 vcm_commonmode a_29322_60186# 0.31fF
C5262 a_31422_15516# a_32426_15516# 0.97fF
C5263 a_14646_29423# a_15548_30761# 0.36fF
C5264 a_5993_32687# a_5449_25071# 0.31fF
C5265 a_1803_20719# VDD 8.29fF
C5266 a_39299_48783# a_44474_68218# 0.38fF
C5267 a_13123_38231# a_32971_35281# 0.42fF
C5268 a_2007_51701# VDD 0.46fF
C5269 a_39223_32463# a_39454_13508# 0.38fF
C5270 a_2794_62697# VDD 1.25fF
C5271 a_10055_58791# a_24740_7638# 0.41fF
C5272 a_8491_27023# a_18370_24552# 0.42fF
C5273 a_25744_7638# a_25398_24552# 0.46fF
C5274 vcm_commonmode a_12985_19087# 6.30fF
C5275 a_18151_52263# a_12869_2741# 0.32fF
C5276 a_1761_25071# a_1803_19087# 2.47fF
C5277 a_18151_52263# a_24394_57174# 0.38fF
C5278 a_1757_14741# VDD 0.62fF
C5279 a_2606_41079# a_18413_47919# 0.38fF
C5280 a_29760_55394# a_29414_70226# 0.38fF
C5281 vcm_commonmode a_36442_69222# 0.87fF
C5282 a_29414_71230# a_30418_71230# 0.97fF
C5283 vcm_commonmode a_16746_8486# 5.34fF
C5284 a_39223_32463# a_12727_15529# 0.41fF
C5285 a_48398_23914# a_48490_23548# 0.32fF
C5286 a_41462_11500# a_42466_11500# 0.97fF
C5287 a_17507_30761# VDD 0.87fF
C5288 a_3295_62083# a_7265_56053# 0.32fF
C5289 a_41261_28335# a_42466_60186# 0.38fF
C5290 a_45386_66210# a_45478_66210# 0.32fF
C5291 vcm_commonmode a_43470_22544# 0.87fF
C5292 a_15851_27791# a_16101_31029# 0.31fF
C5293 a_23567_42035# VDD 1.87fF
C5294 vcm_commonmode a_34434_65206# 0.87fF
C5295 a_31768_55394# a_31422_66210# 0.38fF
C5296 a_7841_12167# a_31659_31751# 0.50fF
C5297 a_36442_18528# VDD 0.51fF
C5298 a_11067_13095# a_6269_43567# 0.65fF
C5299 a_16362_24552# VDD 1.16fF
C5300 vcm_commonmode a_19282_11866# 0.31fF
C5301 a_10515_22671# ctopp 3.22fF
C5302 ctopn a_34434_8488# 3.40fF
C5303 a_12907_56399# a_2021_22325# 0.30fF
C5304 a_45478_24552# a_46482_24552# 0.97fF
C5305 a_5254_67503# VDD 3.36fF
C5306 a_22294_12870# a_22386_12504# 0.32fF
C5307 vcm_commonmode a_43378_18894# 0.31fF
C5308 a_36442_66210# ctopp 3.59fF
C5309 a_25971_52263# a_30418_62194# 0.38fF
C5310 vcm_commonmode a_23298_24918# 0.31fF
C5311 a_39299_48783# a_44474_56170# 0.38fF
C5312 a_7000_43541# a_5831_39189# 0.39fF
C5313 a_17366_59182# a_17366_58178# 1.00fF
C5314 a_27406_55166# VDD 0.60fF
C5315 a_6831_63303# a_17682_50095# 1.08fF
C5316 a_36629_27791# a_12899_10927# 0.41fF
C5317 a_6816_19355# a_7377_18012# 0.92fF
C5318 a_22291_29415# a_26523_29199# 2.22fF
C5319 a_42466_62194# a_43470_62194# 0.97fF
C5320 a_18370_57174# VDD 0.52fF
C5321 vcm_commonmode a_39454_14512# 0.87fF
C5322 a_4571_26677# a_5211_24759# 0.67fF
C5323 vcm_commonmode a_18370_20536# 0.88fF
C5324 vcm_commonmode a_33430_55166# 0.84fF
C5325 a_8583_33551# a_13669_35253# 0.50fF
C5326 a_45478_10496# VDD 0.51fF
C5327 a_22411_40183# VDD 0.61fF
C5328 vcm_commonmode a_25306_57174# 0.31fF
C5329 a_40050_48463# a_12901_66665# 0.40fF
C5330 a_41370_20902# a_41462_20536# 0.32fF
C5331 a_11067_63143# a_1586_18695# 0.53fF
C5332 a_36797_27497# a_12985_7663# 0.41fF
C5333 a_30326_63198# a_30418_63198# 0.32fF
C5334 a_4351_67279# a_10687_52553# 4.63fF
C5335 a_14287_51175# a_4191_33449# 1.34fF
C5336 a_47486_57174# a_48490_57174# 0.97fF
C5337 a_21382_57174# a_21382_56170# 1.00fF
C5338 a_9183_72007# VDD 0.37fF
C5339 vcm_commonmode a_44474_23548# 0.87fF
C5340 a_7571_26151# a_8491_41383# 0.59fF
C5341 a_9484_11989# VDD 1.23fF
C5342 vcm_commonmode a_41462_66210# 0.87fF
C5343 a_17274_21906# a_17366_21540# 0.32fF
C5344 a_32426_62194# VDD 0.51fF
C5345 vcm_commonmode a_18370_12504# 0.88fF
C5346 ctopn a_19374_9492# 3.58fF
C5347 a_11067_13095# a_10515_63143# 4.47fF
C5348 a_11803_64239# a_11053_62607# 0.41fF
C5349 a_27563_35831# VDD 0.64fF
C5350 ctopn a_35438_16520# 3.59fF
C5351 a_3339_32463# a_2339_38129# 0.87fF
C5352 vcm_commonmode a_39362_62194# 0.31fF
C5353 a_2292_17179# a_1929_10651# 0.56fF
C5354 a_40458_15516# VDD 0.51fF
C5355 a_48490_71230# a_49494_71230# 0.97fF
C5356 a_3339_43023# a_3247_20495# 1.18fF
C5357 a_24302_59182# a_24394_59182# 0.32fF
C5358 a_43269_29967# a_12899_11471# 0.41fF
C5359 a_2840_53511# VDD 7.65fF
C5360 a_2012_33927# config_2_in[0] 0.81fF
C5361 vcm_commonmode a_47394_15882# 0.31fF
C5362 a_40458_63198# ctopp 3.64fF
C5363 a_1761_41935# a_14963_39783# 3.95fF
C5364 a_38450_71230# VDD 0.58fF
C5365 a_41427_52263# a_12901_58799# 0.40fF
C5366 a_22294_17890# a_22386_17524# 0.32fF
C5367 a_4495_35925# a_2235_30503# 0.44fF
C5368 a_2216_28309# a_3187_34293# 0.68fF
C5369 a_27535_30503# VDD 9.68fF
C5370 vcm_commonmode a_45386_71230# 0.31fF
C5371 a_4968_60405# VDD 1.00fF
C5372 a_34434_59182# ctopp 3.59fF
C5373 a_5211_24759# a_5963_20149# 0.36fF
C5374 a_28410_64202# a_28410_63198# 1.23fF
C5375 a_15080_32143# VDD 0.42fF
C5376 a_41370_12870# a_41462_12504# 0.32fF
C5377 vcm_commonmode a_18370_17524# 0.88fF
C5378 a_14287_51175# a_12981_59343# 0.40fF
C5379 a_11067_13095# a_3607_34639# 0.68fF
C5380 a_10975_66407# a_9307_30663# 1.05fF
C5381 a_7862_34025# a_10531_31055# 0.89fF
C5382 a_4443_46607# a_4674_40277# 1.12fF
C5383 a_17366_13508# VDD 0.57fF
C5384 a_14258_44527# VDD 1.58fF
C5385 a_36442_59182# a_36442_58178# 1.00fF
C5386 a_2959_47113# a_35039_51335# 0.56fF
C5387 a_27752_7638# a_27406_16520# 0.38fF
C5388 a_20378_22544# a_20378_21540# 1.00fF
C5389 vcm_commonmode a_24302_13874# 0.31fF
C5390 a_6559_59663# a_8123_56399# 2.00fF
C5391 a_14287_51175# a_12447_29199# 0.70fF
C5392 a_5211_24759# a_5085_24759# 2.44fF
C5393 a_11943_69367# VDD 0.39fF
C5394 a_6515_62037# a_7773_63927# 0.55fF
C5395 a_27406_13508# a_28410_13508# 0.97fF
C5396 a_39299_48783# a_12355_15055# 0.40fF
C5397 a_32426_68218# a_33430_68218# 0.97fF
C5398 vcm_commonmode a_45478_63198# 0.92fF
C5399 a_49402_16886# VDD 0.31fF
C5400 a_5239_48767# VDD 0.55fF
C5401 a_28547_51175# a_12516_7093# 0.40fF
C5402 a_1823_76181# a_6515_67477# 0.72fF
C5403 a_8999_61493# VDD 1.40fF
C5404 a_44474_56170# a_44474_55166# 1.00fF
C5405 a_46482_24552# m3_46384_24414# 2.81fF
C5406 a_49402_63198# a_49494_63198# 0.32fF
C5407 a_16955_52047# a_23774_49551# 0.63fF
C5408 a_40458_57174# a_40458_56170# 1.00fF
C5409 a_41370_72234# VDD 0.63fF
C5410 vcm_commonmode a_39454_59182# 0.87fF
C5411 a_12727_15529# a_16362_13508# 19.89fF
C5412 a_33727_43177# VDD 0.65fF
C5413 a_12901_66959# a_16362_69222# 19.89fF
C5414 a_9187_51157# VDD 0.39fF
C5415 a_36350_21906# a_36442_21540# 0.32fF
C5416 a_5405_25615# VDD 0.64fF
C5417 a_17366_58178# a_17366_57174# 1.00fF
C5418 a_38450_60186# ctopp 3.59fF
C5419 a_41462_68218# VDD 0.51fF
C5420 a_5831_39189# a_5915_35943# 1.59fF
C5421 vcm_commonmode a_19374_18528# 0.87fF
C5422 a_41370_7850# VDD 0.63fF
C5423 a_24394_16520# a_24394_15516# 1.00fF
C5424 ctopn a_37446_22544# 3.58fF
C5425 ctopn m3_32328_24414# 0.39fF
C5426 vcm_commonmode a_48398_68218# 0.31fF
C5427 a_34251_52263# a_35438_69222# 0.38fF
C5428 a_39223_32463# a_39454_7484# 0.34fF
C5429 a_43378_59182# a_43470_59182# 0.32fF
C5430 a_12355_65103# a_10407_47607# 0.37fF
C5431 a_23192_27791# VDD 3.45fF
C5432 a_4345_69679# VDD 0.35fF
C5433 a_2787_30503# a_9731_22895# 0.36fF
C5434 a_2927_39733# a_1689_10396# 0.30fF
C5435 a_41370_17890# a_41462_17524# 0.32fF
C5436 a_35601_27497# a_35438_8488# 0.38fF
C5437 a_49402_72234# a_49494_72234# 0.32fF
C5438 a_28318_60186# a_28410_60186# 0.32fF
C5439 vcm_commonmode a_28410_10496# 0.87fF
C5440 a_47486_64202# a_47486_63198# 1.23fF
C5441 ctopn a_33430_14512# 3.59fF
C5442 a_1586_21959# a_8491_27023# 0.61fF
C5443 vcm_commonmode a_43470_60186# 0.87fF
C5444 VDD inn_analog 9.83fF
C5445 a_12901_66665# ctopp 2.95fF
C5446 a_19374_7484# m3_19276_7346# 2.80fF
C5447 a_2292_43291# a_4535_43567# 0.35fF
C5448 a_23298_18894# a_23390_18528# 0.32fF
C5449 a_39454_22544# a_39454_21540# 1.00fF
C5450 a_9135_27239# a_12877_16911# 0.41fF
C5451 a_6417_62215# VDD 2.31fF
C5452 a_41462_56170# VDD 0.52fF
C5453 a_17366_55166# m3_17268_55078# 2.81fF
C5454 a_9670_24527# a_9263_24501# 0.34fF
C5455 a_46482_13508# a_47486_13508# 0.97fF
C5456 a_24394_8488# VDD 0.58fF
C5457 a_18370_68218# a_18370_67214# 1.00fF
C5458 a_41872_29423# a_12257_56623# 0.40fF
C5459 vcm_commonmode a_48398_56170# 0.31fF
C5460 ctopn a_38450_23548# 3.40fF
C5461 a_12877_14441# VDD 7.23fF
C5462 VDD config_2_in[7] 2.42fF
C5463 a_7050_53333# a_10503_52828# 0.52fF
C5464 vcm_commonmode a_31330_8854# 0.31fF
C5465 vcm_commonmode a_23390_15516# 0.87fF
C5466 a_16362_63198# ctopp 1.35fF
C5467 a_1586_21959# a_1757_23445# 0.60fF
C5468 a_34434_57174# ctopp 3.58fF
C5469 a_32426_56170# a_33430_56170# 0.97fF
C5470 a_38557_32143# a_10515_22671# 0.40fF
C5471 a_16955_52047# a_20378_59182# 0.38fF
C5472 ctopn a_47486_19532# 3.58fF
C5473 a_43270_27791# a_45478_9492# 0.38fF
C5474 a_12713_36483# a_13743_35836# 2.80fF
C5475 vcm_commonmode a_21382_71230# 0.86fF
C5476 a_25398_72234# a_26402_72234# 0.97fF
C5477 a_17599_52263# a_25971_52263# 0.38fF
C5478 a_40458_61190# VDD 0.51fF
C5479 VDD result_out[0] 0.74fF
C5480 vcm_commonmode a_33430_11500# 0.87fF
C5481 a_36442_58178# a_36442_57174# 1.00fF
C5482 a_9513_65301# VDD 1.37fF
C5483 vcm_commonmode a_47394_61190# 0.31fF
C5484 a_1770_14441# a_1923_59583# 1.17fF
C5485 a_42709_29199# m2_48260_24282# 0.60fF
C5486 a_43470_16520# a_43470_15516# 1.00fF
C5487 vcm_commonmode a_37446_24552# 0.84fF
C5488 vcm_commonmode a_19282_67214# 0.31fF
C5489 a_28410_19532# a_28410_18528# 1.00fF
C5490 a_2021_17973# a_3417_33231# 0.92fF
C5491 a_32334_10862# a_32426_10496# 0.32fF
C5492 a_48490_62194# ctopp 3.43fF
C5493 a_44474_70226# VDD 0.51fF
C5494 a_19374_68218# ctopp 3.59fF
C5495 vcm_commonmode a_47486_55166# 0.84fF
C5496 a_17507_52047# a_21382_64202# 0.38fF
C5497 a_12341_3311# a_22386_8488# 0.38fF
C5498 vcm_commonmode a_39454_57174# 0.87fF
C5499 a_27535_30503# a_34482_29941# 0.52fF
C5500 a_25398_16520# VDD 0.51fF
C5501 a_19788_48981# VDD 0.88fF
C5502 a_4482_57863# a_17039_51157# 0.65fF
C5503 a_47394_60186# a_47486_60186# 0.32fF
C5504 a_32951_27247# a_33430_21540# 0.38fF
C5505 a_49402_66210# VDD 0.31fF
C5506 a_18278_11866# a_18370_11500# 0.32fF
C5507 vcm_commonmode a_32334_16886# 0.31fF
C5508 a_8531_70543# a_25419_50959# 1.94fF
C5509 a_1586_21959# a_4417_22671# 0.54fF
C5510 a_1761_43567# a_13909_39747# 3.41fF
C5511 a_23390_72234# VDD 1.23fF
C5512 a_1761_52815# a_4887_36495# 0.37fF
C5513 a_21371_52263# a_12727_58255# 0.40fF
C5514 a_1768_16367# config_1_in[11] 1.19fF
C5515 a_23390_15516# a_23390_14512# 1.00fF
C5516 a_42374_18894# a_42466_18528# 0.32fF
C5517 a_13123_38231# a_1761_32143# 1.85fF
C5518 a_1591_18543# VDD 0.37fF
C5519 vcm_commonmode a_28410_72234# 0.69fF
C5520 a_31422_61190# a_32426_61190# 0.97fF
C5521 a_28756_7638# a_12546_22351# 0.41fF
C5522 a_33864_28111# a_34434_23548# 0.36fF
C5523 a_22294_24918# a_22386_24552# 0.32fF
C5524 a_15011_34717# VDD 1.92fF
C5525 a_1761_46287# a_13909_41923# 1.82fF
C5526 a_1803_20719# a_12663_40871# 2.78fF
C5527 a_2021_17973# a_30412_42589# 0.64fF
C5528 a_17366_7484# VDD 1.61fF
C5529 a_37446_68218# a_37446_67214# 1.00fF
C5530 a_8531_70543# a_4339_64521# 0.39fF
C5531 a_3983_48469# a_4149_48469# 0.72fF
C5532 vcm_commonmode a_24394_68218# 0.87fF
C5533 a_33430_58178# VDD 0.51fF
C5534 ctopn a_41967_31375# 2.62fF
C5535 a_2021_22325# a_5211_24759# 0.65fF
C5536 a_3339_43023# a_2143_15271# 2.67fF
C5537 a_8994_63927# VDD 0.72fF
C5538 a_18979_30287# a_25953_32143# 0.63fF
C5539 a_2411_26133# a_1591_36501# 0.34fF
C5540 a_19282_62194# a_19374_62194# 0.32fF
C5541 a_19374_56170# ctopp 3.39fF
C5542 a_6786_37557# VDD 0.58fF
C5543 a_8583_33551# a_12473_36341# 0.74fF
C5544 a_7775_10625# VDD 0.53fF
C5545 a_26417_40193# VDD 1.62fF
C5546 vcm_commonmode a_18278_64202# 0.31fF
C5547 a_22386_69222# a_22386_68218# 1.00fF
C5548 a_18151_52263# a_24394_65206# 0.38fF
C5549 a_1761_50639# a_7387_46831# 0.40fF
C5550 a_39222_48169# a_40458_72234# 0.35fF
C5551 a_42718_27497# a_12727_15529# 0.41fF
C5552 a_16746_60188# a_16362_60186# 2.28fF
C5553 a_34434_8488# a_35438_8488# 0.97fF
C5554 a_36797_27497# a_37446_22544# 0.38fF
C5555 a_31691_32143# VDD 0.57fF
C5556 a_1803_19087# a_14293_41807# 1.12fF
C5557 a_24302_57174# a_24394_57174# 0.32fF
C5558 vcm_commonmode VDD 621.65fF
C5559 a_27314_15882# a_27406_15516# 0.32fF
C5560 ctopn a_45478_21540# 3.59fF
C5561 a_28115_44535# VDD 0.59fF
C5562 a_39222_48169# a_40458_68218# 0.38fF
C5563 a_35438_70226# a_36442_70226# 0.97fF
C5564 a_12985_19087# a_12899_11471# 0.62fF
C5565 a_47486_19532# a_47486_18528# 1.00fF
C5566 a_7756_19087# VDD 0.53fF
C5567 a_6559_59663# a_11067_47695# 0.87fF
C5568 a_3325_18543# VDD 4.61fF
C5569 vcm_commonmode a_38450_13508# 0.87fF
C5570 a_18370_61190# ctopp 3.58fF
C5571 a_46482_59182# a_46482_58178# 1.00fF
C5572 ctopn a_22386_10496# 3.59fF
C5573 a_20378_69222# VDD 0.51fF
C5574 a_12621_44099# a_12381_43957# 3.40fF
C5575 a_23567_44211# a_1803_20719# 0.58fF
C5576 a_47486_9492# VDD 0.51fF
C5577 vcm_commonmode a_24394_56170# 0.87fF
C5578 a_16955_52047# a_20378_57174# 0.38fF
C5579 a_5943_15492# VDD 0.62fF
C5580 vcm_commonmode a_27314_69222# 0.31fF
C5581 a_21371_50959# a_25398_70226# 0.38fF
C5582 a_25306_71230# a_25398_71230# 0.32fF
C5583 a_33430_60186# a_33430_59182# 1.00fF
C5584 a_27406_22544# VDD 0.51fF
C5585 a_18370_65206# VDD 0.52fF
C5586 a_22386_63198# a_22386_62194# 1.00fF
C5587 a_37354_11866# a_37446_11500# 0.32fF
C5588 a_35959_30485# VDD 0.32fF
C5589 a_11067_66191# a_11067_21583# 1.45fF
C5590 a_18611_52047# a_13643_28327# 2.23fF
C5591 a_38557_32143# a_38450_60186# 0.38fF
C5592 a_1929_10651# a_3327_9308# 0.36fF
C5593 a_42466_15516# a_42466_14512# 1.00fF
C5594 vcm_commonmode a_34342_22910# 0.31fF
C5595 a_22386_70226# ctopp 3.58fF
C5596 a_39454_58178# ctopp 3.59fF
C5597 a_23395_52047# a_27406_66210# 0.38fF
C5598 a_41872_29423# a_10975_66407# 0.40fF
C5599 vcm_commonmode a_25306_65206# 0.31fF
C5600 ctopn a_33864_28111# 2.62fF
C5601 a_11067_21583# a_12895_13967# 0.57fF
C5602 a_16362_61190# VDD 2.48fF
C5603 a_27406_9492# a_27406_8488# 1.00fF
C5604 a_41370_24918# a_41462_24552# 0.32fF
C5605 a_19596_34215# VDD 1.22fF
C5606 ctopn a_17366_15516# 3.43fF
C5607 a_22386_67214# a_23390_67214# 0.97fF
C5608 vcm_commonmode a_23390_61190# 0.87fF
C5609 a_21371_52263# a_26402_62194# 0.38fF
C5610 a_39222_48169# a_40458_56170# 0.38fF
C5611 a_23390_14512# VDD 0.51fF
C5612 a_12895_13967# a_16746_18526# 0.41fF
C5613 a_19576_51701# a_20535_51727# 0.73fF
C5614 a_18278_55166# VDD 0.36fF
C5615 a_49494_64202# VDD 1.26fF
C5616 a_12869_2741# a_10515_23975# 2.15fF
C5617 a_38358_62194# a_38450_62194# 0.32fF
C5618 vcm_commonmode a_30326_14878# 0.31fF
C5619 ctopn a_27406_11500# 3.59fF
C5620 a_26748_7638# a_26402_24552# 0.46fF
C5621 a_32031_37683# VDD 2.45fF
C5622 a_1895_38842# VDD 1.24fF
C5623 a_5024_67885# a_7155_55509# 0.38fF
C5624 a_41462_69222# a_41462_68218# 1.00fF
C5625 a_13183_52047# a_12355_15055# 0.40fF
C5626 a_32134_49159# VDD 0.84fF
C5627 a_38557_32143# a_12901_66665# 0.40fF
C5628 vcm_commonmode a_27406_70226# 0.87fF
C5629 a_28410_23548# VDD 0.52fF
C5630 a_31422_8488# a_31422_7484# 1.00fF
C5631 a_25398_66210# VDD 0.51fF
C5632 a_13643_28327# a_28757_27247# 1.22fF
C5633 a_8123_56399# a_7050_53333# 0.45fF
C5634 a_25313_31599# VDD 1.07fF
C5635 a_1761_43567# a_33155_40191# 0.54fF
C5636 a_43378_57174# a_43470_57174# 0.32fF
C5637 a_46390_15882# a_46482_15516# 0.32fF
C5638 vcm_commonmode a_35346_23914# 0.31fF
C5639 a_3339_30503# a_6459_30511# 0.67fF
C5640 a_1775_47381# a_1941_47381# 0.75fF
C5641 a_3162_43023# VDD 0.64fF
C5642 vcm_commonmode a_32334_66210# 0.31fF
C5643 ctopn a_42709_29199# 2.49fF
C5644 a_24394_58178# a_25398_58178# 0.97fF
C5645 a_13123_38231# a_12663_35431# 3.79fF
C5646 a_37446_19532# VDD 0.51fF
C5647 a_8575_74853# a_10883_71855# 0.58fF
C5648 a_32951_27247# a_12877_16911# 0.41fF
C5649 a_8273_42479# a_9367_29397# 0.48fF
C5650 a_19374_9492# a_20378_9492# 0.97fF
C5651 a_20378_13508# a_20378_12504# 1.00fF
C5652 vcm_commonmode a_44382_19898# 0.31fF
C5653 a_28410_67214# ctopp 3.59fF
C5654 a_8583_33551# a_13357_32143# 0.33fF
C5655 a_35438_16520# a_36442_16520# 0.97fF
C5656 a_27393_47919# VDD 0.40fF
C5657 a_44382_71230# a_44474_71230# 0.32fF
C5658 a_6614_21237# VDD 0.46fF
C5659 vcm_commonmode a_45478_8488# 0.86fF
C5660 a_2411_26133# a_1761_37039# 1.04fF
C5661 a_41462_63198# a_41462_62194# 1.00fF
C5662 a_11803_29967# VDD 0.31fF
C5663 a_34780_56398# a_12901_58799# 0.40fF
C5664 vcm_commonmode a_16746_58180# 5.36fF
C5665 a_8197_31599# a_15207_30511# 0.47fF
C5666 a_29414_72234# m3_29316_72146# 2.80fF
C5667 a_6863_42692# a_6269_43567# 0.43fF
C5668 a_24740_7638# a_24394_8488# 0.38fF
C5669 ctopn a_9503_26151# 2.62fF
C5670 a_10543_16580# VDD 0.45fF
C5671 a_31330_72234# a_31422_72234# 0.32fF
C5672 a_39223_32463# a_39454_11500# 0.38fF
C5673 a_24740_7638# a_12877_14441# 0.41fF
C5674 a_3295_54421# a_3141_59887# 0.56fF
C5675 a_45386_24918# VDD 0.36fF
C5676 a_46482_9492# a_46482_8488# 1.00fF
C5677 a_11067_13095# a_2872_44111# 0.44fF
C5678 a_40675_27791# a_41462_22544# 0.38fF
C5679 a_17712_7638# a_17366_22544# 0.38fF
C5680 a_26748_7638# a_12985_7663# 0.41fF
C5681 a_17711_32385# VDD 0.32fF
C5682 a_46482_58178# a_46482_57174# 1.00fF
C5683 a_41462_67214# a_42466_67214# 0.97fF
C5684 a_27387_32373# a_27417_32509# 0.31fF
C5685 a_26514_47375# a_27393_47919# 0.64fF
C5686 vcm_commonmode a_33430_67214# 0.87fF
C5687 a_40458_20536# VDD 0.51fF
C5688 a_43175_28335# a_12877_16911# 0.41fF
C5689 a_29760_7638# a_12899_10927# 0.41fF
C5690 a_29414_63198# VDD 0.57fF
C5691 a_20635_29415# a_12899_2767# 0.62fF
C5692 a_2411_26133# a_1761_32143# 0.80fF
C5693 a_12349_25847# a_11865_24527# 0.31fF
C5694 a_30943_38695# a_30115_38695# 0.52fF
C5695 a_2847_36799# VDD 0.67fF
C5696 a_23298_13874# a_23390_13508# 0.32fF
C5697 vcm_commonmode a_47394_20902# 0.31fF
C5698 a_4443_46607# a_7464_39215# 0.42fF
C5699 a_1761_47919# a_14293_41807# 3.32fF
C5700 vcm_commonmode a_36350_63198# 0.31fF
C5701 a_36613_48169# a_12355_15055# 0.40fF
C5702 a_28318_68218# a_28410_68218# 0.32fF
C5703 a_33681_49373# VDD 0.35fF
C5704 a_21371_50959# a_12516_7093# 0.40fF
C5705 a_23390_59182# VDD 0.51fF
C5706 a_8583_33551# a_18979_30287# 0.95fF
C5707 a_6816_19355# VDD 3.73fF
C5708 a_27406_7484# a_28410_7484# 0.97fF
C5709 vcm_commonmode a_30418_9492# 0.87fF
C5710 m3_33332_72146# VDD 0.41fF
C5711 a_39454_24552# m3_39356_24414# 2.81fF
C5712 vcm_commonmode a_46482_16520# 0.87fF
C5713 a_27406_64202# ctopp 3.59fF
C5714 ctopn a_32426_13508# 3.59fF
C5715 a_34342_72234# VDD 0.61fF
C5716 vcm_commonmode a_30326_59182# 0.31fF
C5717 a_40458_12504# VDD 0.51fF
C5718 a_16891_43177# VDD 0.64fF
C5719 a_12139_18517# VDD 0.51fF
C5720 a_37459_51183# VDD 0.66fF
C5721 a_2775_46025# a_2099_59861# 2.68fF
C5722 a_38450_9492# a_39454_9492# 0.97fF
C5723 vcm_commonmode a_47394_12870# 0.31fF
C5724 a_21382_64202# a_22386_64202# 0.97fF
C5725 a_39454_13508# a_39454_12504# 1.00fF
C5726 a_40050_48463# a_45478_63198# 0.42fF
C5727 a_28524_47919# a_26417_47919# 0.50fF
C5728 a_31768_55394# a_31422_69222# 0.38fF
C5729 a_10515_22671# a_7571_26151# 0.42fF
C5730 a_35438_21540# VDD 0.51fF
C5731 vcm_commonmode a_38450_7484# 0.69fF
C5732 a_18370_22544# a_19374_22544# 0.97fF
C5733 a_12907_27023# a_26523_29199# 0.40fF
C5734 a_17415_29423# VDD 0.30fF
C5735 vcm_commonmode a_42374_21906# 0.31fF
C5736 a_36442_69222# ctopp 3.59fF
C5737 a_5449_25071# a_6649_25615# 0.37fF
C5738 vcm_commonmode a_32426_64202# 0.87fF
C5739 a_40458_17524# VDD 0.51fF
C5740 a_1591_49557# VDD 0.45fF
C5741 a_27406_60186# VDD 0.51fF
C5742 vcm_commonmode a_19282_10862# 0.31fF
C5743 vcm_commonmode a_47394_17890# 0.31fF
C5744 a_34434_65206# ctopp 3.59fF
C5745 a_12641_43124# a_15193_41781# 0.66fF
C5746 a_2971_73493# VDD 0.55fF
C5747 vcm_commonmode a_34342_60186# 0.31fF
C5748 a_29414_67214# a_29414_66210# 1.00fF
C5749 a_1761_43567# VDD 8.85fF
C5750 a_10409_18543# VDD 0.62fF
C5751 a_43270_27791# a_12877_16911# 0.41fF
C5752 a_5963_20149# a_5825_20495# 0.52fF
C5753 a_1761_40847# a_13005_35823# 6.83fF
C5754 a_12641_37684# a_12343_36893# 0.37fF
C5755 a_43362_28879# a_20267_30503# 0.92fF
C5756 a_25398_65206# a_25398_64202# 1.00fF
C5757 a_42374_13874# a_42466_13508# 0.32fF
C5758 vcm_commonmode a_20378_19532# 0.87fF
C5759 a_25971_52263# a_30418_55166# 0.46fF
C5760 a_2021_17973# a_12381_43957# 1.22fF
C5761 a_47394_68218# a_47486_68218# 0.32fF
C5762 vcm_commonmode a_24740_7638# 10.35fF
C5763 a_36717_47375# a_12257_56623# 0.40fF
C5764 vcm_commonmode a_41462_69222# 0.87fF
C5765 a_4482_57863# a_30928_49007# 0.71fF
C5766 a_3295_54421# a_4891_47388# 0.36fF
C5767 a_46482_7484# a_47486_7484# 0.97fF
C5768 a_2952_53333# a_5541_53609# 0.64fF
C5769 a_19374_23548# a_19374_22544# 1.00fF
C5770 ctopp a_33430_55166# 1.70fF
C5771 a_28318_56170# a_28410_56170# 0.32fF
C5772 a_31768_55394# a_10515_22671# 0.40fF
C5773 vcm_commonmode a_48490_22544# 0.87fF
C5774 a_17366_11500# VDD 0.58fF
C5775 a_30418_69222# a_31422_69222# 0.97fF
C5776 vcm_commonmode a_39454_65206# 0.87fF
C5777 a_41462_18528# VDD 0.51fF
C5778 a_17599_52263# a_18611_52047# 0.33fF
C5779 a_29760_7638# a_29414_16520# 0.38fF
C5780 a_25398_61190# a_25398_60186# 1.00fF
C5781 a_21382_24552# VDD 0.60fF
C5782 vcm_commonmode a_24302_11866# 0.31fF
C5783 ctopn a_39454_8488# 3.40fF
C5784 a_40458_64202# a_41462_64202# 0.97fF
C5785 vcm_commonmode a_48398_18894# 0.31fF
C5786 a_41462_66210# ctopp 3.59fF
C5787 vcm_commonmode a_28318_24918# 0.31fF
C5788 a_2007_45717# VDD 0.48fF
C5789 a_11803_55311# a_12901_66959# 1.08fF
C5790 a_16746_20534# VDD 33.20fF
C5791 a_32334_55166# VDD 0.36fF
C5792 a_4758_45369# a_19946_51157# 0.55fF
C5793 a_37446_22544# a_38450_22544# 0.97fF
C5794 a_23390_57174# VDD 0.51fF
C5795 vcm_commonmode a_44474_14512# 0.87fF
C5796 a_40491_27247# a_42718_27497# 1.28fF
C5797 a_28410_65206# a_29414_65206# 0.97fF
C5798 vcm_commonmode a_23390_20536# 0.87fF
C5799 vcm_commonmode a_38358_55166# 0.30fF
C5800 a_16746_68220# a_16362_68218# 2.28fF
C5801 a_24394_17524# a_24394_16520# 1.00fF
C5802 vcm_commonmode a_30326_57174# 0.31fF
C5803 a_20359_29199# a_13643_28327# 1.67fF
C5804 a_16362_16520# VDD 2.47fF
C5805 a_4240_48981# VDD 0.69fF
C5806 a_19374_23548# a_20378_23548# 0.97fF
C5807 a_9955_20969# a_7377_18012# 0.52fF
C5808 VDD dummypin[11] 0.85fF
C5809 a_28410_56170# a_28410_55166# 1.00fF
C5810 a_2004_42453# config_2_in[3] 0.77fF
C5811 a_19720_55394# a_12727_58255# 0.40fF
C5812 a_48490_67214# a_48490_66210# 1.00fF
C5813 vcm_commonmode a_49494_23548# 0.90fF
C5814 a_6727_47607# a_4674_40277# 0.36fF
C5815 a_4563_32900# a_5831_39189# 1.45fF
C5816 a_16746_12502# VDD 33.20fF
C5817 a_23567_43123# VDD 2.06fF
C5818 a_43362_28879# a_12983_63151# 0.40fF
C5819 vcm_commonmode a_46482_66210# 0.87fF
C5820 a_1591_69141# a_1757_69141# 0.72fF
C5821 a_11067_47695# a_10791_15529# 0.37fF
C5822 a_25133_37571# a_31847_36893# 1.06fF
C5823 vcm_commonmode a_21382_72234# 0.69fF
C5824 a_37446_62194# VDD 0.51fF
C5825 a_27314_61190# a_27406_61190# 0.32fF
C5826 vcm_commonmode a_23390_12504# 0.87fF
C5827 ctopn a_24394_9492# 3.58fF
C5828 a_43269_29967# a_12985_7663# 0.41fF
C5829 a_44474_65206# a_44474_64202# 1.00fF
C5830 a_1591_12565# a_1757_12565# 0.75fF
C5831 ctopn a_40458_16520# 3.59fF
C5832 vcm_commonmode a_44382_62194# 0.31fF
C5833 a_45478_15516# VDD 0.51fF
C5834 a_7295_44647# VDD 9.93fF
C5835 a_12901_66665# a_16746_70228# 2.28fF
C5836 a_28410_19532# a_29414_19532# 0.97fF
C5837 a_1683_52271# a_1849_52271# 0.57fF
C5838 a_9135_27239# a_12895_13967# 0.41fF
C5839 a_38450_23548# a_38450_22544# 1.00fF
C5840 a_10680_52245# a_6775_53877# 0.44fF
C5841 a_45478_63198# ctopp 3.64fF
C5842 a_47394_56170# a_47486_56170# 0.32fF
C5843 a_43470_71230# VDD 0.58fF
C5844 a_32426_66210# a_32426_65206# 1.00fF
C5845 a_33430_14512# a_34434_14512# 0.97fF
C5846 vcm_commonmode a_18370_21540# 0.88fF
C5847 a_34759_31029# a_32823_29397# 0.36fF
C5848 a_7847_40847# VDD 0.57fF
C5849 a_16955_52047# a_20378_65206# 0.38fF
C5850 a_12899_11471# VDD 8.07fF
C5851 a_44474_61190# a_44474_60186# 1.00fF
C5852 a_11574_22869# VDD 1.27fF
C5853 a_30326_8854# a_30418_8488# 0.32fF
C5854 a_39454_59182# ctopp 3.59fF
C5855 ctopp m3_17268_56082# 0.46fF
C5856 a_27195_32375# VDD 0.57fF
C5857 vcm_commonmode a_23390_17524# 0.87fF
C5858 a_22386_13508# VDD 0.51fF
C5859 a_31330_70226# a_31422_70226# 0.32fF
C5860 a_36717_47375# a_36442_68218# 0.38fF
C5861 a_30418_62194# a_30418_61190# 1.00fF
C5862 a_21382_10496# a_21382_9492# 1.00fF
C5863 vcm_commonmode a_29322_13874# 0.31fF
C5864 a_2099_59861# a_4427_25071# 1.15fF
C5865 a_47486_65206# a_48490_65206# 0.97fF
C5866 a_19743_36919# VDD 0.62fF
C5867 a_2952_46805# a_2004_42453# 0.39fF
C5868 a_1761_44111# a_13716_43047# 3.55fF
C5869 a_1761_22895# a_12381_43957# 0.49fF
C5870 a_43470_17524# a_43470_16520# 1.00fF
C5871 ctopn a_12947_23413# 1.43fF
C5872 a_16510_8760# a_11067_23759# 9.01fF
C5873 a_27535_30503# a_24959_30503# 0.32fF
C5874 a_10195_48437# VDD 0.43fF
C5875 a_17507_52047# a_21382_70226# 0.38fF
C5876 a_30418_20536# a_30418_19532# 1.00fF
C5877 a_38450_23548# a_39454_23548# 0.97fF
C5878 a_40050_48463# VDD 7.22fF
C5879 a_35438_66210# a_36442_66210# 0.97fF
C5880 a_34780_56398# a_34434_60186# 0.38fF
C5881 vcm_commonmode a_44474_59182# 0.87fF
C5882 a_8531_70543# a_2959_47113# 1.55fF
C5883 a_3607_34639# a_6162_28487# 0.72fF
C5884 a_28757_27247# a_30790_30663# 0.34fF
C5885 a_4674_40277# a_17311_46833# 0.37fF
C5886 a_36717_47375# a_10975_66407# 0.40fF
C5887 a_18611_52047# a_23390_66210# 0.38fF
C5888 a_38115_52263# a_16863_29415# 0.42fF
C5889 a_12341_3311# a_12877_16911# 0.41fF
C5890 a_46390_61190# a_46482_61190# 0.32fF
C5891 a_43470_60186# ctopp 3.59fF
C5892 a_46482_68218# VDD 0.51fF
C5893 a_12970_34191# VDD 0.36fF
C5894 vcm_commonmode a_24394_18528# 0.87fF
C5895 a_46390_7850# VDD 0.62fF
C5896 a_17599_52263# a_22386_62194# 0.38fF
C5897 a_18278_67214# a_18370_67214# 0.32fF
C5898 a_36717_47375# a_36442_56170# 0.38fF
C5899 ctopn a_42466_22544# 3.58fF
C5900 a_2952_66139# a_3143_66972# 0.46fF
C5901 a_35438_71230# a_35438_70226# 1.00fF
C5902 a_5682_69367# a_4351_67279# 1.23fF
C5903 a_47486_19532# a_48490_19532# 0.97fF
C5904 a_8123_56399# a_14831_50095# 1.44fF
C5905 a_19889_27497# a_22026_27497# 0.73fF
C5906 a_10975_55535# a_11141_55535# 0.65fF
C5907 a_10865_69679# VDD 0.67fF
C5908 vcm_commonmode a_17274_55166# 0.30fF
C5909 a_10506_29967# a_13390_29575# 0.40fF
C5910 a_33856_40743# VDD 1.76fF
C5911 a_5160_68315# a_5167_68060# 0.42fF
C5912 a_2952_66139# a_1823_65853# 0.79fF
C5913 a_11067_46823# VDD 19.01fF
C5914 vcm_commonmode a_18278_70226# 0.31fF
C5915 a_31768_55394# a_12901_66665# 0.40fF
C5916 a_31422_20536# a_32426_20536# 0.97fF
C5917 a_7210_55081# a_8491_57487# 0.62fF
C5918 a_49402_8854# a_49494_8488# 0.32fF
C5919 vcm_commonmode a_33430_10496# 0.87fF
C5920 a_12355_65103# VDD 14.59fF
C5921 a_8132_53511# a_9240_53877# 0.41fF
C5922 a_20378_63198# a_21382_63198# 0.97fF
C5923 ctopn a_38450_14512# 3.59fF
C5924 a_7615_73193# VDD 0.44fF
C5925 vcm_commonmode a_48490_60186# 0.87fF
C5926 a_2873_13879# a_3843_13880# 0.33fF
C5927 a_21382_71230# ctopp 3.40fF
C5928 ctopn a_17366_20536# 3.43fF
C5929 a_7571_26151# a_10407_47607# 0.35fF
C5930 a_13067_38517# VDD 8.43fF
C5931 a_20286_58178# a_20378_58178# 0.32fF
C5932 a_28756_7638# a_12985_16367# 0.41fF
C5933 a_49494_62194# a_49494_61190# 1.00fF
C5934 a_40458_10496# a_40458_9492# 1.00fF
C5935 a_46482_56170# VDD 0.52fF
C5936 vcm_commonmode a_43470_58178# 0.87fF
C5937 a_49402_69222# VDD 0.31fF
C5938 ctopn a_12727_13353# 3.23fF
C5939 a_29414_8488# VDD 0.58fF
C5940 vcm_commonmode a_20378_62194# 0.87fF
C5941 a_31330_16886# a_31422_16520# 0.32fF
C5942 ctopn a_43470_23548# 3.40fF
C5943 a_11067_46823# a_26514_47375# 0.51fF
C5944 a_49494_20536# a_49494_19532# 1.00fF
C5945 vcm_commonmode a_36350_8854# 0.31fF
C5946 ctopp a_47486_55166# 0.30fF
C5947 a_3016_60949# a_3295_62083# 0.63fF
C5948 vcm_commonmode a_28410_15516# 0.87fF
C5949 ctopn a_17366_12504# 3.43fF
C5950 a_39454_57174# ctopp 3.58fF
C5951 a_23395_52047# a_12901_58799# 0.40fF
C5952 a_9503_26151# a_20378_9492# 0.38fF
C5953 a_27535_30503# a_22843_29415# 1.62fF
C5954 vcm_commonmode a_26402_71230# 0.86fF
C5955 a_29414_21540# a_29414_20536# 1.00fF
C5956 a_45478_61190# VDD 0.51fF
C5957 vcm_commonmode a_38450_11500# 0.87fF
C5958 a_36629_27791# a_36442_22544# 0.38fF
C5959 a_17366_67214# VDD 0.57fF
C5960 a_31422_12504# a_32426_12504# 0.97fF
C5961 a_32167_29611# a_12899_3855# 0.50fF
C5962 a_3024_67191# a_6095_44807# 0.55fF
C5963 a_2689_65103# a_6831_63303# 0.33fF
C5964 a_37354_67214# a_37446_67214# 0.32fF
C5965 a_12877_16911# a_16746_13506# 2.28fF
C5966 vcm_commonmode a_42466_24552# 0.84fF
C5967 a_16863_29415# a_20267_30503# 0.48fF
C5968 a_34482_29941# a_7295_44647# 2.37fF
C5969 vcm_commonmode a_24302_67214# 0.31fF
C5970 a_16863_29415# a_28963_28853# 0.75fF
C5971 a_49494_70226# VDD 1.10fF
C5972 a_7155_55509# a_7210_55081# 0.39fF
C5973 a_24394_68218# ctopp 3.59fF
C5974 ctopn a_17366_17524# 3.43fF
C5975 a_1761_46287# a_12357_37999# 0.82fF
C5976 a_25971_52263# a_12355_15055# 0.40fF
C5977 a_2411_18517# a_10995_14333# 0.32fF
C5978 a_2292_17179# a_2830_15431# 0.51fF
C5979 vcm_commonmode a_44474_57174# 0.87fF
C5980 ctopn a_10515_23975# 2.99fF
C5981 a_30418_16520# VDD 0.51fF
C5982 a_23847_47919# VDD 0.49fF
C5983 a_14287_51175# a_12516_7093# 0.49fF
C5984 a_33864_28111# a_34434_14512# 0.38fF
C5985 a_5612_58229# VDD 0.42fF
C5986 a_23298_7850# a_23390_7484# 0.32fF
C5987 vcm_commonmode a_21290_9858# 0.31fF
C5988 a_32426_24552# m3_32328_24414# 2.09fF
C5989 a_39454_63198# a_40458_63198# 0.97fF
C5990 a_21273_30485# VDD 0.75fF
C5991 vcm_commonmode a_37354_16886# 0.31fF
C5992 a_4351_67279# a_4215_51157# 0.89fF
C5993 a_15193_41781# a_15459_41781# 0.33fF
C5994 a_27314_72234# VDD 0.61fF
C5995 a_1761_52815# a_13669_37429# 0.51fF
C5996 a_17039_51157# a_22015_50645# 0.34fF
C5997 a_22164_51157# VDD 0.38fF
C5998 a_26402_21540# a_27406_21540# 0.97fF
C5999 a_34342_9858# a_34434_9492# 0.32fF
C6000 ctopp VDD 94.33fF
C6001 a_1768_13103# config_2_in[9] 1.60fF
C6002 a_11619_56615# a_11067_46823# 0.30fF
C6003 a_17274_64202# a_17366_64202# 0.32fF
C6004 a_22386_7484# VDD 1.40fF
C6005 a_44474_58178# a_45478_58178# 0.97fF
C6006 a_11619_56615# a_12355_65103# 3.76fF
C6007 a_41427_52263# a_41462_63198# 0.42fF
C6008 a_18500_47491# VDD 0.50fF
C6009 a_23395_52047# a_27406_69222# 0.38fF
C6010 vcm_commonmode a_29414_68218# 0.87fF
C6011 a_42718_27497# a_44474_13508# 0.38fF
C6012 a_33430_59182# a_34434_59182# 0.97fF
C6013 a_35601_27497# a_12985_19087# 0.41fF
C6014 a_32951_27247# a_12895_13967# 0.41fF
C6015 a_16746_64204# VDD 33.21fF
C6016 a_18979_30287# a_30052_32117# 0.31fF
C6017 a_4095_29423# VDD 0.39fF
C6018 a_23736_7638# a_23390_22544# 0.38fF
C6019 a_12473_41781# a_13909_39747# 0.57fF
C6020 a_24394_56170# ctopp 3.40fF
C6021 a_1761_50639# a_13669_37429# 2.08fF
C6022 a_12907_56399# a_10515_22671# 0.51fF
C6023 ctopn a_18370_18528# 3.58fF
C6024 a_5039_42167# a_5098_41641# 0.48fF
C6025 vcm_commonmode a_23298_64202# 0.31fF
C6026 a_31422_17524# a_32426_17524# 0.97fF
C6027 a_2099_59861# a_2292_43291# 0.42fF
C6028 a_48490_21540# a_48490_20536# 1.00fF
C6029 a_18370_60186# a_19374_60186# 0.97fF
C6030 a_1923_54591# a_4555_55233# 0.33fF
C6031 a_35438_24552# a_35438_23548# 1.00fF
C6032 a_20378_12504# a_20378_11500# 1.00fF
C6033 a_2787_30503# a_20881_28111# 1.62fF
C6034 a_15607_46805# a_18979_30287# 1.29fF
C6035 a_1761_47919# a_1941_47381# 0.59fF
C6036 a_38454_43983# VDD 0.81fF
C6037 a_24740_7638# a_12899_11471# 0.41fF
C6038 a_7078_36103# a_6883_37019# 0.42fF
C6039 a_15439_49525# a_11251_59879# 3.62fF
C6040 vcm_commonmode a_43470_13508# 0.87fF
C6041 a_23390_61190# ctopp 3.59fF
C6042 ctopn a_27406_10496# 3.59fF
C6043 a_25398_69222# VDD 0.51fF
C6044 a_7019_35951# VDD 0.48fF
C6045 a_21371_52263# a_26402_55166# 0.46fF
C6046 a_11067_23759# a_25744_7638# 1.41fF
C6047 a_9963_29967# a_10045_29967# 0.30fF
C6048 a_29760_55394# a_12257_56623# 0.40fF
C6049 vcm_commonmode a_29414_56170# 0.87fF
C6050 a_2235_30503# a_7862_34025# 0.92fF
C6051 a_11067_46823# a_34482_29941# 1.42fF
C6052 vcm_commonmode a_32334_69222# 0.31fF
C6053 a_2339_38129# a_1586_21959# 1.70fF
C6054 a_3339_43023# a_1761_46287# 2.67fF
C6055 a_32426_22544# VDD 0.51fF
C6056 a_42374_7850# a_42466_7484# 0.32fF
C6057 a_4758_45369# a_10680_54171# 0.36fF
C6058 a_43175_28335# a_12895_13967# 0.41fF
C6059 a_42709_29199# a_48490_19532# 0.38fF
C6060 a_23390_65206# VDD 0.51fF
C6061 a_29927_29199# a_30155_32375# 0.39fF
C6062 a_18151_52263# a_10515_22671# 0.55fF
C6063 vcm_commonmode a_39362_22910# 0.31fF
C6064 a_27406_70226# ctopp 3.58fF
C6065 a_16362_72234# m3_16264_72146# 2.81fF
C6066 a_5483_11140# VDD 0.42fF
C6067 a_26310_69222# a_26402_69222# 0.32fF
C6068 vcm_commonmode a_30326_65206# 0.31fF
C6069 a_32426_18528# a_32426_17524# 1.00fF
C6070 a_30762_49641# VDD 0.55fF
C6071 a_18370_72234# a_19374_72234# 0.97fF
C6072 a_45478_21540# a_46482_21540# 0.97fF
C6073 a_36797_27497# a_12727_13353# 0.41fF
C6074 a_8031_24527# VDD 0.37fF
C6075 a_36350_64202# a_36442_64202# 0.32fF
C6076 ctopn a_22386_15516# 3.59fF
C6077 a_13143_29575# a_9731_22895# 0.47fF
C6078 vcm_commonmode a_28410_61190# 0.87fF
C6079 a_14354_32117# a_14298_32143# 0.75fF
C6080 a_28410_14512# VDD 0.51fF
C6081 a_1586_66567# a_4351_67279# 0.76fF
C6082 a_23298_55166# VDD 0.35fF
C6083 a_19720_7638# a_12899_10927# 0.41fF
C6084 a_33338_22910# a_33430_22544# 0.32fF
C6085 a_22386_10496# a_23390_10496# 0.97fF
C6086 vcm_commonmode a_35346_14878# 0.31fF
C6087 ctopn a_32426_11500# 3.59fF
C6088 a_29760_7638# a_30764_7638# 0.41fF
C6089 a_24302_65206# a_24394_65206# 0.32fF
C6090 a_33430_14512# a_33430_13508# 1.00fF
C6091 a_42283_38007# VDD 0.68fF
C6092 a_12283_40183# VDD 0.65fF
C6093 a_11495_16341# VDD 0.54fF
C6094 vcm_commonmode a_32426_70226# 0.87fF
C6095 a_39223_32463# a_39454_10496# 0.38fF
C6096 a_37446_60186# a_38450_60186# 0.97fF
C6097 a_33430_23548# VDD 0.52fF
C6098 a_16746_58180# ctopp 1.68fF
C6099 a_43269_29967# a_47486_19532# 0.38fF
C6100 a_30418_66210# VDD 0.51fF
C6101 a_39454_12504# a_39454_11500# 1.00fF
C6102 a_21371_50959# a_34579_50613# 0.38fF
C6103 vcm_commonmode a_40366_23914# 0.31fF
C6104 a_8117_30287# a_8197_31599# 0.34fF
C6105 a_8383_43255# VDD 0.50fF
C6106 a_26402_70226# a_26402_69222# 1.00fF
C6107 a_39222_48169# a_12983_63151# 0.40fF
C6108 vcm_commonmode a_37354_66210# 0.31fF
C6109 a_32426_18528# a_33430_18528# 0.97fF
C6110 a_1591_36501# a_1757_36501# 0.72fF
C6111 a_42466_19532# VDD 0.51fF
C6112 a_10055_58791# a_17712_7638# 0.40fF
C6113 a_36797_27497# a_10515_23975# 0.41fF
C6114 a_12641_37684# a_1799_29556# 0.99fF
C6115 a_3024_67191# VDD 5.70fF
C6116 a_4339_64521# a_8994_63927# 0.31fF
C6117 vcm_commonmode a_49402_19898# 0.31fF
C6118 a_33430_67214# ctopp 3.59fF
C6119 a_49494_70226# m3_49396_70138# 2.78fF
C6120 a_41261_28335# a_12981_62313# 0.40fF
C6121 a_11803_55311# a_6835_46823# 0.64fF
C6122 a_24302_19898# a_24394_19532# 0.32fF
C6123 a_43270_27791# a_12895_13967# 0.41fF
C6124 a_15439_49525# a_2775_46025# 0.78fF
C6125 a_25398_11500# a_25398_10496# 1.00fF
C6126 vcm_commonmode a_21382_58178# 0.87fF
C6127 a_38315_39141# VDD 1.03fF
C6128 a_29322_14878# a_29414_14512# 0.32fF
C6129 a_12935_31287# a_12999_29423# 0.39fF
C6130 a_32426_72234# m3_32328_72146# 2.80fF
C6131 a_37951_42089# VDD 0.59fF
C6132 a_45386_69222# a_45478_69222# 0.32fF
C6133 a_11067_67279# a_7598_36103# 1.76fF
C6134 a_2283_15797# VDD 1.83fF
C6135 a_25787_28327# a_33430_72234# 0.34fF
C6136 a_6607_42167# a_5441_27791# 1.04fF
C6137 a_23390_55166# a_24394_55166# 0.97fF
C6138 a_9765_32143# VDD 0.95fF
C6139 a_28547_51175# a_35568_49525# 0.87fF
C6140 a_15959_42943# a_15193_42917# 0.32fF
C6141 a_2787_32679# a_4685_37583# 0.51fF
C6142 a_12257_56623# a_16746_57176# 0.41fF
C6143 a_17366_15516# a_18370_15516# 0.97fF
C6144 a_2292_43291# a_1761_25071# 0.43fF
C6145 vcm_commonmode a_38450_67214# 0.87fF
C6146 a_1823_72381# a_1770_14441# 0.71fF
C6147 a_39299_48783# a_12727_67753# 0.40fF
C6148 a_28547_51175# a_32426_68218# 0.38fF
C6149 a_1923_54591# a_2163_57853# 0.31fF
C6150 a_45478_20536# VDD 0.51fF
C6151 a_40491_27247# a_12899_10927# 0.41fF
C6152 a_34434_63198# VDD 0.57fF
C6153 a_41462_10496# a_42466_10496# 0.97fF
C6154 a_12663_39783# a_1761_39215# 0.55fF
C6155 a_2672_69513# VDD 0.30fF
C6156 a_43378_65206# a_43470_65206# 0.32fF
C6157 a_11067_13095# a_11943_63125# 0.41fF
C6158 a_28757_27247# a_28756_7638# 0.42fF
C6159 vcm_commonmode a_41370_63198# 0.31fF
C6160 a_42718_27497# a_44474_7484# 0.35fF
C6161 a_29760_55394# a_8531_70543# 0.34fF
C6162 a_43362_28879# a_47486_71230# 0.38fF
C6163 a_18611_52047# a_4351_67279# 0.46fF
C6164 a_12907_56399# a_12901_66665# 0.36fF
C6165 a_28410_59182# VDD 0.51fF
C6166 vcm_commonmode a_35438_9492# 0.87fF
C6167 a_34342_23914# a_34434_23548# 0.32fF
C6168 a_27406_11500# a_28410_11500# 0.97fF
C6169 a_39035_31055# VDD 0.31fF
C6170 a_32426_64202# ctopp 3.59fF
C6171 ctopn a_37446_13508# 3.59fF
C6172 a_38557_32143# VDD 8.85fF
C6173 a_31330_66210# a_31422_66210# 0.32fF
C6174 a_25971_52263# a_30418_60186# 0.38fF
C6175 vcm_commonmode a_35346_59182# 0.31fF
C6176 vcm_commonmode m3_16264_62106# 3.21fF
C6177 a_45478_12504# VDD 0.51fF
C6178 a_19720_55394# a_19374_66210# 0.38fF
C6179 a_45478_70226# a_45478_69222# 1.00fF
C6180 a_43267_31055# a_46482_67214# 0.38fF
C6181 a_29760_55394# a_10975_66407# 0.40fF
C6182 a_25517_37455# a_1761_31055# 4.44fF
C6183 a_30757_37455# a_31223_36369# 0.32fF
C6184 a_11067_47695# a_21261_47919# 0.59fF
C6185 a_3307_18259# VDD 0.51fF
C6186 vcm_commonmode a_41872_29423# 10.07fF
C6187 a_8039_61493# VDD 0.36fF
C6188 a_9955_20969# VDD 2.32fF
C6189 a_31422_24552# a_32426_24552# 0.97fF
C6190 a_16244_34973# VDD 1.47fF
C6191 a_14287_51175# a_18370_62194# 0.38fF
C6192 a_28547_51175# a_32426_56170# 0.36fF
C6193 a_43267_31055# a_12901_66959# 0.40fF
C6194 a_43378_19898# a_43470_19532# 0.32fF
C6195 a_40458_21540# VDD 0.51fF
C6196 vcm_commonmode a_43470_7484# 0.69fF
C6197 a_12889_39889# a_16043_38825# 0.54fF
C6198 a_3987_19623# a_5346_33775# 0.56fF
C6199 a_19807_28111# a_27016_29587# 0.33fF
C6200 a_28410_62194# a_29414_62194# 0.97fF
C6201 a_44474_11500# a_44474_10496# 1.00fF
C6202 a_4758_45369# a_12659_54965# 2.08fF
C6203 a_48398_14878# a_48490_14512# 0.32fF
C6204 vcm_commonmode a_47394_21906# 0.31fF
C6205 a_41462_69222# ctopp 3.59fF
C6206 a_17366_10496# VDD 0.57fF
C6207 a_16615_41001# VDD 0.65fF
C6208 a_1591_57711# a_1768_16367# 1.66fF
C6209 vcm_commonmode a_37446_64202# 0.87fF
C6210 a_12549_35836# a_15011_34717# 1.11fF
C6211 a_2011_34837# a_3607_34639# 0.37fF
C6212 a_45478_17524# VDD 0.51fF
C6213 a_6559_49557# VDD 0.50fF
C6214 a_18151_52263# a_12901_66665# 0.40fF
C6215 a_43362_28879# a_42985_46831# 5.63fF
C6216 a_27314_20902# a_27406_20536# 0.32fF
C6217 a_32426_60186# VDD 0.51fF
C6218 a_41462_55166# a_42466_55166# 0.97fF
C6219 vcm_commonmode a_24302_10862# 0.31fF
C6220 a_7773_63927# a_9424_60949# 0.33fF
C6221 a_15439_49525# a_12981_62313# 23.42fF
C6222 a_16746_63200# a_16362_63198# 2.28fF
C6223 a_9405_31599# VDD 0.56fF
C6224 a_39454_65206# ctopp 3.59fF
C6225 a_33430_57174# a_34434_57174# 0.97fF
C6226 a_3751_72373# VDD 2.46fF
C6227 vcm_commonmode a_39362_60186# 0.31fF
C6228 a_36442_15516# a_37446_15516# 0.97fF
C6229 vcm_commonmode a_16362_23548# 4.45fF
C6230 a_12907_56399# a_10680_52245# 2.89fF
C6231 a_6269_43567# VDD 0.53fF
C6232 a_1768_16367# a_1803_20719# 3.17fF
C6233 a_1768_16367# a_2007_51701# 0.59fF
C6234 a_14963_39783# a_14293_39631# 1.92fF
C6235 a_7948_38377# a_7187_37583# 0.38fF
C6236 a_28441_36389# VDD 1.65fF
C6237 vcm_commonmode a_25398_19532# 0.87fF
C6238 a_28547_51175# a_32426_55166# 0.42fF
C6239 a_12727_67753# a_16746_67216# 2.28fF
C6240 a_19788_48981# a_20161_48463# 0.62fF
C6241 vcm_commonmode a_46482_69222# 0.87fF
C6242 a_34434_71230# a_35438_71230# 0.97fF
C6243 a_49494_60186# m3_49396_60098# 2.78fF
C6244 a_31898_30761# VDD 0.34fF
C6245 a_46482_11500# a_47486_11500# 0.97fF
C6246 vcm_commonmode a_19282_15882# 0.31fF
C6247 a_20027_27221# a_17712_7638# 0.34fF
C6248 a_1761_41935# a_30943_38695# 0.45fF
C6249 a_16955_52047# a_12901_58799# 0.40fF
C6250 a_28446_31375# a_30790_30663# 0.79fF
C6251 vcm_commonmode m3_16264_9354# 3.20fF
C6252 a_22386_11500# VDD 0.51fF
C6253 a_12473_41781# VDD 6.84fF
C6254 vcm_commonmode a_44474_65206# 0.87fF
C6255 a_46482_18528# VDD 0.51fF
C6256 vcm_commonmode a_17274_71230# 0.33fF
C6257 a_24302_72234# a_24394_72234# 0.32fF
C6258 a_32951_27247# a_33430_16520# 0.38fF
C6259 a_26402_24552# VDD 0.60fF
C6260 vcm_commonmode a_29322_11866# 0.31fF
C6261 ctopn a_44474_8488# 3.40fF
C6262 a_27314_12870# a_27406_12504# 0.32fF
C6263 a_46482_66210# ctopp 3.59fF
C6264 a_1689_10396# a_1887_10422# 0.31fF
C6265 a_49494_55166# m2_48260_54946# 0.60fF
C6266 a_43269_29967# a_42709_29199# 3.15fF
C6267 a_12249_43457# a_12343_42333# 0.71fF
C6268 vcm_commonmode a_33338_24918# 0.31fF
C6269 a_2235_30503# a_7460_31055# 0.65fF
C6270 a_8308_44111# VDD 0.63fF
C6271 a_22386_59182# a_22386_58178# 1.00fF
C6272 a_30573_52271# a_30663_51727# 0.50fF
C6273 a_36442_55166# VDD 0.60fF
C6274 a_12341_3311# a_12895_13967# 0.41fF
C6275 a_10515_63143# VDD 13.81fF
C6276 a_47486_62194# a_48490_62194# 0.97fF
C6277 a_7773_63927# a_8199_58229# 1.32fF
C6278 a_28410_57174# VDD 0.51fF
C6279 vcm_commonmode a_49494_14512# 0.90fF
C6280 a_75794_40594# a_76346_40594# 0.72fF
C6281 a_48490_23548# m2_48260_24282# 0.98fF
C6282 vcm_commonmode a_28410_20536# 0.87fF
C6283 a_11067_67279# a_9751_25071# 0.36fF
C6284 vcm_commonmode a_43378_55166# 0.30fF
C6285 a_18611_52047# a_12355_15055# 0.45fF
C6286 a_18370_68218# a_19374_68218# 0.97fF
C6287 vcm_commonmode a_17366_63198# 1.88fF
C6288 vcm_commonmode a_35346_57174# 0.31fF
C6289 a_14831_50095# a_23019_48463# 0.33fF
C6290 a_4119_70741# a_2689_65103# 0.32fF
C6291 a_46390_20902# a_46482_20536# 0.32fF
C6292 a_11019_59575# VDD 0.71fF
C6293 a_25398_24552# m3_25300_24414# 2.81fF
C6294 a_35346_63198# a_35438_63198# 0.32fF
C6295 a_14097_31375# VDD 1.21fF
C6296 a_12473_42869# a_25221_41281# 0.30fF
C6297 a_26402_57174# a_26402_56170# 1.00fF
C6298 a_20286_72234# VDD 0.62fF
C6299 a_1761_49007# a_12381_43957# 1.94fF
C6300 a_28115_43447# VDD 0.61fF
C6301 a_12895_13967# a_12985_16367# 0.99fF
C6302 a_3247_20495# a_6816_19355# 0.32fF
C6303 a_22294_21906# a_22386_21540# 0.32fF
C6304 a_31768_7638# a_12727_15529# 0.41fF
C6305 a_42466_62194# VDD 0.51fF
C6306 a_35601_27497# VDD 6.11fF
C6307 a_7755_54999# VDD 0.32fF
C6308 vcm_commonmode a_28410_12504# 0.87fF
C6309 ctopn a_29414_9492# 3.58fF
C6310 a_3607_34639# VDD 3.53fF
C6311 ctopn a_45478_16520# 3.59fF
C6312 a_42985_46831# a_49494_55166# 0.30fF
C6313 vcm_commonmode a_49402_62194# 0.30fF
C6314 a_36613_48169# a_37446_63198# 0.42fF
C6315 a_2004_42453# a_1586_18695# 0.44fF
C6316 a_18611_52047# a_23390_69222# 0.38fF
C6317 vcm_commonmode a_20286_68218# 0.31fF
C6318 a_2099_59861# a_3339_32463# 1.50fF
C6319 a_36797_27497# a_37446_13508# 0.38fF
C6320 a_29322_59182# a_29414_59182# 0.32fF
C6321 a_12985_7663# VDD 11.61fF
C6322 a_4608_63811# VDD 0.63fF
C6323 a_38557_32143# a_34482_29941# 1.24fF
C6324 a_48490_71230# VDD 0.61fF
C6325 vcm_commonmode a_23390_21540# 0.87fF
C6326 a_19629_39631# VDD 1.80fF
C6327 a_27314_17890# a_27406_17524# 0.32fF
C6328 a_30764_7638# a_12727_15529# 0.41fF
C6329 a_44474_59182# ctopp 3.59fF
C6330 a_33430_64202# a_33430_63198# 1.23fF
C6331 a_46390_12870# a_46482_12504# 0.32fF
C6332 a_30155_32375# VDD 1.43fF
C6333 vcm_commonmode a_28410_17524# 0.87fF
C6334 a_24893_37429# a_27271_37455# 1.69fF
C6335 vcm_commonmode a_49402_24918# 0.30fF
C6336 a_33694_30761# a_30788_28487# 0.91fF
C6337 a_27406_13508# VDD 0.51fF
C6338 a_22632_42919# VDD 1.57fF
C6339 a_2411_26133# a_1591_26159# 0.34fF
C6340 a_6775_53877# VDD 1.38fF
C6341 a_25398_22544# a_25398_21540# 1.00fF
C6342 vcm_commonmode a_34342_13874# 0.31fF
C6343 a_16746_69224# VDD 33.20fF
C6344 a_32426_13508# a_33430_13508# 0.97fF
C6345 a_32181_36893# VDD 0.97fF
C6346 a_17599_52263# a_22386_55166# 0.47fF
C6347 a_3339_30503# a_24768_27247# 0.57fF
C6348 a_26063_30511# a_25971_29967# 0.33fF
C6349 a_37446_68218# a_38450_68218# 0.97fF
C6350 a_17599_52263# a_12257_56623# 0.40fF
C6351 vcm_commonmode a_20286_56170# 0.31fF
C6352 a_2603_64783# VDD 1.05fF
C6353 a_26523_28111# a_11067_23759# 1.28fF
C6354 a_12869_2741# a_22026_27497# 1.10fF
C6355 a_12355_15055# a_16746_61192# 2.28fF
C6356 a_21057_30669# VDD 0.40fF
C6357 a_2411_26133# a_1591_40303# 0.34fF
C6358 a_45478_57174# a_45478_56170# 1.00fF
C6359 a_18370_56170# a_19374_56170# 0.97fF
C6360 vcm_commonmode a_49494_59182# 0.91fF
C6361 a_11619_56615# a_10515_63143# 2.04fF
C6362 ctopn a_19374_19532# 3.59fF
C6363 a_4443_46607# a_2021_17973# 0.47fF
C6364 a_4446_40553# VDD 0.66fF
C6365 a_41370_21906# a_41462_21540# 0.32fF
C6366 a_5363_25321# VDD 0.62fF
C6367 a_22386_58178# a_22386_57174# 1.00fF
C6368 a_48490_60186# ctopp 3.43fF
C6369 a_41967_31375# a_12985_19087# 0.41fF
C6370 a_6662_34025# VDD 1.37fF
C6371 vcm_commonmode a_29414_18528# 0.87fF
C6372 vcm_commonmode a_19282_61190# 0.31fF
C6373 a_29414_16520# a_29414_15516# 1.00fF
C6374 ctopn a_47486_22544# 3.57fF
C6375 a_13183_52047# a_12727_67753# 0.40fF
C6376 a_43470_58178# ctopp 3.59fF
C6377 a_48398_59182# a_48490_59182# 0.32fF
C6378 a_2971_37589# a_3137_37589# 0.75fF
C6379 a_12447_29199# a_35815_31751# 0.57fF
C6380 a_18278_10862# a_18370_10496# 0.32fF
C6381 a_20378_62194# ctopp 3.59fF
C6382 a_16746_70228# VDD 33.20fF
C6383 a_23599_38007# VDD 0.60fF
C6384 vcm_commonmode a_20378_55166# 0.84fF
C6385 a_77451_38925# VDD 109.09fF
C6386 a_46390_17890# a_46482_17524# 0.32fF
C6387 vcm_commonmode a_23298_70226# 0.31fF
C6388 a_40366_58178# vcm_commonmode 0.31fF
C6389 a_33338_60186# a_33430_60186# 0.32fF
C6390 vcm_commonmode a_38450_10496# 0.87fF
C6391 a_21187_29415# a_36507_31573# 0.39fF
C6392 ctopn a_43470_14512# 3.59fF
C6393 a_17507_52047# a_22989_48437# 0.32fF
C6394 a_16955_52047# a_27869_50095# 1.19fF
C6395 a_1803_19087# a_12801_38517# 1.33fF
C6396 a_1895_71482# VDD 0.85fF
C6397 a_26402_71230# ctopp 3.40fF
C6398 ctopn a_22386_20536# 3.59fF
C6399 a_36395_44265# VDD 0.65fF
C6400 a_25787_28327# a_12983_63151# 0.40fF
C6401 a_42718_27497# a_44474_11500# 0.38fF
C6402 a_28318_18894# a_28410_18528# 0.32fF
C6403 a_31768_7638# a_31422_9492# 0.38fF
C6404 a_26748_7638# a_12727_13353# 0.41fF
C6405 a_44474_22544# a_44474_21540# 1.00fF
C6406 a_18979_30287# a_30565_30199# 1.38fF
C6407 a_17366_61190# a_18370_61190# 0.97fF
C6408 a_2327_27247# VDD 0.51fF
C6409 a_34434_8488# VDD 0.58fF
C6410 a_23390_68218# a_23390_67214# 1.00fF
C6411 a_34251_52263# a_12981_62313# 0.40fF
C6412 vcm_commonmode a_25398_62194# 0.87fF
C6413 ctopn a_48490_23548# 3.46fF
C6414 a_11067_46823# a_24959_30503# 0.77fF
C6415 a_1761_50639# a_8491_41383# 0.50fF
C6416 a_7571_26151# VDD 6.49fF
C6417 a_17712_7638# a_17366_13508# 0.38fF
C6418 a_40675_27791# a_41462_13508# 0.38fF
C6419 vcm_commonmode a_41370_8854# 0.31fF
C6420 a_33864_28111# a_12985_19087# 0.41fF
C6421 vcm_commonmode a_33430_15516# 0.87fF
C6422 ctopn a_22386_12504# 3.59fF
C6423 a_11602_25071# a_11430_26159# 0.61fF
C6424 a_44474_57174# ctopp 3.58fF
C6425 a_37446_56170# a_38450_56170# 0.97fF
C6426 a_23507_42089# VDD 0.59fF
C6427 vcm_commonmode a_31422_71230# 0.86fF
C6428 a_20378_8488# a_21382_8488# 0.97fF
C6429 a_19282_55166# a_19374_55166# 0.32fF
C6430 vcm_commonmode a_43470_11500# 0.87fF
C6431 a_11067_67279# a_17488_48731# 2.39fF
C6432 a_22386_67214# VDD 0.51fF
C6433 a_4674_40277# a_4495_35925# 0.42fF
C6434 a_9135_29423# VDD 0.59fF
C6435 a_8531_70543# a_11145_60431# 0.68fF
C6436 a_48490_16520# a_48490_15516# 1.00fF
C6437 vcm_commonmode a_47486_24552# 0.84fF
C6438 ctopn a_17366_21540# 3.42fF
C6439 a_28756_55394# a_28410_68218# 0.38fF
C6440 vcm_commonmode a_29322_67214# 0.31fF
C6441 a_36613_48169# a_12727_67753# 0.40fF
C6442 a_21382_70226# a_22386_70226# 0.97fF
C6443 a_33430_19532# a_33430_18528# 1.00fF
C6444 a_1586_18695# a_7571_16917# 0.80fF
C6445 a_38450_58178# a_39454_58178# 0.97fF
C6446 a_1803_20719# a_2235_31055# 0.42fF
C6447 a_37354_10862# a_37446_10496# 0.32fF
C6448 a_17869_28585# VDD 0.85fF
C6449 a_26748_7638# a_10515_23975# 0.41fF
C6450 a_29414_68218# ctopp 3.59fF
C6451 ctopn a_22386_17524# 3.59fF
C6452 a_3339_32463# a_8273_42479# 0.91fF
C6453 a_19374_9492# VDD 0.51fF
C6454 a_36797_27497# a_37446_7484# 0.34fF
C6455 vcm_commonmode a_49494_57174# 0.89fF
C6456 a_35438_16520# VDD 0.51fF
C6457 a_30534_49393# VDD 0.36fF
C6458 a_41872_29423# a_43470_71230# 0.38fF
C6459 a_8273_42479# a_7841_29673# 0.47fF
C6460 a_19374_60186# a_19374_59182# 1.00fF
C6461 vcm_commonmode a_26310_9858# 0.31fF
C6462 a_11067_13095# a_7737_16917# 0.58fF
C6463 a_42709_29199# a_12985_19087# 0.40fF
C6464 a_23298_11866# a_23390_11500# 0.32fF
C6465 vcm_commonmode a_42374_16886# 0.31fF
C6466 a_28817_29111# a_33864_28111# 0.51fF
C6467 a_31768_55394# VDD 6.80fF
C6468 a_21371_52263# a_26402_60186# 0.38fF
C6469 a_28410_15516# a_28410_14512# 1.00fF
C6470 a_41261_28335# a_42466_67214# 0.38fF
C6471 a_17599_52263# a_10975_66407# 0.40fF
C6472 a_47394_18894# a_47486_18528# 0.32fF
C6473 a_2843_71829# a_4119_70741# 0.56fF
C6474 vcm_commonmode a_36717_47375# 10.02fF
C6475 a_8583_33551# a_21187_29415# 0.33fF
C6476 a_6467_55527# a_6559_59663# 0.67fF
C6477 a_36442_61190# a_37446_61190# 0.97fF
C6478 a_4482_57863# a_7479_54439# 0.42fF
C6479 a_27314_24918# a_27406_24552# 0.32fF
C6480 a_34297_35516# VDD 1.07fF
C6481 a_11711_12559# a_11455_12157# 0.47fF
C6482 a_12549_44212# a_12713_43011# 0.84fF
C6483 a_27406_7484# VDD 1.23fF
C6484 a_42466_68218# a_42466_67214# 1.00fF
C6485 a_28756_55394# a_28410_56170# 0.38fF
C6486 a_18703_29199# a_15607_46805# 0.95fF
C6487 a_10956_14459# VDD 0.64fF
C6488 vcm_commonmode a_34434_68218# 0.87fF
C6489 a_39389_52271# a_12901_66959# 0.40fF
C6490 a_43270_27791# a_45478_19532# 0.38fF
C6491 a_32772_7638# a_12899_10927# 0.41fF
C6492 a_9503_26151# a_12985_19087# 0.41fF
C6493 a_21382_64202# VDD 0.51fF
C6494 a_24302_62194# a_24394_62194# 0.32fF
C6495 a_49402_58178# VDD 0.31fF
C6496 a_29414_56170# ctopp 3.40fF
C6497 a_2824_70197# VDD 0.43fF
C6498 a_1761_52815# a_13909_35395# 1.16fF
C6499 a_23565_38565# VDD 1.44fF
C6500 ctopn a_23390_18528# 3.59fF
C6501 a_27406_69222# a_27406_68218# 1.00fF
C6502 vcm_commonmode a_28318_64202# 0.31fF
C6503 a_2283_15797# a_3023_16341# 1.02fF
C6504 a_22843_29415# a_11067_46823# 0.69fF
C6505 a_35403_50069# VDD 0.35fF
C6506 a_43470_72234# a_44474_72234# 0.97fF
C6507 a_17712_7638# a_12877_14441# 0.40fF
C6508 a_7571_29199# a_10964_25615# 0.54fF
C6509 a_37354_55166# a_37446_55166# 0.32fF
C6510 a_39454_8488# a_40458_8488# 0.97fF
C6511 a_17366_8488# a_17366_7484# 1.00fF
C6512 a_11619_56615# a_7571_26151# 1.84fF
C6513 a_24740_7638# a_12985_7663# 0.41fF
C6514 a_2021_22325# a_5691_36727# 0.41fF
C6515 a_29322_57174# a_29414_57174# 0.32fF
C6516 a_6835_46823# a_3780_56347# 0.34fF
C6517 a_32334_15882# a_32426_15516# 0.32fF
C6518 a_13357_32143# a_25263_29981# 0.37fF
C6519 a_40458_70226# a_41462_70226# 0.97fF
C6520 a_16362_18528# a_12899_10927# 1.27fF
C6521 a_10791_57711# a_10957_57711# 0.69fF
C6522 a_4379_18756# VDD 0.58fF
C6523 a_1586_69367# a_2686_70223# 0.69fF
C6524 a_18979_30287# a_26523_29199# 0.38fF
C6525 a_7210_55081# a_6559_59879# 0.50fF
C6526 vcm_commonmode a_48490_13508# 0.87fF
C6527 a_28410_61190# ctopp 3.59fF
C6528 ctopn a_32426_10496# 3.59fF
C6529 a_30418_69222# VDD 0.51fF
C6530 a_15959_36415# VDD 0.99fF
C6531 vcm_commonmode a_16362_19532# 4.47fF
C6532 a_21382_16520# a_22386_16520# 0.97fF
C6533 vcm_commonmode a_34434_56170# 0.87fF
C6534 vcm_commonmode a_37354_69222# 0.31fF
C6535 a_30326_71230# a_30418_71230# 0.32fF
C6536 a_38450_60186# a_38450_59182# 1.00fF
C6537 a_37446_22544# VDD 0.51fF
C6538 vcm_commonmode a_17366_8488# 1.81fF
C6539 a_28410_65206# VDD 0.51fF
C6540 a_4563_32900# a_4259_32687# 0.62fF
C6541 a_1586_36727# a_1591_36501# 0.38fF
C6542 a_27406_63198# a_27406_62194# 1.00fF
C6543 a_42374_11866# a_42466_11500# 0.32fF
C6544 a_6162_28487# a_5211_24759# 0.46fF
C6545 a_10975_66407# a_16746_65208# 2.28fF
C6546 a_47486_15516# a_47486_14512# 1.00fF
C6547 a_1929_12131# a_3327_9308# 2.21fF
C6548 vcm_commonmode a_44382_22910# 0.31fF
C6549 a_32426_70226# ctopp 3.58fF
C6550 a_16101_31029# a_14625_30761# 0.45fF
C6551 a_3339_32463# a_2787_32679# 0.35fF
C6552 a_3339_43023# a_5915_30287# 1.39fF
C6553 a_1761_50639# a_12801_38517# 0.49fF
C6554 a_27245_41829# VDD 1.47fF
C6555 vcm_commonmode a_35346_65206# 0.31fF
C6556 a_41872_29423# a_12355_65103# 0.40fF
C6557 a_32426_9492# a_32426_8488# 1.00fF
C6558 a_17274_24918# VDD 0.37fF
C6559 a_46390_24918# a_46482_24552# 0.32fF
C6560 a_9263_24501# a_10073_23439# 0.86fF
C6561 ctopn a_27406_15516# 3.59fF
C6562 a_5449_25071# a_4351_26703# 0.88fF
C6563 vcm_commonmode a_33430_61190# 0.87fF
C6564 a_27406_67214# a_28410_67214# 0.97fF
C6565 a_5755_14709# a_5465_14967# 0.46fF
C6566 a_33430_14512# VDD 0.51fF
C6567 a_13909_38659# a_13097_37455# 1.68fF
C6568 a_11759_51959# a_11855_51959# 0.32fF
C6569 a_28318_55166# VDD 0.35fF
C6570 a_37919_28111# a_12899_10927# 0.41fF
C6571 a_43269_29967# a_12727_13353# 0.41fF
C6572 a_11067_46823# a_41334_29575# 0.68fF
C6573 a_43378_62194# a_43470_62194# 0.32fF
C6574 a_12899_3855# VDD 3.39fF
C6575 vcm_commonmode a_40366_14878# 0.31fF
C6576 ctopn a_37446_11500# 3.59fF
C6577 a_23395_52047# a_26523_28111# 4.90fF
C6578 a_4123_37013# VDD 0.98fF
C6579 vcm_commonmode a_19282_20902# 0.31fF
C6580 a_28757_27247# a_28305_28879# 0.75fF
C6581 a_27183_40229# VDD 1.11fF
C6582 a_46482_69222# a_46482_68218# 1.00fF
C6583 a_40675_27791# a_41462_7484# 0.34fF
C6584 a_17712_7638# a_17366_7484# 0.34fF
C6585 a_3391_15797# VDD 0.43fF
C6586 vcm_commonmode a_37446_70226# 0.87fF
C6587 a_36442_8488# a_36442_7484# 1.00fF
C6588 a_38450_23548# VDD 0.52fF
C6589 a_21382_58178# ctopp 3.59fF
C6590 a_5211_24759# a_7377_18012# 0.37fF
C6591 a_35438_66210# VDD 0.51fF
C6592 a_18370_24552# m3_18272_24702# 2.45fF
C6593 a_42807_31849# VDD 0.59fF
C6594 vcm_commonmode a_18370_16520# 0.88fF
C6595 a_16955_52047# a_14831_50095# 0.58fF
C6596 a_48398_57174# a_48490_57174# 0.32fF
C6597 a_12877_14441# a_16362_14512# 19.89fF
C6598 vcm_commonmode a_45386_23914# 0.31fF
C6599 a_13947_43447# VDD 0.60fF
C6600 vcm_commonmode a_42374_66210# 0.31fF
C6601 a_29414_58178# a_30418_58178# 0.97fF
C6602 a_47486_19532# VDD 0.51fF
C6603 a_2872_44111# VDD 7.12fF
C6604 a_24394_9492# a_25398_9492# 0.97fF
C6605 a_10501_55535# VDD 0.34fF
C6606 vcm_commonmode a_19282_12870# 0.31fF
C6607 a_25398_13508# a_25398_12504# 1.00fF
C6608 a_38450_67214# ctopp 3.59fF
C6609 a_39299_48783# a_44474_55166# 0.54fF
C6610 a_25787_28327# a_33430_63198# 0.42fF
C6611 a_40458_16520# a_41462_16520# 0.97fF
C6612 vcm_commonmode a_17712_7638# 10.74fF
C6613 a_49402_71230# a_49494_71230# 0.32fF
C6614 a_19720_55394# a_19374_69222# 0.38fF
C6615 a_39223_32463# a_39454_15516# 0.38fF
C6616 a_46482_63198# a_46482_62194# 1.00fF
C6617 a_27016_29587# VDD 0.47fF
C6618 a_43269_29967# a_10515_23975# 0.41fF
C6619 a_1761_52815# a_13005_35823# 2.19fF
C6620 vcm_commonmode a_26402_58178# 0.87fF
C6621 a_35438_72234# m3_35340_72146# 2.80fF
C6622 a_1761_40847# VDD 7.88fF
C6623 a_35683_50613# VDD 0.53fF
C6624 a_6737_60431# VDD 0.98fF
C6625 a_5363_30503# a_9765_32143# 0.54fF
C6626 vcm_commonmode a_19282_17890# 0.31fF
C6627 a_46482_67214# a_47486_67214# 0.97fF
C6628 a_41872_29423# ctopp 2.63fF
C6629 a_15775_44581# VDD 0.94fF
C6630 vcm_commonmode a_43470_67214# 0.87fF
C6631 a_5531_53903# VDD 0.32fF
C6632 a_39454_63198# VDD 0.57fF
C6633 a_27132_28585# VDD 0.45fF
C6634 a_6559_59663# a_8132_53511# 0.34fF
C6635 a_6372_38279# a_1761_27791# 0.31fF
C6636 a_7571_29199# a_7841_12167# 0.76fF
C6637 a_28318_13874# a_28410_13508# 0.32fF
C6638 a_14287_51175# a_18370_55166# 0.43fF
C6639 a_33338_68218# a_33430_68218# 0.32fF
C6640 vcm_commonmode a_46390_63198# 0.31fF
C6641 a_4191_33449# a_4443_46607# 0.53fF
C6642 a_49494_72234# a_49494_71230# 1.00fF
C6643 a_33430_59182# VDD 0.51fF
C6644 a_6775_53877# a_9507_53877# 0.33fF
C6645 a_32426_7484# a_33430_7484# 0.97fF
C6646 vcm_commonmode a_40458_9492# 0.87fF
C6647 a_41967_31375# VDD 6.70fF
C6648 a_37446_64202# ctopp 3.59fF
C6649 ctopn a_42466_13508# 3.59fF
C6650 a_12899_2767# a_32951_27247# 0.37fF
C6651 vcm_commonmode a_40366_59182# 0.31fF
C6652 vcm_commonmode a_20378_22544# 0.87fF
C6653 a_36432_42919# VDD 1.67fF
C6654 a_3339_43023# a_12663_39783# 1.71fF
C6655 a_31847_36893# a_1761_30511# 1.14fF
C6656 a_9668_51451# VDD 0.31fF
C6657 a_43470_9492# a_44474_9492# 0.97fF
C6658 a_26402_64202# a_27406_64202# 0.97fF
C6659 a_30412_34337# VDD 1.19fF
C6660 a_44474_13508# a_44474_12504# 1.00fF
C6661 vcm_commonmode a_20286_18894# 0.31fF
C6662 a_12357_37999# a_12473_42869# 0.65fF
C6663 ctopn m3_34336_24702# 0.36fF
C6664 a_24413_39087# a_16152_37601# 0.60fF
C6665 a_45478_21540# VDD 0.51fF
C6666 vcm_commonmode a_48490_7484# 0.68fF
C6667 a_23390_22544# a_24394_22544# 0.97fF
C6668 vcm_commonmode a_16362_14512# 4.47fF
C6669 a_5449_37191# VDD 0.53fF
C6670 a_46482_69222# ctopp 3.59fF
C6671 a_4842_45467# a_1689_10396# 0.42fF
C6672 a_22386_10496# VDD 0.51fF
C6673 vcm_commonmode a_42466_64202# 0.87fF
C6674 a_37446_60186# VDD 0.51fF
C6675 vcm_commonmode a_29322_10862# 0.31fF
C6676 a_23747_31055# VDD 0.59fF
C6677 a_44474_65206# ctopp 3.59fF
C6678 a_2021_22325# a_4685_37583# 0.92fF
C6679 a_12357_37999# a_31004_40743# 0.33fF
C6680 a_4031_73095# VDD 0.39fF
C6681 a_43362_28879# a_12981_59343# 0.40fF
C6682 a_34434_67214# a_34434_66210# 1.00fF
C6683 vcm_commonmode a_44382_60186# 0.31fF
C6684 a_3024_67191# a_4339_64521# 0.57fF
C6685 vcm_commonmode a_21382_23548# 0.87fF
C6686 a_14354_32117# a_10506_29967# 0.38fF
C6687 a_5915_35943# a_11602_25071# 0.36fF
C6688 a_20899_44211# VDD 1.66fF
C6689 a_21371_52263# a_12983_63151# 0.40fF
C6690 vcm_commonmode a_18370_66210# 0.88fF
C6691 a_36797_27497# a_37446_11500# 0.38fF
C6692 a_1853_27247# config_2_in[1] 0.39fF
C6693 a_6883_37019# a_4495_35925# 0.69fF
C6694 a_33864_28111# VDD 6.31fF
C6695 a_32772_7638# a_32426_23548# 0.36fF
C6696 a_30418_65206# a_30418_64202# 1.00fF
C6697 a_47394_13874# a_47486_13508# 0.32fF
C6698 a_32327_35839# VDD 0.69fF
C6699 vcm_commonmode a_30418_19532# 0.87fF
C6700 a_13716_43047# a_13005_43983# 0.35fF
C6701 a_28756_55394# a_12981_62313# 0.40fF
C6702 a_27535_30503# a_34062_47607# 0.31fF
C6703 a_17366_15516# VDD 0.57fF
C6704 VDD clk_vcm 4.02fF
C6705 a_36629_27791# a_36442_13508# 0.38fF
C6706 a_24394_23548# a_24394_22544# 1.00fF
C6707 vcm_commonmode a_24302_15882# 0.31fF
C6708 a_17366_63198# ctopp 3.49fF
C6709 a_19967_41781# a_29269_40741# 0.59fF
C6710 a_33338_56170# a_33430_56170# 0.32fF
C6711 a_12907_56399# VDD 26.81fF
C6712 a_18370_66210# a_18370_65206# 1.00fF
C6713 a_3339_43023# inp_analog 0.57fF
C6714 a_19374_14512# a_20378_14512# 0.97fF
C6715 a_1757_38677# VDD 0.66fF
C6716 a_3339_30503# a_9529_28335# 0.34fF
C6717 a_27406_11500# VDD 0.51fF
C6718 a_3143_66972# a_6515_67477# 0.39fF
C6719 vcm_commonmode a_49494_65206# 0.91fF
C6720 a_35438_69222# a_36442_69222# 0.97fF
C6721 vcm_commonmode a_22294_71230# 0.31fF
C6722 a_21371_52263# a_26402_72234# 0.34fF
C6723 VDD config_2_in[14] 1.69fF
C6724 a_30418_61190# a_30418_60186# 1.00fF
C6725 a_3016_60949# a_3714_58345# 0.91fF
C6726 a_16270_55166# a_16362_55166# 0.32fF
C6727 a_31422_24552# VDD 0.60fF
C6728 vcm_commonmode a_34342_11866# 0.31fF
C6729 a_9135_27239# a_11067_21583# 0.41fF
C6730 a_11659_66567# VDD 1.01fF
C6731 a_45478_64202# a_46482_64202# 0.97fF
C6732 a_5515_32661# VDD 0.35fF
C6733 vcm_commonmode a_38358_24918# 0.31fF
C6734 a_2292_43291# a_2539_42106# 0.37fF
C6735 a_25971_52263# a_12727_67753# 0.40fF
C6736 a_18151_52263# a_24394_68218# 0.38fF
C6737 a_17274_70226# a_17366_70226# 0.32fF
C6738 a_10515_63143# a_5363_30503# 1.45fF
C6739 a_41462_55166# VDD 0.60fF
C6740 a_42466_22544# a_43470_22544# 0.97fF
C6741 a_16746_63200# VDD 33.19fF
C6742 a_42709_29199# VDD 6.85fF
C6743 a_33430_57174# VDD 0.51fF
C6744 a_33430_65206# a_34434_65206# 0.97fF
C6745 a_7580_61751# a_8500_58799# 0.42fF
C6746 vcm_commonmode a_33430_20536# 0.87fF
C6747 vcm_commonmode a_22386_63198# 0.92fF
C6748 a_29414_17524# a_29414_16520# 1.00fF
C6749 vcm_commonmode a_40366_57174# 0.31fF
C6750 a_39389_52271# a_39454_71230# 0.38fF
C6751 a_2695_58951# VDD 0.68fF
C6752 a_6607_42167# a_6752_29941# 0.42fF
C6753 vcm_commonmode a_16746_9490# 5.36fF
C6754 a_24394_23548# a_25398_23548# 0.97fF
C6755 a_18151_52263# VDD 15.64fF
C6756 a_17599_52263# a_22386_60186# 0.38fF
C6757 vcm_commonmode a_16746_59184# 5.36fF
C6758 a_21382_66210# a_22386_66210# 0.97fF
C6759 a_48490_7484# m3_48392_7346# 2.80fF
C6760 a_39244_41953# VDD 1.98fF
C6761 a_2191_68565# a_2927_68565# 0.53fF
C6762 a_38557_32143# a_38450_67214# 0.38fF
C6763 vcm_commonmode a_29760_55394# 10.02fF
C6764 a_23736_7638# a_23390_13508# 0.38fF
C6765 a_47486_62194# VDD 0.51fF
C6766 a_15607_46805# a_29175_28335# 0.44fF
C6767 a_32334_61190# a_32426_61190# 0.32fF
C6768 a_9503_26151# VDD 8.99fF
C6769 a_45478_55166# m3_45380_55078# 2.81fF
C6770 vcm_commonmode a_33430_12504# 0.87fF
C6771 ctopn a_34434_9492# 3.58fF
C6772 a_18370_68218# VDD 0.52fF
C6773 a_20359_29199# a_4811_34855# 0.41fF
C6774 a_49494_65206# a_49494_64202# 1.00fF
C6775 a_19559_35561# VDD 0.61fF
C6776 a_13716_43047# a_30412_42589# 0.46fF
C6777 a_18278_7850# VDD 0.62fF
C6778 a_18151_52263# a_24394_56170# 0.38fF
C6779 a_21382_71230# a_21382_70226# 1.00fF
C6780 a_28547_51175# a_12901_66959# 0.40fF
C6781 vcm_commonmode a_25306_68218# 0.31fF
C6782 a_33430_19532# a_34434_19532# 0.97fF
C6783 a_43470_23548# a_43470_22544# 1.00fF
C6784 a_38959_29967# VDD 0.39fF
C6785 a_37446_66210# a_37446_65206# 1.00fF
C6786 a_1923_59583# a_4647_63937# 0.44fF
C6787 a_38450_14512# a_39454_14512# 0.97fF
C6788 vcm_commonmode a_28410_21540# 0.87fF
C6789 a_1586_18695# a_10995_14333# 0.43fF
C6790 vcm_commonmode a_46482_58178# 0.87fF
C6791 a_13097_35279# a_13909_35395# 0.36fF
C6792 a_26321_50095# VDD 0.32fF
C6793 a_39222_48169# a_41427_52263# 0.33fF
C6794 a_17366_20536# a_18370_20536# 0.97fF
C6795 a_49494_61190# a_49494_60186# 1.00fF
C6796 a_35346_8854# a_35438_8488# 0.32fF
C6797 a_2840_66103# a_3295_54421# 0.91fF
C6798 a_33591_32375# VDD 0.41fF
C6799 vcm_commonmode a_33430_17524# 0.87fF
C6800 a_6162_28487# a_9179_22351# 0.60fF
C6801 a_3339_43023# a_4427_30511# 0.55fF
C6802 a_1591_64239# VDD 2.79fF
C6803 vcm_commonmode a_20378_60186# 0.87fF
C6804 a_1586_9991# a_3413_10389# 0.60fF
C6805 a_3339_30503# a_8753_31055# 0.36fF
C6806 a_1761_52815# a_4314_40821# 0.56fF
C6807 a_32426_13508# VDD 0.51fF
C6808 a_32121_44545# VDD 1.44fF
C6809 a_36350_70226# a_36442_70226# 0.32fF
C6810 a_17712_7638# a_17366_11500# 0.38fF
C6811 a_40675_27791# a_41462_11500# 0.38fF
C6812 a_1586_40455# config_2_in[9] 1.16fF
C6813 a_4482_57863# a_3877_57167# 0.32fF
C6814 a_5909_51433# a_6671_51183# 0.33fF
C6815 a_3295_62083# a_3295_54421# 1.02fF
C6816 a_35438_62194# a_35438_61190# 1.00fF
C6817 a_26402_10496# a_26402_9492# 1.00fF
C6818 a_18370_56170# VDD 0.52fF
C6819 vcm_commonmode a_39362_13874# 0.31fF
C6820 a_12621_44099# a_12549_44212# 0.50fF
C6821 a_17274_16886# a_17366_16520# 0.32fF
C6822 a_48490_17524# a_48490_16520# 1.00fF
C6823 vcm_commonmode a_25306_56170# 0.31fF
C6824 a_5915_30287# a_14361_29967# 0.30fF
C6825 a_21187_29415# a_15607_46805# 3.36fF
C6826 a_35438_20536# a_35438_19532# 1.00fF
C6827 a_43470_23548# a_44474_23548# 0.97fF
C6828 a_40458_66210# a_41462_66210# 0.97fF
C6829 ctopn a_24394_19532# 3.59fF
C6830 a_8491_41383# a_8566_39215# 0.80fF
C6831 a_9642_10357# VDD 0.86fF
C6832 a_36717_47375# a_12355_65103# 0.40fF
C6833 a_42718_27497# a_44474_10496# 0.38fF
C6834 a_17366_61190# VDD 0.57fF
C6835 a_19559_34473# VDD 0.59fF
C6836 a_17366_12504# a_18370_12504# 0.97fF
C6837 vcm_commonmode a_34434_18528# 0.87fF
C6838 vcm_commonmode a_24302_61190# 0.31fF
C6839 a_23298_67214# a_23390_67214# 0.32fF
C6840 a_2292_43291# a_2656_45895# 0.34fF
C6841 a_8531_70543# a_4351_67279# 0.44fF
C6842 a_40458_71230# a_40458_70226# 1.00fF
C6843 a_2223_28617# VDD 2.66fF
C6844 a_25398_62194# ctopp 3.59fF
C6845 a_16955_52047# a_26523_28111# 0.41fF
C6846 a_21382_70226# VDD 0.51fF
C6847 a_35932_37601# VDD 1.42fF
C6848 a_38450_58178# VDD 0.51fF
C6849 vcm_commonmode a_25398_55166# 0.84fF
C6850 a_2419_48783# a_2004_42453# 0.54fF
C6851 a_36629_27791# a_36442_7484# 0.35fF
C6852 vcm_commonmode a_16746_57176# 5.36fF
C6853 a_6619_16341# VDD 0.60fF
C6854 a_32318_48695# VDD 0.93fF
C6855 vcm_commonmode a_28318_70226# 0.31fF
C6856 a_10055_58791# a_7000_43541# 0.44fF
C6857 a_36442_20536# a_37446_20536# 0.97fF
C6858 vcm_commonmode a_43470_10496# 0.87fF
C6859 a_8132_53511# a_7050_53333# 0.96fF
C6860 a_25398_63198# a_26402_63198# 0.97fF
C6861 ctopn a_48490_14512# 3.43fF
C6862 a_4427_30511# a_7111_22351# 0.42fF
C6863 a_5877_70197# VDD 4.69fF
C6864 a_31422_71230# ctopp 3.40fF
C6865 ctopn a_27406_20536# 3.59fF
C6866 a_7571_29199# a_5831_39189# 0.67fF
C6867 a_25306_58178# a_25398_58178# 0.32fF
C6868 a_9314_69367# a_1950_59887# 0.61fF
C6869 a_17712_7638# a_12899_11471# 0.40fF
C6870 a_12907_27023# a_43495_28487# 0.46fF
C6871 a_8273_42479# a_4903_31849# 0.65fF
C6872 a_20286_9858# a_20378_9492# 0.32fF
C6873 a_45478_10496# a_45478_9492# 1.00fF
C6874 a_3301_26703# VDD 1.09fF
C6875 a_28410_55166# m3_28312_55078# 2.81fF
C6876 a_2840_66103# a_6467_55527# 1.67fF
C6877 a_39222_48169# a_40458_55166# 0.48fF
C6878 a_7571_26151# a_5363_30503# 0.71fF
C6879 a_39454_8488# VDD 0.58fF
C6880 a_29760_55394# a_29414_63198# 0.42fF
C6881 vcm_commonmode a_30418_62194# 0.87fF
C6882 a_36350_16886# a_36442_16520# 0.32fF
C6883 a_2235_30503# a_7281_29423# 0.96fF
C6884 a_1761_49007# a_4443_46607# 0.39fF
C6885 a_31753_47919# VDD 0.32fF
C6886 a_1923_73087# a_7580_61751# 0.37fF
C6887 a_19374_59182# a_20378_59182# 0.97fF
C6888 vcm_commonmode a_46390_8854# 0.31fF
C6889 a_2840_53511# a_5749_60039# 0.31fF
C6890 a_11067_13095# a_11251_59879# 1.02fF
C6891 vcm_commonmode a_38450_15516# 0.87fF
C6892 ctopn a_27406_12504# 3.59fF
C6893 a_8935_27791# a_9135_27239# 0.50fF
C6894 vcm_commonmode a_17274_58178# 0.33fF
C6895 a_29943_39141# VDD 0.98fF
C6896 a_2952_46805# a_2539_42106# 0.35fF
C6897 a_35601_27497# a_35438_9492# 0.38fF
C6898 a_17366_17524# a_18370_17524# 0.97fF
C6899 a_1908_17141# VDD 0.51fF
C6900 a_10055_58791# a_12877_16911# 24.49fF
C6901 vcm_commonmode a_36442_71230# 0.86fF
C6902 a_34434_21540# a_34434_20536# 1.00fF
C6903 vcm_commonmode a_48490_11500# 0.87fF
C6904 a_4339_64521# a_6775_53877# 0.57fF
C6905 a_32951_27247# a_11067_21583# 0.41fF
C6906 a_21382_24552# a_21382_23548# 1.00fF
C6907 a_27406_67214# VDD 0.51fF
C6908 a_36442_12504# a_37446_12504# 0.97fF
C6909 a_42374_67214# a_42466_67214# 0.32fF
C6910 a_36717_47375# ctopp 2.62fF
C6911 ctopn a_22386_21540# 3.59fF
C6912 a_15607_46805# a_26523_28111# 0.45fF
C6913 a_1761_47919# a_6863_42692# 0.51fF
C6914 a_16863_29415# a_12447_29199# 0.76fF
C6915 vcm_commonmode a_34342_67214# 0.31fF
C6916 a_23736_7638# a_23390_7484# 0.34fF
C6917 a_32582_51701# a_33360_51701# 0.30fF
C6918 a_10055_58791# a_28756_7638# 0.41fF
C6919 a_39223_32463# a_39454_20536# 0.38fF
C6920 a_34434_68218# ctopp 3.59fF
C6921 ctopn a_27406_17524# 3.59fF
C6922 a_28446_31375# a_28305_28879# 0.83fF
C6923 a_24394_9492# VDD 0.51fF
C6924 a_29863_39913# VDD 0.63fF
C6925 a_40458_16520# VDD 0.51fF
C6926 a_28318_7850# a_28410_7484# 0.32fF
C6927 a_8015_21807# VDD 0.37fF
C6928 vcm_commonmode a_31330_9858# 0.31fF
C6929 a_12907_27023# a_33694_30761# 0.59fF
C6930 a_7773_63927# a_1586_51335# 0.52fF
C6931 a_44474_63198# a_45478_63198# 0.97fF
C6932 vcm_commonmode a_47394_16886# 0.31fF
C6933 a_15681_27497# a_18307_27791# 0.45fF
C6934 a_19596_42919# VDD 1.56fF
C6935 a_18370_18528# a_18370_17524# 1.00fF
C6936 a_13669_37429# a_1761_35407# 1.14fF
C6937 a_39223_32463# a_39454_12504# 0.38fF
C6938 a_31422_21540# a_32426_21540# 0.97fF
C6939 a_39362_9858# a_39454_9492# 0.32fF
C6940 a_5211_24759# VDD 4.80fF
C6941 a_43175_28335# a_11067_21583# 0.41fF
C6942 a_42709_29199# a_48490_22544# 0.38fF
C6943 a_22294_64202# a_22386_64202# 0.32fF
C6944 a_1761_34319# VDD 7.43fF
C6945 a_32426_7484# VDD 1.25fF
C6946 a_3280_70501# a_3372_70197# 0.59fF
C6947 vcm_commonmode a_39454_68218# 0.87fF
C6948 a_38450_59182# a_39454_59182# 0.97fF
C6949 a_19282_22910# a_19374_22544# 0.32fF
C6950 a_9503_26151# a_20378_19532# 0.38fF
C6951 a_26402_64202# VDD 0.51fF
C6952 a_18703_29199# a_26523_29199# 0.85fF
C6953 a_18829_29423# VDD 0.51fF
C6954 a_12801_38517# a_19919_38695# 0.80fF
C6955 a_34434_56170# ctopp 3.44fF
C6956 a_35033_38780# VDD 0.87fF
C6957 a_19374_14512# a_19374_13508# 1.00fF
C6958 ctopn a_28410_18528# 3.59fF
C6959 vcm_commonmode a_33338_64202# 0.31fF
C6960 a_12341_3311# a_22386_9492# 0.38fF
C6961 a_36442_17524# a_37446_17524# 0.97fF
C6962 a_1757_49557# VDD 0.65fF
C6963 a_17507_52047# a_11803_55311# 0.57fF
C6964 a_23390_60186# a_24394_60186# 0.97fF
C6965 a_12947_23413# VDD 3.60fF
C6966 a_40458_24552# a_40458_23548# 1.00fF
C6967 a_39223_32463# a_39454_17524# 0.38fF
C6968 a_2939_31573# VDD 0.41fF
C6969 a_25398_12504# a_25398_11500# 1.00fF
C6970 a_20747_27765# a_15681_27497# 1.06fF
C6971 a_12641_43124# a_15459_41781# 2.94fF
C6972 a_39222_48169# a_12981_59343# 0.40fF
C6973 a_4701_43567# VDD 0.31fF
C6974 a_19720_55394# a_12983_63151# 0.40fF
C6975 a_18370_18528# a_19374_18528# 0.97fF
C6976 a_12815_19319# VDD 0.55fF
C6977 a_12818_52521# VDD 0.65fF
C6978 a_1799_29556# a_12473_37429# 0.91fF
C6979 a_33430_61190# ctopp 3.59fF
C6980 ctopn a_37446_10496# 3.59fF
C6981 a_43269_29967# a_47486_22544# 0.38fF
C6982 a_35438_69222# VDD 0.51fF
C6983 a_4563_32900# a_5631_38127# 0.51fF
C6984 a_21856_36513# VDD 1.66fF
C6985 vcm_commonmode a_21290_19898# 0.31fF
C6986 m2_48260_24282# m3_48968_24414# 0.60fF
C6987 a_2021_17973# a_12549_44212# 0.47fF
C6988 a_12757_8207# VDD 0.70fF
C6989 a_17507_52047# a_12981_62313# 0.40fF
C6990 a_11067_13095# a_5691_36727# 0.46fF
C6991 vcm_commonmode a_39454_56170# 0.87fF
C6992 a_1761_34319# a_33486_34191# 0.33fF
C6993 a_9083_13879# VDD 1.20fF
C6994 vcm_commonmode a_42374_69222# 0.31fF
C6995 a_7107_58487# a_8199_58229# 0.47fF
C6996 a_47394_7850# a_47486_7484# 0.32fF
C6997 a_42466_22544# VDD 0.51fF
C6998 vcm_commonmode a_22386_8488# 0.86fF
C6999 a_33430_65206# VDD 0.51fF
C7000 a_4351_67279# a_16219_51183# 0.49fF
C7001 vcm_commonmode a_49402_22910# 0.30fF
C7002 a_37446_70226# ctopp 3.58fF
C7003 a_14625_30761# a_17358_31069# 0.70fF
C7004 a_2656_45895# a_2952_46805# 0.97fF
C7005 a_37491_42359# VDD 0.60fF
C7006 a_31330_69222# a_31422_69222# 0.32fF
C7007 vcm_commonmode a_40366_65206# 0.31fF
C7008 a_37446_18528# a_37446_17524# 1.00fF
C7009 a_37287_51433# VDD 0.40fF
C7010 a_22294_24918# VDD 0.36fF
C7011 a_9135_27239# a_12546_22351# 0.41fF
C7012 a_43270_27791# a_11067_21583# 0.41fF
C7013 a_41370_64202# a_41462_64202# 0.32fF
C7014 a_3339_30503# VDD 11.88fF
C7015 ctopn a_32426_15516# 3.59fF
C7016 a_12663_40871# a_39244_41953# 0.44fF
C7017 a_2124_56891# a_2163_56765# 0.56fF
C7018 vcm_commonmode a_38450_61190# 0.87fF
C7019 a_22015_28111# a_8491_41383# 0.57fF
C7020 a_38450_14512# VDD 0.51fF
C7021 a_1867_45743# VDD 0.36fF
C7022 a_16955_52047# a_20378_68218# 0.38fF
C7023 a_18611_52047# a_12727_67753# 0.40fF
C7024 a_17366_20536# VDD 0.57fF
C7025 a_38358_22910# a_38450_22544# 0.32fF
C7026 a_7295_44647# a_29667_31055# 0.34fF
C7027 a_6835_46823# a_23774_49551# 0.39fF
C7028 a_27406_10496# a_28410_10496# 0.97fF
C7029 vcm_commonmode a_45386_14878# 0.31fF
C7030 ctopn a_42466_11500# 3.59fF
C7031 a_29322_65206# a_29414_65206# 0.32fF
C7032 a_13097_37455# VDD 1.88fF
C7033 a_38450_14512# a_38450_13508# 1.00fF
C7034 vcm_commonmode a_24302_20902# 0.31fF
C7035 a_1761_25071# a_1761_44111# 1.04fF
C7036 a_35647_40229# VDD 0.99fF
C7037 a_11803_55311# a_11067_13095# 1.04fF
C7038 a_20359_29199# a_20635_29415# 0.68fF
C7039 a_12727_13353# VDD 7.23fF
C7040 vcm_commonmode a_42466_70226# 0.87fF
C7041 a_34251_52263# a_35438_71230# 0.38fF
C7042 a_42466_60186# a_43470_60186# 0.97fF
C7043 a_43470_23548# VDD 0.52fF
C7044 a_26402_58178# ctopp 3.59fF
C7045 a_11067_23759# a_12727_15529# 0.35fF
C7046 a_49494_61190# m3_49396_61102# 2.78fF
C7047 a_20286_23914# a_20378_23548# 0.32fF
C7048 a_40458_66210# VDD 0.51fF
C7049 VDD config_1_in[4] 0.80fF
C7050 a_44474_12504# a_44474_11500# 1.00fF
C7051 vcm_commonmode a_23390_16520# 0.87fF
C7052 a_41967_31375# a_42466_24552# 0.45fF
C7053 a_26350_28585# a_26748_7638# 0.36fF
C7054 a_12139_71829# VDD 0.45fF
C7055 a_17274_66210# a_17366_66210# 0.32fF
C7056 a_43267_31055# a_46482_61190# 0.38fF
C7057 a_14287_51175# a_18370_60186# 0.38fF
C7058 a_41462_7484# m3_41364_7346# 2.80fF
C7059 a_7000_43541# a_1803_20719# 0.49fF
C7060 a_17366_12504# VDD 0.57fF
C7061 a_13835_43177# VDD 3.29fF
C7062 a_31422_70226# a_31422_69222# 1.00fF
C7063 vcm_commonmode a_47394_66210# 0.31fF
C7064 a_34780_56398# a_34434_67214# 0.38fF
C7065 a_37446_18528# a_38450_18528# 0.97fF
C7066 a_25419_50959# a_35403_50069# 0.47fF
C7067 vcm_commonmode a_17599_52263# 10.02fF
C7068 a_25462_27497# VDD 0.66fF
C7069 a_38450_55166# m3_38352_55078# 2.81fF
C7070 vcm_commonmode a_24302_12870# 0.31fF
C7071 a_4891_47388# a_6835_46823# 0.64fF
C7072 a_17366_24552# a_18370_24552# 0.97fF
C7073 a_5024_67885# VDD 3.42fF
C7074 a_43470_67214# ctopp 3.59fF
C7075 VDD dummypin[9] 0.97fF
C7076 a_16955_52047# a_20378_56170# 0.38fF
C7077 a_1775_47381# VDD 0.46fF
C7078 a_21371_50959# a_12901_66959# 0.40fF
C7079 a_29322_19898# a_29414_19532# 0.32fF
C7080 a_14287_51175# a_7598_36103# 2.16fF
C7081 ctopn a_23736_7638# 2.62fF
C7082 a_11943_63125# VDD 1.86fF
C7083 a_12355_15055# a_10055_58791# 12.16fF
C7084 a_30418_11500# a_30418_10496# 1.00fF
C7085 vcm_commonmode a_31422_58178# 0.87fF
C7086 a_34342_14878# a_34434_14512# 0.32fF
C7087 a_42283_39095# VDD 0.70fF
C7088 vcm_commonmode a_19282_21906# 0.31fF
C7089 a_38450_72234# m3_38352_72146# 2.80fF
C7090 a_17039_51157# a_21003_49007# 0.34fF
C7091 a_17366_17524# VDD 0.57fF
C7092 a_34359_50639# VDD 0.39fF
C7093 a_36442_72234# a_37446_72234# 0.97fF
C7094 a_4891_47388# a_5612_52520# 0.76fF
C7095 a_10667_60735# VDD 0.36fF
C7096 a_28410_55166# a_29414_55166# 0.97fF
C7097 a_10515_23975# VDD 10.51fF
C7098 vcm_commonmode a_24302_17890# 0.31fF
C7099 a_21371_50959# a_17039_51157# 0.44fF
C7100 a_19374_57174# a_20378_57174# 0.97fF
C7101 a_5599_74549# VDD 1.40fF
C7102 a_22386_15516# a_23390_15516# 0.97fF
C7103 a_2012_33927# a_3143_22364# 0.45fF
C7104 vcm_commonmode a_48490_67214# 0.87fF
C7105 a_36629_27791# a_36442_11500# 0.38fF
C7106 a_2775_46025# a_33360_51701# 0.49fF
C7107 a_30764_7638# a_30418_18528# 0.38fF
C7108 a_44474_63198# VDD 0.57fF
C7109 a_3339_32463# a_6459_30511# 0.32fF
C7110 a_46482_10496# a_47486_10496# 0.97fF
C7111 a_48398_65206# a_48490_65206# 0.32fF
C7112 a_23749_36929# VDD 1.88fF
C7113 a_2927_68565# a_1823_66941# 1.50fF
C7114 a_3911_16065# a_3872_15939# 0.75fF
C7115 a_11619_56615# a_3339_30503# 0.32fF
C7116 vcm_commonmode a_18370_69222# 0.88fF
C7117 a_20378_71230# a_21382_71230# 0.97fF
C7118 a_38450_59182# VDD 0.51fF
C7119 a_11251_59879# a_10515_22671# 2.11fF
C7120 vcm_commonmode a_45478_9492# 0.87fF
C7121 a_39362_23914# a_39454_23548# 0.32fF
C7122 a_2099_64757# VDD 0.50fF
C7123 a_32426_11500# a_33430_11500# 0.97fF
C7124 a_9161_30511# VDD 0.47fF
C7125 a_42466_64202# ctopp 3.59fF
C7126 ctopn a_47486_13508# 3.58fF
C7127 a_45478_72234# VDD 1.65fF
C7128 vcm_commonmode a_45386_59182# 0.31fF
C7129 a_36350_66210# a_36442_66210# 0.32fF
C7130 a_42985_46831# a_12727_58255# 0.40fF
C7131 vcm_commonmode a_25398_22544# 0.87fF
C7132 a_12677_42333# VDD 1.00fF
C7133 vcm_commonmode a_16746_65208# 5.36fF
C7134 a_29760_55394# a_12355_65103# 0.40fF
C7135 a_36797_27497# a_37446_10496# 0.38fF
C7136 a_24740_7638# a_24394_9492# 0.38fF
C7137 a_18370_18528# VDD 0.52fF
C7138 a_5653_60039# VDD 0.52fF
C7139 ctopn a_16362_8488# 1.17fF
C7140 a_39223_32463# a_12899_10927# 0.41fF
C7141 a_36442_24552# a_37446_24552# 0.97fF
C7142 vcm_commonmode a_25306_18894# 0.31fF
C7143 a_18370_66210# ctopp 3.58fF
C7144 a_2012_33927# a_2317_28892# 1.40fF
C7145 a_13643_28327# a_7295_44647# 0.34fF
C7146 ctopn m3_48968_24414# 0.39fF
C7147 a_40783_46831# VDD 0.34fF
C7148 a_48398_19898# a_48490_19532# 0.32fF
C7149 a_12869_2741# a_28959_49783# 0.36fF
C7150 a_1591_59343# a_1775_60663# 0.36fF
C7151 a_33430_62194# a_34434_62194# 0.97fF
C7152 a_49494_11500# a_49494_10496# 1.00fF
C7153 a_33008_28853# VDD 0.31fF
C7154 vcm_commonmode a_21382_14512# 0.87fF
C7155 a_14919_37683# VDD 1.48fF
C7156 a_4842_45467# a_1761_25071# 0.68fF
C7157 a_27406_10496# VDD 0.51fF
C7158 vcm_commonmode a_47486_64202# 0.87fF
C7159 a_32334_20902# a_32426_20536# 0.32fF
C7160 a_23736_7638# a_23390_11500# 0.38fF
C7161 a_32772_7638# a_32426_14512# 0.38fF
C7162 a_42466_60186# VDD 0.51fF
C7163 a_46482_55166# a_47486_55166# 0.97fF
C7164 vcm_commonmode a_34342_10862# 0.31fF
C7165 a_12341_3311# a_11067_21583# 1.00fF
C7166 a_16362_66210# VDD 2.48fF
C7167 a_21290_63198# a_21382_63198# 0.32fF
C7168 a_38450_57174# a_39454_57174# 0.97fF
C7169 a_10509_73193# VDD 0.55fF
C7170 a_11067_66191# a_10975_66407# 2.43fF
C7171 a_2952_66139# a_3295_62083# 0.85fF
C7172 vcm_commonmode a_49402_60186# 0.30fF
C7173 a_41462_15516# a_42466_15516# 0.97fF
C7174 vcm_commonmode a_26402_23548# 0.87fF
C7175 a_1915_35015# a_4095_29423# 0.37fF
C7176 a_1591_12565# VDD 0.44fF
C7177 vcm_commonmode a_23390_66210# 0.87fF
C7178 a_1683_52271# VDD 0.41fF
C7179 a_27752_7638# a_12727_15529# 0.41fF
C7180 a_21382_55166# m3_21284_55078# 2.81fF
C7181 vcm_commonmode a_35438_19532# 0.87fF
C7182 a_41462_58178# a_41462_59182# 1.00fF
C7183 ctopn a_17366_16520# 3.43fF
C7184 a_36717_47375# a_36442_55166# 0.47fF
C7185 vcm_commonmode a_21290_62194# 0.31fF
C7186 a_21371_50959# a_25398_63198# 0.42fF
C7187 a_22386_15516# VDD 0.51fF
C7188 a_39454_71230# a_40458_71230# 0.97fF
C7189 a_2099_59861# a_2419_48783# 1.39fF
C7190 m3_22288_7346# VDD 0.33fF
C7191 vcm_commonmode a_29322_15882# 0.31fF
C7192 a_22386_63198# ctopp 3.64fF
C7193 a_3949_41935# a_3305_38671# 0.85fF
C7194 a_20378_71230# VDD 0.58fF
C7195 a_32426_11500# VDD 0.51fF
C7196 a_16744_41605# VDD 1.79fF
C7197 a_2689_65103# a_1770_14441# 0.41fF
C7198 a_2473_34293# a_2011_34837# 0.81fF
C7199 vcm_commonmode a_27314_71230# 0.31fF
C7200 a_36442_24552# VDD 0.60fF
C7201 vcm_commonmode a_39362_11866# 0.31fF
C7202 a_16746_59184# ctopp 1.68fF
C7203 a_32951_27247# a_12546_22351# 0.41fF
C7204 a_19374_64202# a_19374_63198# 1.23fF
C7205 a_32334_12870# a_32426_12504# 0.32fF
C7206 a_1586_36727# a_2411_26133# 1.03fF
C7207 a_1586_66567# a_2163_63293# 0.35fF
C7208 vcm_commonmode a_43378_24918# 0.31fF
C7209 a_29760_55394# ctopp 2.62fF
C7210 a_6559_45205# VDD 0.41fF
C7211 a_27406_59182# a_27406_58178# 1.00fF
C7212 a_46482_55166# VDD 0.60fF
C7213 a_9135_27239# a_21382_18528# 0.38fF
C7214 a_10680_52245# a_32582_51701# 0.50fF
C7215 a_9179_22351# VDD 2.85fF
C7216 a_38450_57174# VDD 0.51fF
C7217 a_30757_37455# VDD 1.80fF
C7218 a_18370_13508# a_19374_13508# 0.97fF
C7219 vcm_commonmode a_38450_20536# 0.87fF
C7220 a_1761_46287# a_13067_38517# 1.81fF
C7221 a_12757_9295# VDD 0.71fF
C7222 vcm_commonmode a_27406_63198# 0.92fF
C7223 a_23390_68218# a_24394_68218# 0.97fF
C7224 a_2292_17179# a_1895_14906# 0.50fF
C7225 vcm_commonmode a_45386_57174# 0.31fF
C7226 a_26218_48981# VDD 1.04fF
C7227 a_17488_48731# a_13357_32143# 1.82fF
C7228 a_35438_56170# a_35438_55166# 1.00fF
C7229 a_40366_63198# a_40458_63198# 0.32fF
C7230 a_1823_66941# a_1923_54591# 0.41fF
C7231 a_11902_27497# a_11602_25071# 0.33fF
C7232 a_31422_57174# a_31422_56170# 1.00fF
C7233 a_46482_58178# ctopp 3.59fF
C7234 vcm_commonmode a_21382_59182# 0.87fF
C7235 a_2292_17179# a_7203_10383# 0.50fF
C7236 a_2511_42479# VDD 0.48fF
C7237 a_40675_27791# a_41462_10496# 0.38fF
C7238 a_17712_7638# a_17366_10496# 0.38fF
C7239 a_5331_18517# VDD 0.48fF
C7240 a_27314_21906# a_27406_21540# 0.32fF
C7241 a_24740_7638# a_12727_13353# 0.41fF
C7242 a_9669_26703# VDD 1.13fF
C7243 vcm_commonmode a_38450_12504# 0.87fF
C7244 a_20378_60186# ctopp 3.59fF
C7245 ctopn a_39454_9492# 3.58fF
C7246 a_43175_28335# a_12546_22351# 0.41fF
C7247 a_2317_28892# a_4839_21495# 0.41fF
C7248 a_23390_68218# VDD 0.51fF
C7249 a_1803_20719# a_12473_42869# 0.88fF
C7250 a_12381_43957# a_32327_40191# 0.75fF
C7251 a_23298_7850# VDD 0.61fF
C7252 a_45386_58178# a_45478_58178# 0.32fF
C7253 a_13183_52047# a_17366_62194# 0.38fF
C7254 a_8772_63927# a_7803_55509# 0.46fF
C7255 ctopn a_19374_22544# 3.58fF
C7256 a_2606_41079# a_4676_47607# 0.30fF
C7257 vcm_commonmode a_30326_68218# 0.31fF
C7258 a_34342_59182# a_34434_59182# 0.32fF
C7259 a_6743_29673# VDD 0.32fF
C7260 a_11803_55311# a_10515_22671# 2.52fF
C7261 vcm_commonmode a_33430_21540# 0.87fF
C7262 a_1761_50639# a_13909_39747# 1.07fF
C7263 a_32334_17890# a_32426_17524# 0.32fF
C7264 a_42374_72234# a_42466_72234# 0.32fF
C7265 a_8491_27023# a_12727_15529# 0.41fF
C7266 a_19282_60186# a_19374_60186# 0.32fF
C7267 a_2847_23743# VDD 0.60fF
C7268 a_10515_63143# a_8295_47388# 0.54fF
C7269 a_11067_66191# a_10055_58791# 13.42fF
C7270 a_38450_64202# a_38450_63198# 1.23fF
C7271 vcm_commonmode a_38450_17524# 0.87fF
C7272 a_14471_28585# a_12985_25615# 0.50fF
C7273 a_12473_42869# a_23567_42035# 0.39fF
C7274 a_25787_28327# a_12981_59343# 0.40fF
C7275 vcm_commonmode a_25398_60186# 0.87fF
C7276 a_3339_30503# a_12120_29941# 0.61fF
C7277 a_37446_13508# VDD 0.51fF
C7278 a_41462_58178# a_41462_57174# 1.00fF
C7279 a_30418_22544# a_30418_21540# 1.00fF
C7280 a_4839_21495# a_4792_20443# 0.70fF
C7281 a_1823_63677# a_1923_54591# 0.37fF
C7282 a_23390_56170# VDD 0.52fF
C7283 vcm_commonmode a_44382_13874# 0.31fF
C7284 a_24740_7638# a_10515_23975# 0.41fF
C7285 a_13909_39747# a_14963_39783# 3.79fF
C7286 a_2473_34293# VDD 3.55fF
C7287 a_37446_13508# a_38450_13508# 0.97fF
C7288 a_12725_44527# a_12357_37999# 0.53fF
C7289 a_42466_68218# a_43470_68218# 0.97fF
C7290 vcm_commonmode a_30326_56170# 0.31fF
C7291 ctopn a_20378_23548# 3.40fF
C7292 a_2606_41079# a_4443_46607# 0.44fF
C7293 a_43362_28879# a_12516_7093# 0.40fF
C7294 a_11067_13095# a_2292_43291# 0.31fF
C7295 a_19967_41781# a_49876_41198# 1.54fF
C7296 a_16746_57176# ctopp 1.67fF
C7297 a_23390_56170# a_24394_56170# 0.97fF
C7298 ctopn a_29414_19532# 3.59fF
C7299 a_6559_22671# a_1761_44111# 0.30fF
C7300 ctopn a_39673_28111# 2.62fF
C7301 a_19720_55394# a_19374_72234# 0.34fF
C7302 a_46390_21906# a_46482_21540# 0.32fF
C7303 a_28756_7638# a_12877_14441# 0.41fF
C7304 a_22386_61190# VDD 0.51fF
C7305 a_9263_24501# VDD 0.77fF
C7306 a_27406_58178# a_27406_57174# 1.00fF
C7307 a_43270_27791# a_12546_22351# 0.41fF
C7308 a_1915_67477# VDD 0.82fF
C7309 vcm_commonmode a_39454_18528# 0.87fF
C7310 a_13835_43177# a_12663_40871# 4.13fF
C7311 vcm_commonmode a_29322_61190# 0.31fF
C7312 a_34434_16520# a_34434_15516# 1.00fF
C7313 vcm_commonmode a_19374_24552# 0.84fF
C7314 a_26465_48463# a_27509_47695# 0.32fF
C7315 a_5039_42167# a_4674_40277# 0.50fF
C7316 a_19374_19532# a_19374_18528# 1.00fF
C7317 a_5825_20495# VDD 0.92fF
C7318 a_23298_10862# a_23390_10496# 0.32fF
C7319 a_30418_62194# ctopp 3.59fF
C7320 a_26402_70226# VDD 0.51fF
C7321 vcm_commonmode a_30418_55166# 0.84fF
C7322 a_15775_40229# VDD 1.02fF
C7323 vcm_commonmode a_21382_57174# 0.87fF
C7324 a_4495_35925# a_7281_29423# 0.94fF
C7325 a_12815_16519# VDD 0.36fF
C7326 a_31768_55394# a_31422_71230# 0.38fF
C7327 vcm_commonmode a_33338_70226# 0.31fF
C7328 a_42718_27497# a_44474_15516# 0.38fF
C7329 a_38358_60186# a_38450_60186# 0.32fF
C7330 vcm_commonmode a_48490_10496# 0.87fF
C7331 a_17712_7638# a_12985_7663# 0.40fF
C7332 a_4443_46607# a_5595_33205# 0.32fF
C7333 a_41261_28335# a_42466_61190# 0.38fF
C7334 a_36442_71230# ctopp 3.40fF
C7335 ctopn a_32426_20536# 3.59fF
C7336 a_34434_7484# m3_34336_7346# 2.80fF
C7337 a_1803_19087# VDD 8.11fF
C7338 a_1950_59887# a_1923_59583# 0.96fF
C7339 a_25971_52263# a_30418_67214# 0.38fF
C7340 a_33338_18894# a_33430_18528# 0.32fF
C7341 a_19478_51959# VDD 1.21fF
C7342 a_6327_72917# a_6453_71855# 0.47fF
C7343 a_2775_46025# a_6646_50639# 1.50fF
C7344 a_49494_22544# a_49494_21540# 1.00fF
C7345 a_22386_61190# a_23390_61190# 0.97fF
C7346 a_43175_28335# a_46482_23548# 0.38fF
C7347 a_8491_41383# a_13484_39325# 0.33fF
C7348 a_11710_58487# a_10055_58791# 1.00fF
C7349 a_1761_47919# a_33155_40191# 0.42fF
C7350 a_44474_8488# VDD 0.58fF
C7351 a_28410_68218# a_28410_67214# 1.00fF
C7352 vcm_commonmode a_35438_62194# 0.87fF
C7353 a_1823_76181# VDD 3.07fF
C7354 a_14287_51175# a_12901_66959# 0.40fF
C7355 a_2163_64381# VDD 0.56fF
C7356 a_20505_29967# VDD 0.94fF
C7357 vcm_commonmode a_43470_15516# 0.87fF
C7358 ctopn a_32426_12504# 3.59fF
C7359 a_42466_56170# a_43470_56170# 0.97fF
C7360 a_3983_65327# a_4149_65327# 0.72fF
C7361 vcm_commonmode a_22294_58178# 0.31fF
C7362 a_36579_39095# VDD 0.64fF
C7363 a_4674_40277# a_3987_19623# 5.91fF
C7364 a_41443_41855# VDD 0.98fF
C7365 a_25971_52263# a_32823_29397# 1.28fF
C7366 a_7737_16917# VDD 0.34fF
C7367 a_22989_48437# VDD 1.80fF
C7368 vcm_commonmode a_41462_71230# 0.86fF
C7369 a_1923_54591# a_4831_52413# 0.71fF
C7370 a_25398_8488# a_26402_8488# 0.97fF
C7371 a_24302_55166# a_24394_55166# 0.32fF
C7372 a_43270_27791# a_45478_22544# 0.38fF
C7373 a_32426_67214# VDD 0.51fF
C7374 a_27535_30503# a_31659_31751# 0.76fF
C7375 vcm_commonmode a_12877_16911# 6.29fF
C7376 a_18278_15882# a_18370_15516# 0.32fF
C7377 ctopn a_27406_21540# 3.59fF
C7378 a_2292_43291# a_1591_44655# 0.34fF
C7379 a_12559_44527# VDD 0.37fF
C7380 vcm_commonmode a_39362_67214# 0.31fF
C7381 a_26402_70226# a_27406_70226# 0.97fF
C7382 a_38450_19532# a_38450_18528# 1.00fF
C7383 a_32582_51701# a_33748_51727# 0.35fF
C7384 a_2163_54589# VDD 0.53fF
C7385 a_42718_27497# a_12899_10927# 0.41fF
C7386 a_3305_38671# a_1761_37039# 0.68fF
C7387 a_42374_10862# a_42466_10496# 0.32fF
C7388 vcm_commonmode a_20378_13508# 0.87fF
C7389 a_9135_27239# a_12341_3311# 0.53fF
C7390 a_5295_69135# VDD 0.54fF
C7391 a_7479_36495# VDD 0.34fF
C7392 a_39454_68218# ctopp 3.59fF
C7393 ctopn a_32426_17524# 3.59fF
C7394 a_29414_9492# VDD 0.51fF
C7395 vcm_commonmode a_28756_7638# 10.39fF
C7396 a_22989_48437# a_26514_47375# 0.35fF
C7397 a_45478_16520# VDD 0.51fF
C7398 a_47486_72234# a_47486_71230# 1.00fF
C7399 a_11803_55311# a_12901_66665# 1.07fF
C7400 a_16746_71232# a_16362_71230# 2.28fF
C7401 a_7571_29199# a_12341_3311# 0.65fF
C7402 a_24394_60186# a_24394_59182# 1.00fF
C7403 a_1591_21807# VDD 0.39fF
C7404 vcm_commonmode a_36350_9858# 0.31fF
C7405 m3_16264_71142# VDD 0.30fF
C7406 a_31768_7638# a_31422_19532# 0.38fF
C7407 a_7213_62215# a_4298_58951# 0.69fF
C7408 a_28318_11866# a_28410_11500# 0.32fF
C7409 a_17599_52263# a_11067_46823# 0.88fF
C7410 a_32695_43455# a_33155_40191# 0.40fF
C7411 a_38450_72234# VDD 1.36fF
C7412 a_41427_52263# a_12727_58255# 0.40fF
C7413 a_33430_15516# a_33430_14512# 1.00fF
C7414 vcm_commonmode a_16362_22544# 4.47fF
C7415 vcm_commonmode m3_16264_61102# 3.21fF
C7416 a_24893_37429# VDD 1.70fF
C7417 a_17599_52263# a_12355_65103# 0.40fF
C7418 a_30757_37455# a_31280_36165# 0.38fF
C7419 a_8295_47388# a_7571_26151# 0.40fF
C7420 a_35568_49525# a_21187_29415# 0.48fF
C7421 a_4719_71855# a_5023_72068# 0.62fF
C7422 vcm_commonmode a_43470_72234# 0.69fF
C7423 a_9135_27239# a_12985_16367# 0.41fF
C7424 a_7210_55081# VDD 5.29fF
C7425 a_41462_61190# a_42466_61190# 0.97fF
C7426 a_18370_9492# a_18370_8488# 1.00fF
C7427 a_32334_24918# a_32426_24552# 0.33fF
C7428 a_18611_52047# a_10687_52553# 1.13fF
C7429 a_21371_52263# a_10503_52828# 0.46fF
C7430 a_37446_7484# VDD 1.63fF
C7431 a_47486_68218# a_47486_67214# 1.00fF
C7432 a_7862_34025# a_25321_29673# 0.69fF
C7433 a_7623_13621# VDD 0.54fF
C7434 vcm_commonmode a_44474_68218# 0.87fF
C7435 a_31422_64202# VDD 0.51fF
C7436 a_7295_44647# a_19626_31751# 0.83fF
C7437 a_29322_62194# a_29414_62194# 0.32fF
C7438 a_39223_32463# a_39454_21540# 0.38fF
C7439 a_4314_40821# a_4685_37583# 0.81fF
C7440 a_39454_56170# ctopp 3.40fF
C7441 a_7755_70223# VDD 1.13fF
C7442 a_2971_37589# VDD 0.49fF
C7443 ctopn a_33430_18528# 3.59fF
C7444 a_19596_40743# VDD 1.87fF
C7445 vcm_commonmode a_38358_64202# 0.31fF
C7446 a_32426_69222# a_32426_68218# 1.00fF
C7447 a_22386_8488# a_22386_7484# 1.00fF
C7448 a_44474_8488# a_45478_8488# 0.97fF
C7449 a_42374_55166# a_42466_55166# 0.32fF
C7450 a_2419_48783# a_10975_55535# 0.56fF
C7451 a_12341_3311# a_12546_22351# 0.82fF
C7452 a_12981_62313# a_16362_63198# 19.89fF
C7453 a_11143_31599# VDD 0.34fF
C7454 a_34342_57174# a_34434_57174# 0.32fF
C7455 a_37354_15882# a_37446_15516# 0.32fF
C7456 vcm_commonmode a_17274_23914# 0.33fF
C7457 a_3607_34639# a_4248_29967# 0.92fF
C7458 a_45478_70226# a_46482_70226# 0.97fF
C7459 a_19374_19532# VDD 0.51fF
C7460 a_1761_52815# VDD 15.26fF
C7461 a_1644_62037# VDD 0.31fF
C7462 a_38450_61190# ctopp 3.59fF
C7463 ctopn a_42466_10496# 3.59fF
C7464 a_28756_7638# a_28410_23548# 0.38fF
C7465 a_40458_69222# VDD 0.51fF
C7466 a_30139_36649# VDD 0.63fF
C7467 vcm_commonmode a_26310_19898# 0.31fF
C7468 a_17507_52047# a_21382_63198# 0.42fF
C7469 a_12727_67753# a_16362_67214# 1.15fF
C7470 a_26402_16520# a_27406_16520# 0.97fF
C7471 vcm_commonmode a_44474_56170# 0.87fF
C7472 a_1761_47919# VDD 10.44fF
C7473 a_35346_71230# a_35438_71230# 0.32fF
C7474 vcm_commonmode a_47394_69222# 0.31fF
C7475 a_12546_22351# a_12985_16367# 23.46fF
C7476 a_7963_58255# VDD 0.59fF
C7477 a_43470_60186# a_43470_59182# 1.00fF
C7478 a_47486_22544# VDD 0.51fF
C7479 vcm_commonmode a_27406_8488# 0.86fF
C7480 a_38450_65206# VDD 0.51fF
C7481 a_20267_30503# a_7862_34025# 0.34fF
C7482 a_16863_29415# a_38210_30199# 0.60fF
C7483 a_32426_63198# a_32426_62194# 1.00fF
C7484 a_47394_11866# a_47486_11500# 0.32fF
C7485 a_43175_28335# a_43270_27791# 2.50fF
C7486 a_12355_65103# a_16746_65208# 0.41fF
C7487 a_42466_70226# ctopp 3.58fF
C7488 vcm_commonmode m3_16264_8350# 3.05fF
C7489 a_12641_42036# VDD 2.85fF
C7490 vcm_commonmode a_45386_65206# 0.31fF
C7491 a_3987_19623# a_5671_21495# 0.39fF
C7492 a_1761_50639# VDD 8.21fF
C7493 a_11067_67279# ctopn 3.23fF
C7494 a_4674_40277# a_5795_27497# 0.40fF
C7495 a_5363_30503# a_3339_30503# 0.70fF
C7496 a_37446_9492# a_37446_8488# 1.00fF
C7497 a_27314_24918# VDD 0.36fF
C7498 a_7479_67075# VDD 0.32fF
C7499 ctopn a_37446_15516# 3.59fF
C7500 a_32426_67214# a_33430_67214# 0.97fF
C7501 vcm_commonmode a_43470_61190# 0.87fF
C7502 a_17599_52263# ctopp 2.62fF
C7503 a_43470_14512# VDD 0.51fF
C7504 a_22386_20536# VDD 0.51fF
C7505 a_37354_55166# VDD 0.35fF
C7506 a_2959_47113# a_2872_44111# 0.68fF
C7507 a_48398_62194# a_48490_62194# 0.32fF
C7508 ctopn a_47486_11500# 3.58fF
C7509 vcm_commonmode a_29322_20902# 0.31fF
C7510 a_14963_39783# VDD 3.43fF
C7511 vcm_commonmode a_18278_63198# 0.31fF
C7512 a_19282_68218# a_19374_68218# 0.32fF
C7513 vcm_commonmode inp_analog 3.02fF
C7514 a_17843_48981# VDD 0.63fF
C7515 vcm_commonmode a_47486_70226# 0.87fF
C7516 a_1689_10396# a_2315_24540# 0.46fF
C7517 a_12447_29199# a_37919_28111# 0.34fF
C7518 a_41462_8488# a_41462_7484# 1.00fF
C7519 a_18370_7484# a_19374_7484# 0.97fF
C7520 a_48490_23548# VDD 0.56fF
C7521 a_31422_58178# ctopp 3.59fF
C7522 a_45478_66210# VDD 0.51fF
C7523 a_27535_30503# a_34759_31029# 1.15fF
C7524 a_16101_31029# VDD 0.96fF
C7525 vcm_commonmode a_28410_16520# 0.87fF
C7526 a_22386_12504# VDD 0.51fF
C7527 a_32695_43455# VDD 1.10fF
C7528 a_1586_66567# a_2927_68565# 0.70fF
C7529 a_36629_27791# a_36442_10496# 0.38fF
C7530 a_34434_58178# a_35438_58178# 0.97fF
C7531 a_11759_51959# VDD 0.36fF
C7532 a_2775_46025# a_22181_50645# 0.53fF
C7533 a_6559_22671# a_7755_26703# 0.80fF
C7534 a_29414_9492# a_30418_9492# 0.97fF
C7535 a_2913_54991# VDD 0.73fF
C7536 vcm_commonmode a_29322_12870# 0.31fF
C7537 a_2840_66103# a_19576_51701# 0.32fF
C7538 a_30418_13508# a_30418_12504# 1.00fF
C7539 a_48490_67214# ctopp 3.43fF
C7540 a_1954_61677# a_1770_14441# 0.95fF
C7541 a_45478_16520# a_46482_16520# 0.97fF
C7542 a_2004_42453# a_2315_24540# 0.47fF
C7543 a_3247_20495# a_5211_24759# 0.42fF
C7544 a_17366_21540# VDD 0.58fF
C7545 vcm_commonmode a_20378_7484# 0.69fF
C7546 a_33839_28309# VDD 0.94fF
C7547 a_11619_56615# a_1761_52815# 3.16fF
C7548 a_7373_40847# a_7097_40303# 0.36fF
C7549 a_49402_71230# VDD 0.31fF
C7550 vcm_commonmode a_36442_58178# 0.87fF
C7551 vcm_commonmode a_24302_21906# 0.31fF
C7552 a_18370_69222# ctopp 3.58fF
C7553 a_41462_72234# m3_41364_72146# 2.80fF
C7554 a_23789_39100# VDD 1.91fF
C7555 vcm_commonmode a_12355_15055# 6.21fF
C7556 a_37919_28111# a_38450_8488# 0.38fF
C7557 a_22386_17524# VDD 0.51fF
C7558 vcm_commonmode a_29322_17890# 0.31fF
C7559 a_16746_65208# ctopp 1.68fF
C7560 vcm_commonmode a_16746_60188# 5.36fF
C7561 a_20378_67214# a_20378_66210# 1.00fF
C7562 a_21371_52263# a_12981_59343# 0.40fF
C7563 a_12907_27023# a_8491_41383# 0.31fF
C7564 a_22132_44129# VDD 1.66fF
C7565 a_7764_53877# VDD 0.61fF
C7566 a_6224_73095# a_6098_73095# 1.06fF
C7567 a_49494_63198# VDD 1.22fF
C7568 a_41261_28335# a_18979_30287# 0.58fF
C7569 a_16362_69222# VDD 2.49fF
C7570 a_33338_13874# a_33430_13508# 0.32fF
C7571 a_30875_36919# VDD 0.63fF
C7572 a_11719_28023# a_9179_22351# 0.61fF
C7573 a_33641_29967# a_28841_29575# 0.52fF
C7574 a_38358_68218# a_38450_68218# 0.32fF
C7575 a_39222_48169# a_12516_7093# 0.40fF
C7576 vcm_commonmode a_23390_69222# 0.87fF
C7577 a_23736_7638# a_23390_10496# 0.38fF
C7578 a_43470_59182# VDD 0.51fF
C7579 a_37446_7484# a_38450_7484# 0.97fF
C7580 a_12355_15055# a_16362_61190# 1.15fF
C7581 a_47486_64202# ctopp 3.58fF
C7582 a_4427_25071# a_5085_23047# 0.61fF
C7583 a_19282_56170# a_19374_56170# 0.32fF
C7584 a_49494_72234# VDD 2.17fF
C7585 a_7797_13885# a_7917_13885# 0.33fF
C7586 vcm_commonmode a_30418_22544# 0.87fF
C7587 a_7281_29423# a_6752_29941# 0.36fF
C7588 a_21382_69222# a_22386_69222# 0.97fF
C7589 vcm_commonmode a_21382_65206# 0.87fF
C7590 a_35676_49525# a_36821_50095# 0.64fF
C7591 a_23390_18528# VDD 0.51fF
C7592 a_32951_27247# a_12985_16367# 0.41fF
C7593 a_12981_59343# a_12727_58255# 23.54fF
C7594 a_48490_9492# a_49494_9492# 0.97fF
C7595 a_6143_25321# VDD 0.40fF
C7596 ctopn a_21382_8488# 3.40fF
C7597 a_31422_64202# a_32426_64202# 0.97fF
C7598 a_49494_13508# a_49494_12504# 1.00fF
C7599 VDD result_out[3] 0.68fF
C7600 vcm_commonmode a_30326_18894# 0.31fF
C7601 a_23390_66210# ctopp 3.59fF
C7602 a_2021_17973# a_2411_26133# 3.35fF
C7603 a_7050_53333# a_17039_51157# 0.54fF
C7604 a_16270_55166# VDD 0.47fF
C7605 a_28410_22544# a_29414_22544# 0.97fF
C7606 a_3247_20495# a_3339_30503# 0.58fF
C7607 a_6072_56872# VDD 0.39fF
C7608 vcm_commonmode a_26402_14512# 0.87fF
C7609 a_18127_35797# a_13669_39605# 1.30fF
C7610 a_19374_65206# a_20378_65206# 0.97fF
C7611 a_11067_67279# a_36797_27497# 0.41fF
C7612 vcm_commonmode a_21290_55166# 0.30fF
C7613 a_33641_29967# a_30565_30199# 0.58fF
C7614 a_7000_43541# a_7847_40847# 0.37fF
C7615 a_32426_10496# VDD 0.51fF
C7616 VDD result_out[12] 0.49fF
C7617 a_40491_27247# a_43470_8488# 0.38fF
C7618 a_2686_70223# a_5213_70223# 0.43fF
C7619 a_23395_52047# a_27406_71230# 0.38fF
C7620 a_36797_27497# a_37446_15516# 0.38fF
C7621 a_47486_60186# VDD 0.51fF
C7622 vcm_commonmode a_39362_10862# 0.31fF
C7623 a_12947_23413# a_16362_23548# 19.83fF
C7624 a_3339_43023# a_4839_21495# 0.33fF
C7625 a_19374_56170# a_19374_55166# 1.00fF
C7626 a_14926_31849# VDD 4.58fF
C7627 a_12257_56623# a_16746_56172# 2.28fF
C7628 a_39454_67214# a_39454_66210# 1.00fF
C7629 a_38557_32143# a_38450_61190# 0.38fF
C7630 a_12877_16911# a_16746_12502# 0.41fF
C7631 vcm_commonmode a_31422_23548# 0.87fF
C7632 a_27406_7484# m3_27308_7346# 2.80fF
C7633 a_21371_52263# a_26402_67214# 0.38fF
C7634 vcm_commonmode a_28410_66210# 0.87fF
C7635 vcm_commonmode a_16362_72234# 1.71fF
C7636 a_43175_28335# a_12985_16367# 0.41fF
C7637 a_19374_62194# VDD 0.51fF
C7638 a_22291_29415# a_32167_29611# 0.47fF
C7639 a_18278_61190# a_18370_61190# 0.32fF
C7640 a_7803_55509# a_4758_45369# 0.76fF
C7641 a_35438_65206# a_35438_64202# 1.00fF
C7642 a_8531_70543# a_11080_58229# 0.37fF
C7643 vcm_commonmode a_40458_19532# 0.87fF
C7644 ctopn a_22386_16520# 3.59fF
C7645 vcm_commonmode a_26310_62194# 0.31fF
C7646 a_16863_29415# a_15607_46805# 1.53fF
C7647 a_27406_15516# VDD 0.51fF
C7648 a_19374_19532# a_20378_19532# 0.97fF
C7649 a_4482_57863# VDD 11.53fF
C7650 m3_37348_7346# VDD 0.41fF
C7651 a_29414_23548# a_29414_22544# 1.00fF
C7652 a_42718_27497# a_44474_20536# 0.38fF
C7653 vcm_commonmode a_34342_15882# 0.31fF
C7654 a_27406_63198# ctopp 3.64fF
C7655 a_38358_56170# a_38450_56170# 0.32fF
C7656 a_25398_71230# VDD 0.58fF
C7657 a_23390_66210# a_23390_65206# 1.00fF
C7658 a_43267_31055# a_10515_22671# 0.40fF
C7659 a_24394_14512# a_25398_14512# 0.97fF
C7660 a_37446_11500# VDD 0.51fF
C7661 a_40458_69222# a_41462_69222# 0.97fF
C7662 a_2595_47653# a_6559_49557# 0.46fF
C7663 a_19591_50943# VDD 0.33fF
C7664 a_29414_72234# a_30418_72234# 0.97fF
C7665 vcm_commonmode a_32334_71230# 0.31fF
C7666 a_23395_52047# a_25787_28327# 5.02fF
C7667 a_35438_61190# a_35438_60186# 1.00fF
C7668 a_21290_8854# a_21382_8488# 0.32fF
C7669 a_41462_24552# VDD 0.60fF
C7670 vcm_commonmode a_44382_11866# 0.31fF
C7671 a_21382_59182# ctopp 3.59fF
C7672 a_9367_29397# VDD 1.10fF
C7673 a_12381_43957# a_19967_41781# 0.55fF
C7674 a_22294_70226# a_22386_70226# 0.32fF
C7675 a_42718_27497# a_44474_12504# 0.38fF
C7676 a_39362_58178# a_39454_58178# 0.32fF
C7677 a_28756_7638# a_12899_11471# 0.41fF
C7678 a_47486_22544# a_48490_22544# 0.97fF
C7679 a_7479_54439# a_23774_49551# 0.54fF
C7680 a_10680_52245# a_32612_51727# 0.31fF
C7681 a_21382_62194# a_21382_61190# 1.00fF
C7682 a_26350_28585# VDD 0.96fF
C7683 a_43470_57174# VDD 0.51fF
C7684 a_4685_37583# a_7244_39189# 0.57fF
C7685 a_38450_65206# a_39454_65206# 0.97fF
C7686 a_34251_52263# a_35438_58178# 0.38fF
C7687 vcm_commonmode a_43470_20536# 0.87fF
C7688 a_14926_31849# a_18053_28879# 0.31fF
C7689 a_1761_44111# a_2021_22325# 0.86fF
C7690 a_22319_39913# VDD 0.65fF
C7691 vcm_commonmode a_32426_63198# 0.92fF
C7692 a_34434_17524# a_34434_16520# 1.00fF
C7693 a_22015_28111# a_19807_28111# 1.02fF
C7694 a_43470_72234# a_43470_71230# 1.00fF
C7695 a_42709_29199# a_48490_13508# 0.38fF
C7696 a_21382_20536# a_21382_19532# 1.00fF
C7697 m3_22288_72146# VDD 0.33fF
C7698 a_29414_23548# a_30418_23548# 0.97fF
C7699 a_18944_31055# VDD 0.44fF
C7700 a_15459_41781# a_13909_41923# 1.36fF
C7701 a_31422_72234# VDD 1.23fF
C7702 a_26402_66210# a_27406_66210# 0.97fF
C7703 a_34780_56398# a_12727_58255# 0.40fF
C7704 vcm_commonmode a_26402_59182# 0.87fF
C7705 a_28757_27247# a_32823_29397# 0.54fF
C7706 a_12889_40977# VDD 0.74fF
C7707 a_32582_51701# VDD 0.34fF
C7708 vcm_commonmode a_36442_72234# 0.69fF
C7709 a_43270_27791# a_12985_16367# 0.41fF
C7710 a_42718_27497# a_44474_17524# 0.38fF
C7711 a_18979_30287# a_41597_29967# 0.73fF
C7712 a_37354_61190# a_37446_61190# 0.32fF
C7713 vcm_commonmode a_43470_12504# 0.87fF
C7714 a_25398_60186# ctopp 3.59fF
C7715 ctopn a_44474_9492# 3.58fF
C7716 a_28410_68218# VDD 0.51fF
C7717 a_12907_56399# a_8295_47388# 5.06fF
C7718 a_1761_43567# a_12473_42869# 3.14fF
C7719 a_28318_7850# VDD 0.62fF
C7720 ctopn a_24394_22544# 3.58fF
C7721 vcm_commonmode a_35346_68218# 0.31fF
C7722 a_26402_71230# a_26402_70226# 1.00fF
C7723 a_38450_19532# a_39454_19532# 0.97fF
C7724 a_48490_23548# a_48490_22544# 1.00fF
C7725 a_18979_30287# a_33694_30761# 0.45fF
C7726 a_3280_70501# VDD 0.82fF
C7727 a_42466_66210# a_42466_65206# 1.00fF
C7728 a_43470_14512# a_44474_14512# 0.97fF
C7729 a_25263_38825# VDD 0.61fF
C7730 vcm_commonmode a_38450_21540# 0.87fF
C7731 a_39299_48783# a_44474_72234# 0.35fF
C7732 a_17712_7638# a_17366_15516# 0.38fF
C7733 a_22386_20536# a_23390_20536# 0.97fF
C7734 a_43269_29967# a_47486_13508# 0.38fF
C7735 a_40675_27791# a_41462_15516# 0.38fF
C7736 a_40366_8854# a_40458_8488# 0.32fF
C7737 a_7187_23439# VDD 2.08fF
C7738 a_1923_54591# a_8453_51727# 0.37fF
C7739 a_11619_3303# a_12985_7663# 0.51fF
C7740 a_10515_23975# a_16362_23548# 1.27fF
C7741 a_1591_66415# VDD 0.37fF
C7742 vcm_commonmode a_43470_17524# 0.87fF
C7743 ctopn a_20378_14512# 3.59fF
C7744 a_12663_40871# a_12641_42036# 0.56fF
C7745 vcm_commonmode a_30418_60186# 0.87fF
C7746 a_10791_15529# a_10995_14333# 0.34fF
C7747 a_42466_13508# VDD 0.51fF
C7748 a_41370_70226# a_41462_70226# 0.32fF
C7749 a_10791_57711# a_2419_48783# 0.63fF
C7750 a_13669_37429# a_25133_37571# 0.66fF
C7751 a_1923_73087# a_2971_73493# 0.34fF
C7752 a_10275_21495# a_7377_18012# 0.59fF
C7753 a_7523_62581# VDD 0.46fF
C7754 a_40458_62194# a_40458_61190# 1.00fF
C7755 a_31422_10496# a_31422_9492# 1.00fF
C7756 a_28410_56170# VDD 0.52fF
C7757 vcm_commonmode a_49402_13874# 0.30fF
C7758 a_4528_26159# a_7111_22351# 0.46fF
C7759 a_9955_20969# a_11069_23983# 0.46fF
C7760 a_13097_35279# VDD 1.28fF
C7761 vcm_commonmode a_12895_13967# 6.32fF
C7762 a_18151_52263# a_8295_47388# 2.26fF
C7763 a_22294_16886# a_22386_16520# 0.32fF
C7764 vcm_commonmode a_35346_56170# 0.31fF
C7765 ctopn a_25398_23548# 3.40fF
C7766 a_40458_20536# a_40458_19532# 1.00fF
C7767 vcm_commonmode a_18278_8854# 0.31fF
C7768 a_48490_23548# a_49494_23548# 0.97fF
C7769 a_29927_29199# a_30788_28487# 0.38fF
C7770 a_19807_28111# a_23736_7638# 0.31fF
C7771 a_21382_57174# ctopp 3.58fF
C7772 a_45478_66210# a_46482_66210# 0.97fF
C7773 ctopn a_34434_19532# 3.59fF
C7774 vcm_commonmode m3_16264_22406# 3.20fF
C7775 a_2606_41079# a_3949_41935# 1.06fF
C7776 a_29513_42333# VDD 0.88fF
C7777 a_22015_50645# a_22181_50645# 0.75fF
C7778 a_20378_21540# a_20378_20536# 1.00fF
C7779 a_27406_61190# VDD 0.51fF
C7780 a_7479_54439# a_23929_47381# 0.70fF
C7781 vcm_commonmode a_20378_11500# 0.87fF
C7782 a_22386_12504# a_23390_12504# 0.97fF
C7783 a_36890_34191# VDD 0.37fF
C7784 vcm_commonmode a_44474_18528# 0.87fF
C7785 vcm_commonmode a_34342_61190# 0.31fF
C7786 a_28318_67214# a_28410_67214# 0.32fF
C7787 vcm_commonmode a_24394_24552# 0.84fF
C7788 a_45478_71230# a_45478_70226# 1.00fF
C7789 a_22015_28111# a_9529_28335# 0.51fF
C7790 a_22577_29111# VDD 0.62fF
C7791 a_35438_62194# ctopp 3.59fF
C7792 a_49494_65206# m3_49396_65118# 2.78fF
C7793 a_31422_70226# VDD 0.51fF
C7794 vcm_commonmode a_34434_55166# 0.84fF
C7795 a_8583_33551# a_1761_32143# 0.78fF
C7796 a_25355_40183# VDD 0.64fF
C7797 vcm_commonmode a_26402_57174# 0.87fF
C7798 a_3911_16065# VDD 0.48fF
C7799 a_43267_31055# a_12901_66665# 0.40fF
C7800 vcm_commonmode a_38358_70226# 0.31fF
C7801 a_41462_20536# a_42466_20536# 0.97fF
C7802 a_43175_28335# a_46482_14512# 0.38fF
C7803 a_11251_59879# VDD 8.26fF
C7804 a_30418_63198# a_31422_63198# 0.97fF
C7805 vcm_commonmode a_19282_16886# 0.31fF
C7806 a_13067_38517# a_12663_39783# 3.93fF
C7807 a_41462_71230# ctopp 3.40fF
C7808 ctopn a_37446_20536# 3.59fF
C7809 a_16152_43677# VDD 2.75fF
C7810 a_18151_52263# a_14646_29423# 0.84fF
C7811 a_30326_58178# a_30418_58178# 0.32fF
C7812 a_13123_38231# a_14258_34191# 0.36fF
C7813 a_28423_52245# VDD 0.38fF
C7814 a_17366_21540# a_18370_21540# 0.97fF
C7815 a_20359_29199# a_9135_27239# 3.13fF
C7816 a_25306_9858# a_25398_9492# 0.32fF
C7817 a_22026_27497# VDD 0.83fF
C7818 a_11141_55535# VDD 0.37fF
C7819 a_5167_68060# VDD 0.46fF
C7820 a_33155_35839# VDD 1.25fF
C7821 a_49494_8488# VDD 1.18fF
C7822 vcm_commonmode a_40458_62194# 0.87fF
C7823 a_41370_16886# a_41462_16520# 0.32fF
C7824 a_22015_28111# a_29927_29199# 0.92fF
C7825 a_19807_28111# a_22291_29415# 0.85fF
C7826 a_20378_58178# VDD 0.51fF
C7827 a_24394_59182# a_25398_59182# 0.97fF
C7828 a_3983_20719# VDD 0.41fF
C7829 vcm_commonmode a_48490_15516# 0.87fF
C7830 ctopn a_37446_12504# 3.59fF
C7831 vcm_commonmode a_27314_58178# 0.31fF
C7832 a_41261_28335# a_12901_58799# 0.40fF
C7833 a_22386_17524# a_23390_17524# 0.97fF
C7834 a_42709_29199# a_48490_7484# 0.35fF
C7835 a_35346_72234# a_35438_72234# 0.32fF
C7836 vcm_commonmode a_46482_71230# 0.86fF
C7837 a_39454_21540# a_39454_20536# 1.00fF
C7838 a_12341_3311# a_12985_16367# 0.41fF
C7839 a_7059_24135# VDD 0.94fF
C7840 a_9503_26151# a_20378_22544# 0.38fF
C7841 a_26402_24552# a_26402_23548# 1.00fF
C7842 a_37446_67214# VDD 0.51fF
C7843 a_41462_12504# a_42466_12504# 0.97fF
C7844 a_19720_55394# a_12981_59343# 0.40fF
C7845 a_47394_67214# a_47486_67214# 0.32fF
C7846 ctopn a_32426_21540# 3.59fF
C7847 vcm_commonmode a_44382_67214# 0.31fF
C7848 vcm_commonmode a_25398_13508# 0.87fF
C7849 a_13576_37149# VDD 2.26fF
C7850 a_44474_68218# ctopp 3.59fF
C7851 ctopn a_37446_17524# 3.59fF
C7852 a_12725_44527# a_1803_20719# 0.63fF
C7853 a_22132_44129# a_23567_44211# 0.87fF
C7854 a_34434_9492# VDD 0.51fF
C7855 a_40050_48463# a_12355_15055# 0.40fF
C7856 a_25787_28327# a_12516_7093# 0.40fF
C7857 a_33338_7850# a_33430_7484# 0.32fF
C7858 vcm_commonmode a_41370_9858# 0.31fF
C7859 m3_49396_64114# VDD 0.35fF
C7860 a_12231_65301# VDD 0.40fF
C7861 a_47486_24552# m3_47388_24414# 2.81fF
C7862 a_42374_72234# VDD 0.61fF
C7863 a_2952_66139# a_3938_61493# 0.62fF
C7864 vcm_commonmode a_21290_22910# 0.31fF
C7865 a_7000_43541# a_8383_43255# 0.48fF
C7866 a_17274_69222# a_17366_69222# 0.32fF
C7867 a_23390_18528# a_23390_17524# 1.00fF
C7868 a_43269_29967# a_47486_7484# 0.34fF
C7869 a_17039_51157# a_14831_50095# 1.45fF
C7870 a_36442_21540# a_37446_21540# 0.97fF
C7871 a_2775_46025# VDD 14.94fF
C7872 a_44382_9858# a_44474_9492# 0.32fF
C7873 a_12394_25615# VDD 0.57fF
C7874 a_11067_13095# a_1586_18695# 0.72fF
C7875 a_23736_7638# a_12985_19087# 0.41fF
C7876 a_27314_64202# a_27406_64202# 0.32fF
C7877 a_42466_7484# VDD 1.36fF
C7878 a_16746_67216# a_16362_67214# 2.28fF
C7879 a_8566_39215# VDD 1.38fF
C7880 vcm_commonmode a_49494_68218# 0.91fF
C7881 a_43470_59182# a_44474_59182# 0.97fF
C7882 a_19478_51959# a_25419_50959# 1.24fF
C7883 a_35601_27497# a_35438_19532# 0.38fF
C7884 a_24302_22910# a_24394_22544# 0.32fF
C7885 a_36442_64202# VDD 0.51fF
C7886 a_31117_28879# VDD 0.50fF
C7887 a_7479_57175# VDD 0.30fF
C7888 vcm_commonmode a_17274_14878# 0.33fF
C7889 a_44474_56170# ctopp 3.40fF
C7890 a_43362_28879# a_47486_59182# 0.38fF
C7891 a_12355_65103# a_12355_15055# 2.05fF
C7892 a_24394_14512# a_24394_13508# 1.00fF
C7893 a_5691_36727# VDD 1.83fF
C7894 ctopn a_38450_18528# 3.59fF
C7895 a_19919_38695# VDD 1.49fF
C7896 vcm_commonmode a_43378_64202# 0.31fF
C7897 a_41462_17524# a_42466_17524# 0.97fF
C7898 ctopn a_18370_24552# 0.57fF
C7899 a_3247_20495# a_5825_20495# 0.86fF
C7900 a_1761_30511# a_1867_32839# 0.42fF
C7901 a_27535_30503# a_20635_29415# 0.43fF
C7902 a_18611_52047# a_23390_71230# 0.38fF
C7903 a_28756_7638# a_28410_14512# 0.38fF
C7904 a_28410_60186# a_29414_60186# 0.97fF
C7905 a_45478_24552# a_45478_23548# 1.00fF
C7906 a_7213_62215# VDD 1.31fF
C7907 a_12357_37999# a_15305_38543# 0.54fF
C7908 a_6835_46823# a_7050_53333# 0.34fF
C7909 a_30418_12504# a_30418_11500# 1.00fF
C7910 a_6327_72917# VDD 1.03fF
C7911 a_34780_56398# a_34434_61190# 0.38fF
C7912 vcm_commonmode a_22294_23914# 0.31fF
C7913 a_20378_7484# m3_20280_7346# 2.80fF
C7914 a_20839_44265# VDD 0.58fF
C7915 a_17599_52263# a_22386_67214# 0.38fF
C7916 a_17366_70226# a_17366_69222# 1.00fF
C7917 vcm_commonmode a_19282_66210# 0.31fF
C7918 a_23390_18528# a_24394_18528# 0.97fF
C7919 a_24394_19532# VDD 0.51fF
C7920 a_35550_27791# VDD 0.33fF
C7921 a_43470_61190# ctopp 3.59fF
C7922 ctopn a_47486_10496# 3.58fF
C7923 a_45478_69222# VDD 0.51fF
C7924 a_12381_35836# VDD 7.51fF
C7925 vcm_commonmode a_31330_19898# 0.31fF
C7926 a_42985_46831# a_48490_64202# 0.38fF
C7927 vcm_commonmode a_16362_62194# 4.47fF
C7928 vcm_commonmode a_49494_56170# 0.90fF
C7929 a_39299_48783# a_12257_56623# 0.40fF
C7930 vcm_commonmode a_32426_8488# 0.86fF
C7931 m3_49396_11362# VDD 0.34fF
C7932 a_36797_27497# a_37446_20536# 0.38fF
C7933 a_43470_65206# VDD 0.51fF
C7934 a_11803_55311# VDD 7.61fF
C7935 ctopp inp_analog 1.03fF
C7936 a_39389_52271# a_10515_22671# 0.40fF
C7937 a_1768_13103# config_1_in[12] 1.32fF
C7938 a_20286_14878# a_20378_14512# 0.32fF
C7939 a_12985_19087# a_16362_8488# 19.89fF
C7940 a_11067_67279# a_26748_7638# 0.41fF
C7941 a_47486_70226# ctopp 3.57fF
C7942 a_15009_40193# VDD 1.39fF
C7943 a_36350_69222# a_36442_69222# 0.32fF
C7944 a_43470_59182# a_43470_58178# 1.00fF
C7945 a_42466_18528# a_42466_17524# 1.00fF
C7946 VDD config_2_in[13] 0.98fF
C7947 a_16362_8488# a_16746_8486# 2.28fF
C7948 a_32334_24918# VDD 0.36fF
C7949 a_11711_67325# VDD 0.39fF
C7950 a_46390_64202# a_46482_64202# 0.32fF
C7951 ctopn a_42466_15516# 3.59fF
C7952 a_12663_40871# a_12889_40977# 0.60fF
C7953 vcm_commonmode a_48490_61190# 0.87fF
C7954 a_22291_29415# a_29927_29199# 0.48fF
C7955 a_48490_14512# VDD 0.54fF
C7956 a_2927_39733# VDD 1.17fF
C7957 vcm_commonmode a_20378_67214# 0.87fF
C7958 a_36797_27497# a_37446_12504# 0.38fF
C7959 a_27406_20536# VDD 0.51fF
C7960 a_42374_55166# VDD 0.35fF
C7961 a_12341_3311# a_22386_19532# 0.38fF
C7962 a_33864_28111# a_34434_18528# 0.38fF
C7963 a_43378_22910# a_43470_22544# 0.32fF
C7964 a_12981_62313# VDD 7.11fF
C7965 a_7295_44647# a_34759_31029# 0.33fF
C7966 a_32426_10496# a_33430_10496# 0.97fF
C7967 a_31768_55394# a_31422_58178# 0.38fF
C7968 a_34342_65206# a_34434_65206# 0.32fF
C7969 a_43470_14512# a_43470_13508# 1.00fF
C7970 vcm_commonmode a_34342_20902# 0.31fF
C7971 a_12725_44527# a_14258_44527# 1.20fF
C7972 a_7187_37583# VDD 0.52fF
C7973 vcm_commonmode a_23298_63198# 0.31fF
C7974 a_17039_51157# a_21261_47919# 0.64fF
C7975 a_23830_49525# a_23774_49551# 0.96fF
C7976 a_39454_72234# a_39454_71230# 1.00fF
C7977 a_1761_25071# a_2315_24540# 0.92fF
C7978 a_47486_60186# a_48490_60186# 0.97fF
C7979 vcm_commonmode a_17366_9492# 1.82fF
C7980 a_36442_58178# ctopp 3.59fF
C7981 a_25306_23914# a_25398_23548# 0.32fF
C7982 a_4443_46607# a_17672_32259# 0.61fF
C7983 a_33430_56170# a_33430_55166# 1.00fF
C7984 a_49494_12504# a_49494_11500# 1.00fF
C7985 a_18370_11500# a_19374_11500# 0.97fF
C7986 a_17358_31069# VDD 2.23fF
C7987 vcm_commonmode a_33430_16520# 0.87fF
C7988 a_12355_15055# ctopp 3.23fF
C7989 ctopn a_19374_13508# 3.59fF
C7990 a_12899_3855# a_11619_3303# 0.58fF
C7991 a_24394_72234# VDD 1.24fF
C7992 a_23395_52047# a_12727_58255# 0.40fF
C7993 a_22294_66210# a_22386_66210# 0.32fF
C7994 vcm_commonmode a_17274_59182# 0.33fF
C7995 a_27406_12504# VDD 0.51fF
C7996 a_4351_67279# a_3024_67191# 0.87fF
C7997 a_36442_70226# a_36442_69222# 1.00fF
C7998 a_42466_18528# a_43470_18528# 0.97fF
C7999 a_2411_18517# VDD 5.02fF
C8000 a_20535_51727# VDD 0.40fF
C8001 a_6453_71855# a_5023_72068# 0.53fF
C8002 vcm_commonmode a_29414_72234# 0.69fF
C8003 a_36797_27497# a_37446_17524# 0.38fF
C8004 a_22291_29415# a_28817_29111# 0.30fF
C8005 a_13643_28327# a_33864_28111# 0.58fF
C8006 vcm_commonmode a_34342_12870# 0.31fF
C8007 a_16746_60188# ctopp 1.68fF
C8008 a_22386_24552# a_23390_24552# 0.97fF
C8009 a_43362_28879# a_47486_57174# 0.38fF
C8010 a_34342_19898# a_34434_19532# 0.32fF
C8011 a_6559_59663# a_8491_57487# 0.74fF
C8012 a_22386_21540# VDD 0.51fF
C8013 vcm_commonmode a_25398_7484# 0.69fF
C8014 a_7676_61493# VDD 1.05fF
C8015 a_12907_27023# a_43680_29941# 0.44fF
C8016 a_16863_29415# a_30565_30199# 1.09fF
C8017 a_19374_62194# a_20378_62194# 0.97fF
C8018 a_35438_11500# a_35438_10496# 1.00fF
C8019 a_14287_51175# a_8491_57487# 0.59fF
C8020 a_39362_14878# a_39454_14512# 0.32fF
C8021 vcm_commonmode a_29322_21906# 0.31fF
C8022 a_23390_69222# ctopp 3.59fF
C8023 a_14646_29423# a_18829_29423# 0.33fF
C8024 a_44474_72234# m3_44376_72146# 2.80fF
C8025 a_10259_10703# VDD 0.38fF
C8026 vcm_commonmode a_19374_64202# 0.87fF
C8027 a_39673_28111# a_40458_8488# 0.38fF
C8028 vcm_commonmode a_47394_58178# 0.31fF
C8029 a_31223_36369# a_13669_35253# 0.33fF
C8030 a_27406_17524# VDD 0.51fF
C8031 a_36629_27791# a_36442_15516# 0.38fF
C8032 a_18278_20902# a_18370_20536# 0.32fF
C8033 a_49494_19532# m3_49396_19394# 2.78fF
C8034 a_33338_55166# a_33430_55166# 0.33fF
C8035 a_1803_20719# a_2012_33927# 1.32fF
C8036 a_30788_28487# VDD 3.14fF
C8037 vcm_commonmode a_34342_17890# 0.31fF
C8038 a_21382_65206# ctopp 3.59fF
C8039 a_24394_57174# a_25398_57174# 0.97fF
C8040 a_3275_73658# VDD 0.52fF
C8041 vcm_commonmode a_21290_60186# 0.31fF
C8042 a_27406_15516# a_28410_15516# 0.97fF
C8043 a_33856_44869# VDD 1.51fF
C8044 a_6008_69679# a_5924_69135# 0.36fF
C8045 a_10515_63143# a_7000_43541# 0.47fF
C8046 a_4427_25071# VDD 1.54fF
C8047 a_3339_30503# a_17712_7638# 0.83fF
C8048 a_2952_66139# a_6515_62037# 0.45fF
C8049 a_5915_30287# a_14097_31375# 1.05fF
C8050 a_6895_15253# VDD 0.36fF
C8051 a_25398_71230# a_26402_71230# 0.97fF
C8052 vcm_commonmode a_28410_69222# 0.87fF
C8053 a_11067_13095# a_6372_38279# 1.33fF
C8054 a_48490_59182# VDD 0.55fF
C8055 a_43470_58178# a_43470_57174# 1.00fF
C8056 a_44382_23914# a_44474_23548# 0.32fF
C8057 a_40675_27791# a_41462_20536# 0.38fF
C8058 a_17712_7638# a_17366_20536# 0.38fF
C8059 a_37446_11500# a_38450_11500# 0.97fF
C8060 a_15681_27497# a_12349_25847# 0.72fF
C8061 a_41370_66210# a_41462_66210# 0.32fF
C8062 vcm_commonmode a_35438_22544# 0.87fF
C8063 a_28446_31375# a_32823_29397# 0.37fF
C8064 vcm_commonmode a_26402_65206# 0.87fF
C8065 a_39299_48783# a_10975_66407# 0.40fF
C8066 a_28410_18528# VDD 0.51fF
C8067 a_19894_51433# VDD 0.44fF
C8068 a_17712_7638# a_12727_13353# 0.40fF
C8069 ctopn a_26402_8488# 3.40fF
C8070 a_41462_24552# a_42466_24552# 0.97fF
C8071 a_18278_12870# a_18370_12504# 0.32fF
C8072 vcm_commonmode a_35346_18894# 0.31fF
C8073 a_28410_66210# ctopp 3.59fF
C8074 a_18611_52047# a_4215_51157# 1.55fF
C8075 a_1586_18695# a_10883_11177# 0.41fF
C8076 a_6224_73095# a_5254_67503# 0.73fF
C8077 a_42709_29199# a_48490_11500# 0.38fF
C8078 a_17712_7638# a_17366_12504# 0.38fF
C8079 a_40675_27791# a_41462_12504# 0.38fF
C8080 a_19374_55166# VDD 0.60fF
C8081 a_23736_7638# a_23390_15516# 0.38fF
C8082 a_38450_62194# a_39454_62194# 0.97fF
C8083 a_4151_28879# VDD 0.55fF
C8084 vcm_commonmode a_31422_14512# 0.87fF
C8085 a_11067_63143# a_11480_23957# 1.01fF
C8086 vcm_commonmode a_26310_55166# 0.30fF
C8087 a_37446_10496# VDD 0.51fF
C8088 a_4685_37583# VDD 3.40fF
C8089 vcm_commonmode a_17274_57174# 0.33fF
C8090 a_12621_36091# a_20715_34717# 0.74fF
C8091 a_4495_35925# a_7695_31573# 0.35fF
C8092 a_22015_28111# VDD 10.48fF
C8093 a_39389_52271# a_12901_66665# 0.40fF
C8094 a_37354_20902# a_37446_20536# 0.32fF
C8095 a_3339_43023# a_7571_29199# 1.30fF
C8096 a_7210_55081# a_4674_57685# 0.96fF
C8097 vcm_commonmode a_44382_10862# 0.31fF
C8098 a_26310_63198# a_26402_63198# 0.32fF
C8099 a_12263_4391# a_25744_7638# 1.29fF
C8100 a_1803_20719# a_2052_38377# 0.61fF
C8101 a_43470_57174# a_44474_57174# 0.97fF
C8102 a_17366_57174# a_17366_56170# 1.00fF
C8103 a_13183_52047# a_17366_60186# 0.38fF
C8104 a_46482_15516# a_47486_15516# 0.97fF
C8105 vcm_commonmode a_36442_23548# 0.87fF
C8106 a_11067_67279# a_43269_29967# 0.41fF
C8107 vcm_commonmode a_33430_66210# 0.87fF
C8108 a_2775_46025# a_4057_50645# 0.58fF
C8109 a_35601_27497# a_12877_16911# 0.41fF
C8110 a_17712_7638# a_17366_17524# 0.38fF
C8111 a_40675_27791# a_41462_17524# 0.38fF
C8112 a_24394_62194# VDD 0.51fF
C8113 a_17712_7638# a_10515_23975# 0.40fF
C8114 vcm_commonmode a_45478_19532# 0.87fF
C8115 ctopn a_27406_16520# 3.59fF
C8116 vcm_commonmode a_31330_62194# 0.31fF
C8117 a_32426_15516# VDD 0.51fF
C8118 a_37557_32463# VDD 3.34fF
C8119 a_1923_73087# a_3024_67191# 0.38fF
C8120 a_44474_71230# a_45478_71230# 0.97fF
C8121 a_43270_27791# a_45478_13508# 0.38fF
C8122 a_43269_29967# a_47486_11500# 0.38fF
C8123 a_10957_57711# VDD 0.41fF
C8124 a_20286_59182# a_20378_59182# 0.32fF
C8125 a_10275_21495# VDD 0.49fF
C8126 a_39673_28111# a_12985_19087# 0.41fF
C8127 a_31768_7638# a_12899_10927# 0.41fF
C8128 a_24740_7638# a_24394_19532# 0.38fF
C8129 a_24959_30503# a_14926_31849# 0.76fF
C8130 vcm_commonmode a_39362_15882# 0.31fF
C8131 a_32426_63198# ctopp 3.64fF
C8132 a_30418_71230# VDD 0.58fF
C8133 a_34251_52263# a_12901_58799# 0.40fF
C8134 a_27379_39095# VDD 0.65fF
C8135 a_1689_10396# a_1929_10651# 0.76fF
C8136 a_42466_11500# VDD 0.51fF
C8137 a_33764_41831# VDD 1.61fF
C8138 a_18278_17890# a_18370_17524# 0.32fF
C8139 a_22015_50645# VDD 0.46fF
C8140 vcm_commonmode a_37354_71230# 0.31fF
C8141 a_5363_30503# a_9367_29397# 0.38fF
C8142 a_46482_24552# VDD 0.60fF
C8143 vcm_commonmode a_49402_11866# 0.30fF
C8144 a_26402_59182# ctopp 3.59fF
C8145 a_28756_7638# a_12985_7663# 0.41fF
C8146 a_24394_64202# a_24394_63198# 1.23fF
C8147 a_37354_12870# a_37446_12504# 0.32fF
C8148 a_19439_32143# VDD 0.30fF
C8149 a_5024_67885# a_8896_65015# 0.37fF
C8150 a_10515_63143# a_5915_35943# 1.18fF
C8151 a_32426_59182# a_32426_58178# 1.00fF
C8152 a_2959_47113# a_27793_51733# 0.53fF
C8153 a_11067_21583# a_16362_21540# 19.89fF
C8154 a_30764_7638# a_12899_10927# 0.41fF
C8155 a_12447_29199# a_32970_31145# 1.10fF
C8156 a_11067_46823# a_28305_28879# 0.39fF
C8157 a_48490_57174# VDD 0.54fF
C8158 a_23390_13508# a_24394_13508# 0.97fF
C8159 vcm_commonmode a_48490_20536# 0.87fF
C8160 a_32795_39679# VDD 0.99fF
C8161 a_38557_32143# a_12355_15055# 0.40fF
C8162 a_28410_68218# a_29414_68218# 0.97fF
C8163 vcm_commonmode a_37446_63198# 0.92fF
C8164 a_2292_17179# a_1591_14741# 0.36fF
C8165 a_13183_52047# a_12257_56623# 0.40fF
C8166 a_21371_52263# a_12516_7093# 0.47fF
C8167 a_4482_57863# a_26397_51183# 0.43fF
C8168 a_8671_22671# VDD 0.41fF
C8169 a_10055_58791# a_11067_21583# 0.72fF
C8170 m3_37348_72146# VDD 0.41fF
C8171 a_42718_27497# a_44474_21540# 0.38fF
C8172 a_39223_32463# a_39454_16520# 0.38fF
C8173 a_34482_29941# a_30788_28487# 0.43fF
C8174 a_20635_29415# a_25313_31599# 1.04fF
C8175 a_40458_56170# a_40458_55166# 1.00fF
C8176 a_40458_24552# m3_40360_24414# 2.81fF
C8177 a_45386_63198# a_45478_63198# 0.32fF
C8178 a_23736_7638# VDD 8.91fF
C8179 a_8132_53511# a_7749_55535# 0.31fF
C8180 a_36442_57174# a_36442_56170# 1.00fF
C8181 a_35346_72234# VDD 0.61fF
C8182 vcm_commonmode a_31422_59182# 0.87fF
C8183 a_3339_30503# a_4248_29967# 0.68fF
C8184 a_23763_47381# a_23929_47381# 0.46fF
C8185 a_19559_43177# VDD 0.60fF
C8186 a_32612_51727# VDD 0.67fF
C8187 a_32334_21906# a_32426_21540# 0.32fF
C8188 a_1775_60663# VDD 0.81fF
C8189 vcm_commonmode a_48490_12504# 0.87fF
C8190 a_30418_60186# ctopp 3.59fF
C8191 a_33430_68218# VDD 0.51fF
C8192 a_33338_7850# VDD 0.63fF
C8193 a_20378_16520# a_20378_15516# 1.00fF
C8194 ctopn a_29414_22544# 3.58fF
C8195 vcm_commonmode a_40366_68218# 0.31fF
C8196 a_2143_15271# a_5320_18231# 0.30fF
C8197 a_39362_59182# a_39454_59182# 0.32fF
C8198 a_6835_46823# a_14831_50095# 0.30fF
C8199 a_19459_29423# VDD 0.34fF
C8200 a_7097_40303# a_6372_38279# 0.33fF
C8201 a_15189_39889# a_14963_39783# 0.32fF
C8202 a_41872_29423# a_43470_59182# 0.38fF
C8203 vcm_commonmode a_43470_21540# 0.87fF
C8204 a_37354_17890# a_37446_17524# 0.32fF
C8205 a_25744_7638# a_25398_8488# 0.38fF
C8206 a_8491_27023# a_18370_8488# 0.38fF
C8207 a_2292_43291# VDD 4.17fF
C8208 a_19720_55394# a_19374_71230# 0.38fF
C8209 a_4482_57863# a_25419_50959# 0.52fF
C8210 a_24302_60186# a_24394_60186# 0.32fF
C8211 vcm_commonmode a_20378_10496# 0.87fF
C8212 a_43470_64202# a_43470_63198# 1.23fF
C8213 a_3668_56311# a_4298_58951# 0.39fF
C8214 a_10515_22671# a_4903_31849# 0.59fF
C8215 vcm_commonmode a_48490_17524# 0.87fF
C8216 a_11067_67279# a_7377_18012# 0.68fF
C8217 ctopn a_25398_14512# 3.59fF
C8218 a_2191_68565# a_3325_49551# 0.40fF
C8219 a_4351_67279# a_6775_53877# 0.93fF
C8220 a_12473_42869# a_12473_41781# 1.56fF
C8221 a_4227_73791# VDD 0.48fF
C8222 vcm_commonmode a_35438_60186# 0.87fF
C8223 a_25971_52263# a_30418_61190# 0.38fF
C8224 a_47486_13508# VDD 0.51fF
C8225 a_14287_51175# a_18370_67214# 0.38fF
C8226 a_19282_18894# a_19374_18528# 0.32fF
C8227 a_10961_19087# VDD 0.62fF
C8228 a_1761_25071# config_1_in[15] 0.42fF
C8229 a_35438_22544# a_35438_21540# 1.00fF
C8230 a_6835_46823# a_19333_48463# 0.40fF
C8231 a_33430_56170# VDD 0.52fF
C8232 a_42466_13508# a_43470_13508# 0.97fF
C8233 a_24055_36415# VDD 1.09fF
C8234 a_16362_8488# VDD 2.54fF
C8235 a_39299_48783# a_44474_64202# 0.38fF
C8236 a_47486_68218# a_48490_68218# 0.97fF
C8237 vcm_commonmode a_40366_56170# 0.31fF
C8238 a_36613_48169# a_12257_56623# 0.40fF
C8239 ctopn a_30418_23548# 3.40fF
C8240 a_19807_28111# a_12907_27023# 1.44fF
C8241 a_22291_29415# VDD 14.64fF
C8242 a_39454_58178# a_39389_52271# 0.38fF
C8243 vcm_commonmode a_23298_8854# 0.31fF
C8244 ctopp a_34434_55166# 0.65fF
C8245 a_1823_62589# a_3016_60949# 0.64fF
C8246 a_28410_56170# a_29414_56170# 0.97fF
C8247 a_26402_57174# ctopp 3.58fF
C8248 a_28547_51175# a_10515_22671# 0.40fF
C8249 ctopn a_39454_19532# 3.59fF
C8250 a_14625_30761# a_13353_30511# 0.89fF
C8251 a_8197_31599# a_6459_30511# 1.26fF
C8252 a_22386_72234# a_23390_72234# 0.97fF
C8253 a_1768_13103# a_1586_36727# 0.66fF
C8254 a_32426_61190# VDD 0.51fF
C8255 vcm_commonmode a_25398_11500# 0.87fF
C8256 a_32426_58178# a_32426_57174# 1.00fF
C8257 a_12355_15055# a_10515_63143# 0.69fF
C8258 vcm_commonmode a_49494_18528# 1.01fF
C8259 a_31768_55394# a_28881_52271# 0.95fF
C8260 vcm_commonmode a_39362_61190# 0.31fF
C8261 a_39454_16520# a_39454_15516# 1.00fF
C8262 vcm_commonmode a_29414_24552# 0.84fF
C8263 a_24394_19532# a_24394_18528# 1.00fF
C8264 a_33338_55166# VDD 0.36fF
C8265 a_2959_47113# a_19478_51959# 0.38fF
C8266 a_28318_10862# a_28410_10496# 0.32fF
C8267 a_40458_62194# ctopp 3.59fF
C8268 a_1761_40847# a_12641_37684# 0.31fF
C8269 a_36442_70226# VDD 0.51fF
C8270 a_23395_52047# a_27406_58178# 0.38fF
C8271 vcm_commonmode a_39454_55166# 0.84fF
C8272 a_31084_30485# a_30565_30199# 0.30fF
C8273 a_30788_28487# a_36904_28879# 0.46fF
C8274 a_43362_28879# a_47486_65206# 0.38fF
C8275 a_43270_27791# a_45478_7484# 0.34fF
C8276 vcm_commonmode a_31422_57174# 0.87fF
C8277 a_17366_16520# VDD 0.58fF
C8278 a_7557_49007# VDD 0.41fF
C8279 vcm_commonmode a_43378_70226# 0.31fF
C8280 a_35438_72234# a_35438_71230# 1.00fF
C8281 a_5190_59575# VDD 5.05fF
C8282 a_43378_60186# a_43470_60186# 0.32fF
C8283 VDD dummypin[12] 0.79fF
C8284 vcm_commonmode a_24302_16886# 0.31fF
C8285 a_17366_72234# VDD 1.61fF
C8286 a_1761_52815# a_37733_37477# 0.62fF
C8287 a_16955_52047# a_12727_58255# 0.40fF
C8288 a_19374_15516# a_19374_14512# 1.00fF
C8289 a_46482_71230# ctopp 3.40fF
C8290 ctopn a_42466_20536# 3.59fF
C8291 a_5039_42167# a_2021_17973# 0.32fF
C8292 a_42985_46831# a_12983_63151# 0.40fF
C8293 a_13183_52047# a_10975_66407# 0.40fF
C8294 a_38358_18894# a_38450_18528# 0.32fF
C8295 vcm_commonmode a_22386_72234# 0.69fF
C8296 a_6095_44807# a_6725_45205# 0.60fF
C8297 a_22291_29415# a_18053_28879# 0.66fF
C8298 a_22015_28111# a_24740_7638# 1.84fF
C8299 a_27406_61190# a_28410_61190# 0.97fF
C8300 a_1644_54965# VDD 0.31fF
C8301 a_18278_24918# a_18370_24552# 0.33fF
C8302 a_31768_7638# a_31422_22544# 0.38fF
C8303 a_8675_68047# VDD 0.47fF
C8304 a_1887_34863# VDD 0.37fF
C8305 vcm_commonmode a_45478_62194# 0.87fF
C8306 a_33430_68218# a_33430_67214# 1.00fF
C8307 a_4119_70741# a_3016_60949# 0.33fF
C8308 a_41872_29423# a_43470_57174# 0.38fF
C8309 a_42985_46831# a_48490_70226# 0.38fF
C8310 vcm_commonmode a_12727_67753# 6.23fF
C8311 a_25398_58178# VDD 0.51fF
C8312 vcm_commonmode a_16270_7850# 0.33fF
C8313 a_8491_41383# a_13357_32143# 0.35fF
C8314 ctopn a_42466_12504# 3.59fF
C8315 a_34251_52263# a_18703_29199# 0.40fF
C8316 a_4314_40821# a_6372_38279# 0.44fF
C8317 a_47486_56170# a_48490_56170# 0.97fF
C8318 vcm_commonmode a_32334_58178# 0.31fF
C8319 a_12985_16367# a_16746_11498# 2.28fF
C8320 a_3607_34639# a_7461_27247# 0.53fF
C8321 a_7373_40847# VDD 1.13fF
C8322 a_18370_69222# a_18370_68218# 1.00fF
C8323 VDD config_2_in[3] 2.16fF
C8324 a_36613_48169# a_37446_72234# 0.34fF
C8325 a_29322_55166# a_29414_55166# 0.32fF
C8326 a_30418_8488# a_31422_8488# 0.97fF
C8327 a_42466_67214# VDD 0.51fF
C8328 a_13643_28327# a_3339_30503# 0.39fF
C8329 ctopp m3_18272_55078# 0.35fF
C8330 a_1586_21959# a_3972_25615# 0.38fF
C8331 a_20286_57174# a_20378_57174# 0.32fF
C8332 a_1586_69367# VDD 7.48fF
C8333 a_23298_15882# a_23390_15516# 0.32fF
C8334 ctopn a_37446_21540# 3.59fF
C8335 a_2012_33927# a_3325_18543# 0.45fF
C8336 a_31422_70226# a_32426_70226# 0.97fF
C8337 vcm_commonmode a_49402_67214# 0.30fF
C8338 a_43470_19532# a_43470_18528# 1.00fF
C8339 a_77451_38925# inp_analog 0.44fF
C8340 a_1770_14441# a_1586_36727# 0.47fF
C8341 a_12907_27023# a_9529_28335# 0.69fF
C8342 a_47394_10862# a_47486_10496# 0.32fF
C8343 a_3780_56347# VDD 1.87fF
C8344 vcm_commonmode a_30418_13508# 0.87fF
C8345 a_6733_69135# VDD 0.49fF
C8346 a_25484_37253# VDD 1.59fF
C8347 ctopn a_42466_17524# 3.59fF
C8348 m2_48260_54946# m3_48968_55078# 0.62fF
C8349 a_39454_9492# VDD 0.51fF
C8350 a_12546_22351# a_16746_10494# 2.28fF
C8351 vcm_commonmode a_16746_56172# 5.35fF
C8352 a_14287_51175# a_7479_54439# 2.01fF
C8353 vcm_commonmode a_19282_69222# 0.31fF
C8354 a_21290_71230# a_21382_71230# 0.32fF
C8355 a_29414_60186# a_29414_59182# 1.00fF
C8356 a_19374_22544# VDD 0.51fF
C8357 vcm_commonmode a_46390_9858# 0.31fF
C8358 a_36629_27791# a_36442_20536# 0.38fF
C8359 a_18370_63198# a_18370_62194# 1.00fF
C8360 a_33338_11866# a_33430_11500# 0.32fF
C8361 a_11155_30663# VDD 0.43fF
C8362 a_10975_66407# a_12546_22351# 1.07fF
C8363 a_43267_31055# VDD 8.37fF
C8364 a_38450_15516# a_38450_14512# 1.00fF
C8365 vcm_commonmode a_26310_22910# 0.31fF
C8366 a_3339_30503# a_23195_29967# 0.43fF
C8367 a_4674_40277# a_12447_29199# 0.45fF
C8368 a_18979_30287# a_8491_41383# 1.76fF
C8369 vcm_commonmode a_17274_65206# 0.33fF
C8370 a_36613_48169# a_10975_66407# 0.40fF
C8371 a_2872_44111# a_7000_43541# 0.70fF
C8372 a_14859_51183# VDD 0.36fF
C8373 a_46482_61190# a_47486_61190# 0.97fF
C8374 a_23390_9492# a_23390_8488# 1.00fF
C8375 a_37354_24918# a_37446_24552# 0.32fF
C8376 a_9955_20969# a_8933_22583# 0.36fF
C8377 a_11067_13095# a_6773_27805# 0.53fF
C8378 a_23736_7638# a_24740_7638# 0.30fF
C8379 a_47486_7484# VDD 1.23fF
C8380 a_25787_28327# a_6467_55527# 1.03fF
C8381 a_18370_67214# a_19374_67214# 0.97fF
C8382 a_20635_29415# a_7295_44647# 0.76fF
C8383 a_12907_27023# a_29927_29199# 0.30fF
C8384 a_2952_46805# VDD 2.35fF
C8385 a_1591_57711# a_2191_68565# 0.90fF
C8386 a_36629_27791# a_36442_12504# 0.38fF
C8387 a_7050_53333# a_14983_51157# 0.86fF
C8388 a_12869_2741# a_27869_50095# 0.50fF
C8389 a_2959_47113# a_1761_52815# 2.41fF
C8390 a_41462_64202# VDD 0.51fF
C8391 a_34342_62194# a_34434_62194# 0.32fF
C8392 a_2163_56765# VDD 0.47fF
C8393 vcm_commonmode a_22294_14878# 0.31fF
C8394 a_16362_62194# ctopp 1.35fF
C8395 ctopn a_19374_11500# 3.59fF
C8396 a_18045_38017# VDD 1.50fF
C8397 ctopn a_43470_18528# 3.59fF
C8398 a_15851_27791# a_13390_29575# 0.76fF
C8399 a_30943_38695# VDD 1.82fF
C8400 vcm_commonmode a_48398_64202# 0.31fF
C8401 a_37446_69222# a_37446_68218# 1.00fF
C8402 a_4495_35925# a_5595_33205# 0.34fF
C8403 vcm_commonmode a_19374_70226# 0.87fF
C8404 a_28547_51175# a_12901_66665# 0.40fF
C8405 a_47394_55166# a_47486_55166# 0.32fF
C8406 a_27406_8488# a_27406_7484# 1.00fF
C8407 a_20378_23548# VDD 0.52fF
C8408 a_4891_47388# a_10680_52245# 2.38fF
C8409 a_17366_66210# VDD 0.57fF
C8410 a_17366_56170# a_17366_55166# 1.00fF
C8411 a_2317_28892# a_3143_22364# 1.38fF
C8412 a_39362_57174# a_39454_57174# 0.32fF
C8413 a_1770_14441# a_1768_13103# 0.94fF
C8414 a_42374_15882# a_42466_15516# 0.32fF
C8415 vcm_commonmode a_27314_23914# 0.31fF
C8416 a_32795_44031# VDD 1.02fF
C8417 vcm_commonmode a_24302_66210# 0.31fF
C8418 a_20378_58178# a_21382_58178# 0.97fF
C8419 a_29414_19532# VDD 0.51fF
C8420 a_2775_46025# a_26397_51183# 1.61fF
C8421 a_36629_27791# a_36442_17524# 0.38fF
C8422 a_39673_28111# VDD 7.04fF
C8423 a_10055_58791# a_9135_27239# 0.41fF
C8424 a_48490_61190# ctopp 3.43fF
C8425 a_23736_7638# a_23390_20536# 0.38fF
C8426 a_1761_35407# VDD 9.93fF
C8427 vcm_commonmode a_36350_19898# 0.31fF
C8428 a_20378_67214# ctopp 3.59fF
C8429 a_26523_29199# a_12899_3311# 0.35fF
C8430 a_31422_16520# a_32426_16520# 0.97fF
C8431 a_15617_47919# VDD 0.59fF
C8432 a_40366_71230# a_40458_71230# 0.32fF
C8433 a_48490_60186# a_48490_59182# 1.00fF
C8434 vcm_commonmode a_37446_8488# 0.86fF
C8435 a_48490_65206# VDD 0.54fF
C8436 a_12447_29199# a_7862_34025# 1.43fF
C8437 a_37446_63198# a_37446_62194# 1.00fF
C8438 a_40050_48463# a_20635_29415# 0.44fF
C8439 a_4314_40821# a_4259_40847# 0.51fF
C8440 a_28756_55394# a_12901_58799# 0.40fF
C8441 a_13484_39325# VDD 2.59fF
C8442 a_13097_35279# a_12549_35836# 0.38fF
C8443 a_2473_34293# a_1915_35015# 2.12fF
C8444 a_7019_50639# VDD 0.34fF
C8445 a_28318_72234# a_28410_72234# 0.32fF
C8446 a_23736_7638# a_23390_12504# 0.38fF
C8447 a_42466_9492# a_42466_8488# 1.00fF
C8448 a_37354_24918# VDD 0.36fF
C8449 a_7841_12167# inn_analog 0.43fF
C8450 ctopn a_47486_15516# 3.58fF
C8451 a_6559_42479# a_6725_42479# 0.68fF
C8452 a_37446_67214# a_38450_67214# 0.97fF
C8453 a_2473_34293# a_4248_29967# 0.40fF
C8454 vcm_commonmode a_25398_67214# 0.87fF
C8455 a_32426_20536# VDD 0.51fF
C8456 a_47394_55166# VDD 0.35fF
C8457 a_6831_63303# a_2606_41079# 1.09fF
C8458 a_21382_63198# VDD 0.57fF
C8459 a_41261_28335# a_26523_28111# 0.95fF
C8460 a_1761_27791# config_2_in[1] 0.35fF
C8461 a_11067_66191# a_10515_63143# 1.17fF
C8462 a_19282_13874# a_19374_13508# 0.32fF
C8463 a_31971_37737# VDD 0.59fF
C8464 vcm_commonmode a_39362_20902# 0.31fF
C8465 a_12809_8945# VDD 0.39fF
C8466 a_24302_68218# a_24394_68218# 0.32fF
C8467 a_31768_55394# a_12355_15055# 0.40fF
C8468 vcm_commonmode a_28318_63198# 0.31fF
C8469 a_2292_17179# a_5639_15279# 0.96fF
C8470 a_11067_46823# a_20635_29415# 6.21fF
C8471 a_19720_55394# a_12516_7093# 0.40fF
C8472 a_6559_59879# a_2419_48783# 0.58fF
C8473 a_23390_7484# a_24394_7484# 0.97fF
C8474 a_46482_8488# a_46482_7484# 1.00fF
C8475 vcm_commonmode a_22386_9492# 0.87fF
C8476 a_23736_7638# a_23390_17524# 0.38fF
C8477 a_36797_27497# a_37446_21540# 0.38fF
C8478 a_41967_31375# a_12877_16911# 0.41fF
C8479 a_33430_24552# m3_33332_24990# 1.39fF
C8480 a_27797_29423# VDD 0.53fF
C8481 vcm_commonmode a_38450_16520# 0.87fF
C8482 a_19374_64202# ctopp 3.59fF
C8483 ctopn a_24394_13508# 3.59fF
C8484 a_4351_67279# a_2872_44111# 0.35fF
C8485 a_28318_72234# VDD 0.62fF
C8486 vcm_commonmode a_22294_59182# 0.31fF
C8487 a_32426_12504# VDD 0.51fF
C8488 a_6559_42479# VDD 0.42fF
C8489 a_4758_45369# a_5039_42167# 0.79fF
C8490 a_22291_29415# a_36904_28879# 0.62fF
C8491 a_34434_9492# a_35438_9492# 0.97fF
C8492 vcm_commonmode a_39362_12870# 0.31fF
C8493 a_17366_64202# a_18370_64202# 0.97fF
C8494 a_35438_13508# a_35438_12504# 1.00fF
C8495 a_7841_29673# a_8383_27247# 0.41fF
C8496 a_4443_46607# a_1761_27791# 1.26fF
C8497 a_7155_55509# a_2840_66103# 1.34fF
C8498 a_3339_32463# VDD 10.84fF
C8499 a_27406_21540# VDD 0.51fF
C8500 vcm_commonmode a_30418_7484# 0.69fF
C8501 a_6467_55527# a_29361_51727# 2.32fF
C8502 a_35601_27497# a_12895_13967# 0.41fF
C8503 a_7841_29673# VDD 0.75fF
C8504 a_45478_58178# VDD 0.51fF
C8505 a_11067_66191# a_12985_7663# 1.68fF
C8506 a_1761_40847# a_12663_39783# 0.54fF
C8507 a_13349_37973# a_16744_40517# 0.32fF
C8508 a_39389_52271# a_39454_59182# 0.38fF
C8509 vcm_commonmode a_34342_21906# 0.31fF
C8510 a_28410_69222# ctopp 3.59fF
C8511 a_47486_72234# m3_47388_72146# 2.80fF
C8512 a_40527_41271# VDD 0.60fF
C8513 vcm_commonmode a_24394_64202# 0.87fF
C8514 a_32426_17524# VDD 0.51fF
C8515 a_19374_60186# VDD 0.51fF
C8516 a_20359_29199# a_28757_27247# 1.44fF
C8517 a_21187_29415# a_33694_30761# 0.50fF
C8518 vcm_commonmode a_39362_17890# 0.31fF
C8519 a_26402_65206# ctopp 3.59fF
C8520 a_12641_43124# a_23567_42035# 0.44fF
C8521 a_25398_67214# a_25398_66210# 1.00fF
C8522 vcm_commonmode a_26310_60186# 0.31fF
C8523 a_21371_52263# a_26402_61190# 0.38fF
C8524 a_42709_29199# a_48490_10496# 0.38fF
C8525 a_43270_27791# a_45478_11500# 0.38fF
C8526 a_33864_28111# a_12877_16911# 0.41fF
C8527 a_6835_46823# a_7387_48469# 0.33fF
C8528 a_21382_65206# a_21382_64202# 1.00fF
C8529 a_38358_13874# a_38450_13508# 0.32fF
C8530 a_12725_44527# a_13067_38517# 1.03fF
C8531 a_16955_52047# a_6831_63303# 0.35fF
C8532 a_39222_48169# a_40458_64202# 0.38fF
C8533 a_43378_68218# a_43470_68218# 0.32fF
C8534 a_25971_52263# a_12257_56623# 0.40fF
C8535 a_2595_47653# a_1775_47381# 0.34fF
C8536 a_27509_47695# VDD 0.47fF
C8537 vcm_commonmode a_33430_69222# 0.87fF
C8538 a_18151_52263# a_5915_30287# 0.33fF
C8539 a_42466_7484# a_43470_7484# 0.97fF
C8540 a_24302_56170# a_24394_56170# 0.32fF
C8541 a_21371_50959# a_10515_22671# 0.40fF
C8542 vcm_commonmode a_40458_22544# 0.87fF
C8543 a_6435_10901# VDD 0.49fF
C8544 a_26402_69222# a_27406_69222# 0.97fF
C8545 vcm_commonmode a_31422_65206# 0.87fF
C8546 a_26748_7638# a_26402_8488# 0.38fF
C8547 ctopn a_40675_27791# 2.62fF
C8548 a_33430_18528# VDD 0.51fF
C8549 a_33041_51157# VDD 0.61fF
C8550 a_19720_55394# a_16955_52047# 0.31fF
C8551 a_21382_61190# a_21382_60186# 1.00fF
C8552 ctopn a_31422_8488# 3.40fF
C8553 a_2559_67477# VDD 0.42fF
C8554 a_36442_64202# a_37446_64202# 0.97fF
C8555 vcm_commonmode a_40366_18894# 0.31fF
C8556 a_33430_66210# ctopp 3.59fF
C8557 vcm_commonmode a_20286_24918# 0.31fF
C8558 a_43269_29967# a_47486_10496# 0.38fF
C8559 a_24394_55166# VDD 0.60fF
C8560 a_33430_22544# a_34434_22544# 0.97fF
C8561 a_42709_29199# a_12877_16911# 0.40fF
C8562 vcm_commonmode a_36442_14512# 0.87fF
C8563 a_18611_52047# a_23390_58178# 0.38fF
C8564 a_24394_65206# a_25398_65206# 0.97fF
C8565 vcm_commonmode a_31330_55166# 0.30fF
C8566 a_42466_10496# VDD 0.51fF
C8567 a_41872_29423# a_43470_65206# 0.38fF
C8568 a_20378_17524# a_20378_16520# 1.00fF
C8569 vcm_commonmode a_22294_57174# 0.31fF
C8570 a_4191_33449# a_5039_42167# 0.72fF
C8571 a_31422_72234# a_31422_71230# 1.00fF
C8572 a_2959_47113# a_4482_57863# 0.38fF
C8573 vcm_commonmode a_49402_10862# 0.30fF
C8574 a_12355_15055# a_2872_44111# 0.89fF
C8575 a_40675_27791# a_41462_21540# 0.38fF
C8576 a_17712_7638# a_17366_21540# 0.38fF
C8577 a_24394_56170# a_24394_55166# 1.00fF
C8578 a_5023_72068# VDD 0.61fF
C8579 a_44474_67214# a_44474_66210# 1.00fF
C8580 vcm_commonmode a_41462_23548# 0.87fF
C8581 a_14919_43421# VDD 1.63fF
C8582 a_5682_69367# a_7580_61751# 0.88fF
C8583 vcm_commonmode a_38450_66210# 0.87fF
C8584 a_41427_52263# a_12983_63151# 0.40fF
C8585 a_13669_37429# a_1761_30511# 0.43fF
C8586 a_33041_51157# a_33313_51157# 0.49fF
C8587 a_22921_52245# VDD 0.54fF
C8588 a_2775_46025# a_9963_50959# 1.49fF
C8589 a_9503_26151# a_12877_16911# 0.41fF
C8590 a_29414_62194# VDD 0.51fF
C8591 a_23298_61190# a_23390_61190# 0.32fF
C8592 a_32426_55166# m3_32328_55078# 2.09fF
C8593 a_10055_58791# a_32951_27247# 0.41fF
C8594 ctopn a_16362_9492# 1.35fF
C8595 a_19720_7638# a_19374_23548# 0.38fF
C8596 a_11067_67279# VDD 17.23fF
C8597 a_40458_65206# a_40458_64202# 1.00fF
C8598 ctopn a_32426_16520# 3.59fF
C8599 vcm_commonmode a_36350_62194# 0.31fF
C8600 a_41872_29423# a_12981_62313# 0.40fF
C8601 a_39389_52271# a_39454_57174# 0.38fF
C8602 a_22015_28111# a_24959_30503# 2.56fF
C8603 a_37446_15516# VDD 0.51fF
C8604 a_39299_48783# a_44474_70226# 0.38fF
C8605 a_9503_26151# a_20378_13508# 0.38fF
C8606 a_24394_19532# a_25398_19532# 0.97fF
C8607 a_34434_23548# a_34434_22544# 1.00fF
C8608 vcm_commonmode a_44382_15882# 0.31fF
C8609 a_37446_63198# ctopp 3.64fF
C8610 a_43378_56170# a_43470_56170# 0.32fF
C8611 a_35438_71230# VDD 0.58fF
C8612 a_28410_66210# a_28410_65206# 1.00fF
C8613 a_29414_14512# a_30418_14512# 0.97fF
C8614 a_40403_37683# VDD 2.01fF
C8615 a_1823_66941# a_5252_56891# 0.60fF
C8616 a_47486_11500# VDD 0.51fF
C8617 a_42375_42089# VDD 0.67fF
C8618 a_43267_31055# a_46482_66210# 0.38fF
C8619 a_45478_69222# a_46482_69222# 0.97fF
C8620 a_12381_35836# a_12549_35836# 2.73fF
C8621 a_28959_49783# VDD 0.89fF
C8622 vcm_commonmode a_42374_71230# 0.31fF
C8623 a_40458_61190# a_40458_60186# 1.00fF
C8624 a_26310_8854# a_26402_8488# 0.32fF
C8625 a_31422_59182# ctopp 3.59fF
C8626 a_40050_48463# a_45478_62194# 0.38fF
C8627 a_27314_70226# a_27406_70226# 0.32fF
C8628 a_40050_48463# a_12727_67753# 0.40fF
C8629 a_26402_62194# a_26402_61190# 1.00fF
C8630 a_17366_10496# a_17366_9492# 1.00fF
C8631 vcm_commonmode a_21290_13874# 0.31fF
C8632 a_10055_58791# a_43175_28335# 0.41fF
C8633 a_7755_68591# VDD 0.72fF
C8634 a_43470_65206# a_44474_65206# 0.97fF
C8635 vcm_commonmode a_42466_63198# 0.92fF
C8636 a_39454_17524# a_39454_16520# 1.00fF
C8637 a_42985_46831# m2_48260_54946# 0.61fF
C8638 a_12907_27023# VDD 18.14fF
C8639 a_12901_66665# a_16362_71230# 19.89fF
C8640 a_2099_59861# a_4443_46607# 0.90fF
C8641 a_26402_20536# a_26402_19532# 1.00fF
C8642 a_3247_20495# a_4427_25071# 0.34fF
C8643 a_1757_21807# VDD 0.61fF
C8644 a_34434_23548# a_35438_23548# 0.97fF
C8645 a_39389_52271# VDD 6.63fF
C8646 vcm_commonmode a_36442_59182# 0.87fF
C8647 a_31422_66210# a_32426_66210# 0.97fF
C8648 vcm_commonmode a_11067_21583# 6.32fF
C8649 vcm_commonmode m3_16264_60098# 3.21fF
C8650 a_25971_52263# a_10975_66407# 0.40fF
C8651 a_25419_50959# a_22015_28111# 0.80fF
C8652 a_5271_17999# VDD 0.60fF
C8653 a_5023_72068# a_4885_71855# 0.70fF
C8654 vcm_commonmode a_39299_48783# 10.07fF
C8655 a_4482_57863# a_8295_47388# 0.39fF
C8656 a_1761_27791# a_13097_36367# 0.80fF
C8657 a_42374_61190# a_42466_61190# 0.32fF
C8658 a_5653_60039# a_5749_60039# 0.34fF
C8659 a_35438_60186# ctopp 3.59fF
C8660 a_6095_44807# a_9240_53877# 0.62fF
C8661 a_38450_68218# VDD 0.51fF
C8662 a_21049_34717# VDD 0.87fF
C8663 vcm_commonmode a_16746_18526# 5.36fF
C8664 a_38358_7850# VDD 0.62fF
C8665 ctopn a_34434_22544# 3.58fF
C8666 a_7917_13885# VDD 0.68fF
C8667 a_40691_47375# VDD 0.35fF
C8668 a_43362_28879# a_12901_66959# 0.40fF
C8669 a_31422_71230# a_31422_70226# 1.00fF
C8670 vcm_commonmode a_45386_68218# 0.31fF
C8671 a_43470_19532# a_44474_19532# 0.97fF
C8672 a_22921_52245# a_23193_52245# 0.50fF
C8673 a_6467_55527# a_21267_52047# 0.38fF
C8674 a_28547_51175# a_29927_29199# 1.58fF
C8675 VDD rst_n 1.77fF
C8676 a_3143_66972# VDD 3.36fF
C8677 a_47486_66210# a_47486_65206# 1.00fF
C8678 a_48490_14512# a_49494_14512# 0.97fF
C8679 vcm_commonmode a_48490_21540# 0.87fF
C8680 a_11067_67279# a_11619_56615# 0.73fF
C8681 a_17039_51157# a_4443_46607# 0.46fF
C8682 a_22843_29415# a_22015_28111# 0.37fF
C8683 a_7815_49855# VDD 0.57fF
C8684 a_21371_50959# a_12901_66665# 0.40fF
C8685 a_47486_72234# a_48490_72234# 0.97fF
C8686 a_27406_20536# a_28410_20536# 0.97fF
C8687 a_45386_8854# a_45478_8488# 0.32fF
C8688 vcm_commonmode a_25398_10496# 0.87fF
C8689 a_1823_65853# VDD 1.61fF
C8690 a_2787_32679# a_2216_28309# 0.54fF
C8691 a_22015_28111# a_23395_32463# 1.07fF
C8692 ctopn a_30418_14512# 3.59fF
C8693 a_2401_41941# a_1761_41935# 0.58fF
C8694 vcm_commonmode a_40458_60186# 0.87fF
C8695 a_14646_29423# a_14926_31849# 1.07fF
C8696 a_46390_70226# a_46482_70226# 0.32fF
C8697 a_3231_53047# VDD 0.39fF
C8698 a_12641_37684# a_13097_37455# 0.80fF
C8699 a_6835_46823# a_25015_48437# 1.04fF
C8700 a_45478_62194# a_45478_61190# 1.00fF
C8701 a_36442_10496# a_36442_9492# 1.00fF
C8702 a_38450_56170# VDD 0.52fF
C8703 a_10055_58791# a_43270_27791# 0.41fF
C8704 a_14963_39783# a_19203_39958# 0.32fF
C8705 a_32795_36415# VDD 0.96fF
C8706 a_21382_8488# VDD 0.58fF
C8707 a_12907_56399# a_12355_15055# 0.77fF
C8708 a_27314_16886# a_27406_16520# 0.32fF
C8709 vcm_commonmode a_45386_56170# 0.31fF
C8710 ctopn a_35438_23548# 3.40fF
C8711 a_5451_14735# VDD 0.35fF
C8712 a_5179_47919# VDD 0.42fF
C8713 a_45478_20536# a_45478_19532# 1.00fF
C8714 a_8592_58255# VDD 0.45fF
C8715 vcm_commonmode a_28318_8854# 0.31fF
C8716 a_13349_37973# a_13837_38772# 1.18fF
C8717 vcm_commonmode a_20378_15516# 0.87fF
C8718 a_38557_32143# a_20635_29415# 6.58fF
C8719 a_31422_57174# ctopp 3.58fF
C8720 a_17507_52047# a_12901_58799# 0.40fF
C8721 a_75475_38962# VDD 1.05fF
C8722 ctopn a_44474_19532# 3.59fF
C8723 a_4811_34855# a_17869_28585# 0.69fF
C8724 a_20267_30503# a_12447_29199# 0.52fF
C8725 a_28959_49783# a_29055_49525# 0.76fF
C8726 a_17039_51157# a_20195_49793# 0.71fF
C8727 a_3983_50095# VDD 0.56fF
C8728 vcm_commonmode a_18370_71230# 0.87fF
C8729 a_25398_21540# a_25398_20536# 1.00fF
C8730 a_37446_61190# VDD 0.51fF
C8731 vcm_commonmode a_30418_11500# 0.87fF
C8732 a_3668_56311# VDD 6.78fF
C8733 a_27406_12504# a_28410_12504# 0.97fF
C8734 a_5449_25071# a_5211_24759# 0.50fF
C8735 a_33338_67214# a_33430_67214# 0.32fF
C8736 vcm_commonmode a_44382_61190# 0.31fF
C8737 vcm_commonmode a_34434_24552# 0.84fF
C8738 a_24959_30503# a_22291_29415# 2.42fF
C8739 vcm_commonmode a_16746_67216# 5.36fF
C8740 a_1770_14441# a_2021_17973# 1.37fF
C8741 a_7097_63151# VDD 0.32fF
C8742 a_11067_46823# a_12899_2767# 0.46fF
C8743 a_45478_62194# ctopp 3.59fF
C8744 a_27752_7638# a_27406_23548# 0.38fF
C8745 a_41462_70226# VDD 0.51fF
C8746 a_1770_14441# a_2605_60975# 0.61fF
C8747 a_10317_13647# a_10351_12879# 0.40fF
C8748 a_12985_16367# a_16746_10494# 0.41fF
C8749 a_19283_37737# VDD 0.61fF
C8750 a_12727_67753# ctopp 3.23fF
C8751 vcm_commonmode a_44474_55166# 0.84fF
C8752 a_18151_52263# a_12355_15055# 0.43fF
C8753 a_9503_26151# a_20378_7484# 0.34fF
C8754 vcm_commonmode a_36442_57174# 0.87fF
C8755 a_14831_50095# a_28108_48463# 1.37fF
C8756 a_22386_16520# VDD 0.51fF
C8757 vcm_commonmode a_48398_70226# 0.31fF
C8758 a_46482_20536# a_47486_20536# 0.97fF
C8759 a_10649_58947# VDD 0.40fF
C8760 a_19282_7850# a_19374_7484# 0.32fF
C8761 a_26402_24552# m3_26304_24414# 2.81fF
C8762 a_35438_63198# a_36442_63198# 0.97fF
C8763 vcm_commonmode a_29322_16886# 0.31fF
C8764 a_21290_72234# VDD 0.62fF
C8765 ctopn a_47486_20536# 3.58fF
C8766 a_1761_47919# a_1761_46287# 2.79fF
C8767 a_31611_43447# VDD 0.63fF
C8768 a_35346_58178# a_35438_58178# 0.32fF
C8769 a_1768_13103# a_1761_22895# 7.89fF
C8770 a_6831_63303# a_26417_47919# 1.11fF
C8771 a_22386_21540# a_23390_21540# 0.97fF
C8772 a_30326_9858# a_30418_9492# 0.32fF
C8773 a_11067_66191# a_2872_44111# 0.63fF
C8774 a_46390_16886# a_46482_16520# 0.32fF
C8775 a_1761_50639# a_1761_46287# 0.42fF
C8776 a_12907_27023# a_34482_29941# 6.59fF
C8777 vcm_commonmode a_21382_68218# 0.87fF
C8778 a_2143_15271# a_2411_18517# 1.06fF
C8779 a_30418_58178# VDD 0.51fF
C8780 a_29414_59182# a_30418_59182# 0.97fF
C8781 ctopn a_47486_12504# 3.58fF
C8782 a_16746_56172# ctopp 1.42fF
C8783 a_34251_52263# a_35438_59182# 0.38fF
C8784 a_11067_67279# a_24740_7638# 0.41fF
C8785 a_27406_17524# a_28410_17524# 0.97fF
C8786 a_5915_30287# a_3339_30503# 1.27fF
C8787 a_9135_27239# a_12877_14441# 0.41fF
C8788 a_44474_21540# a_44474_20536# 1.00fF
C8789 a_3141_59887# VDD 0.88fF
C8790 a_31422_24552# a_31422_23548# 1.00fF
C8791 a_35601_27497# a_35438_22544# 0.38fF
C8792 a_47486_67214# VDD 0.51fF
C8793 ctopp m3_33332_55078# 0.31fF
C8794 a_46482_12504# a_47486_12504# 0.97fF
C8795 a_1761_46287# a_14963_39783# 0.98fF
C8796 vcm_commonmode a_16362_60186# 4.47fF
C8797 a_17599_52263# a_22386_61190# 0.38fF
C8798 ctopn a_42466_21540# 3.59fF
C8799 a_1761_52815# a_12341_41281# 0.45fF
C8800 a_11067_47695# a_5039_42167# 0.30fF
C8801 a_1586_18695# VDD 11.41fF
C8802 a_9240_53877# VDD 1.00fF
C8803 a_11251_59879# a_8295_47388# 1.20fF
C8804 a_18979_30287# a_43680_29941# 0.46fF
C8805 a_2959_47113# a_2775_46025# 1.64fF
C8806 vcm_commonmode a_35438_13508# 0.87fF
C8807 ctopn a_19374_10496# 3.59fF
C8808 a_17366_69222# VDD 0.58fF
C8809 a_7295_44647# a_7841_12167# 0.57fF
C8810 a_33080_37149# VDD 1.57fF
C8811 ctopn a_47486_17524# 3.58fF
C8812 a_8583_33551# a_7862_34025# 0.40fF
C8813 a_2021_22325# a_12381_43957# 4.24fF
C8814 a_33856_44869# a_24800_43041# 0.41fF
C8815 a_44474_9492# VDD 0.51fF
C8816 a_36717_47375# a_36442_64202# 0.38fF
C8817 a_18611_52047# a_12257_56623# 0.40fF
C8818 vcm_commonmode a_21382_56170# 0.87fF
C8819 a_22843_29415# a_22291_29415# 7.17fF
C8820 a_18413_47919# VDD 0.99fF
C8821 vcm_commonmode a_24302_69222# 0.31fF
C8822 a_2419_48783# a_6646_50639# 0.69fF
C8823 a_38358_7850# a_38450_7484# 0.32fF
C8824 a_24394_22544# VDD 0.51fF
C8825 a_5085_23047# a_6773_27805# 0.83fF
C8826 a_12357_37999# a_1799_29556# 3.16fF
C8827 a_14287_51175# a_10515_22671# 0.42fF
C8828 vcm_commonmode a_31330_22910# 0.31fF
C8829 a_19374_70226# ctopp 3.58fF
C8830 a_2473_34293# a_2899_28111# 0.35fF
C8831 a_4811_34855# a_12899_3855# 0.87fF
C8832 a_22294_69222# a_22386_69222# 0.32fF
C8833 vcm_commonmode a_22294_65206# 0.31fF
C8834 a_28410_18528# a_28410_17524# 1.00fF
C8835 a_10883_71855# a_11049_71855# 0.72fF
C8836 a_41462_21540# a_42466_21540# 0.97fF
C8837 a_49402_9858# a_49494_9492# 0.32fF
C8838 a_10055_58791# a_12341_3311# 0.46fF
C8839 a_41967_31375# a_12895_13967# 0.41fF
C8840 a_4563_32900# a_4123_37013# 0.81fF
C8841 a_32334_64202# a_32426_64202# 0.32fF
C8842 a_1770_14441# a_2411_19605# 0.87fF
C8843 a_12725_44527# a_12473_41781# 0.35fF
C8844 vcm_commonmode a_20378_61190# 0.87fF
C8845 a_20378_14512# VDD 0.51fF
C8846 a_48490_59182# a_49494_59182# 0.97fF
C8847 a_29322_22910# a_29414_22544# 0.32fF
C8848 a_46482_64202# VDD 0.51fF
C8849 a_18370_10496# a_19374_10496# 0.97fF
C8850 vcm_commonmode a_27314_14878# 0.31fF
C8851 ctopn a_24394_11500# 3.59fF
C8852 a_19629_39631# a_20713_40193# 0.62fF
C8853 a_19720_55394# a_19374_58178# 0.38fF
C8854 a_20286_65206# a_20378_65206# 0.32fF
C8855 a_29414_14512# a_29414_13508# 1.00fF
C8856 a_27652_38237# VDD 2.10fF
C8857 ctopn a_48490_18528# 3.43fF
C8858 VDD result_out[10] 1.18fF
C8859 a_12677_40157# VDD 1.11fF
C8860 a_39389_52271# a_39454_65206# 0.38fF
C8861 a_12877_16911# a_12727_13353# 1.02fF
C8862 a_46482_17524# a_47486_17524# 0.97fF
C8863 a_10055_58791# a_12985_16367# 23.90fF
C8864 a_23774_49551# VDD 1.08fF
C8865 a_27406_72234# a_27406_71230# 1.00fF
C8866 vcm_commonmode a_24394_70226# 0.87fF
C8867 a_41462_58178# vcm_commonmode 0.87fF
C8868 a_33430_60186# a_34434_60186# 0.97fF
C8869 a_25398_23548# VDD 0.52fF
C8870 a_36629_27791# a_36442_21540# 0.38fF
C8871 a_12341_3311# a_22386_22544# 0.38fF
C8872 a_22386_66210# VDD 0.51fF
C8873 a_35438_12504# a_35438_11500# 1.00fF
C8874 a_6162_28487# a_6773_27805# 0.30fF
C8875 vcm_commonmode a_32334_23914# 0.31fF
C8876 a_4443_46607# a_2787_32679# 1.30fF
C8877 a_10351_12879# VDD 0.40fF
C8878 a_12249_43457# VDD 1.76fF
C8879 a_22386_70226# a_22386_69222# 1.00fF
C8880 vcm_commonmode a_29322_66210# 0.31fF
C8881 a_34780_56398# a_12983_63151# 0.40fF
C8882 a_28410_18528# a_29414_18528# 0.97fF
C8883 a_34434_19532# VDD 0.51fF
C8884 vcm_commonmode a_13183_52047# 10.36fF
C8885 a_28756_7638# a_12727_13353# 0.41fF
C8886 a_11067_23759# a_12899_10927# 0.37fF
C8887 vcm_commonmode a_41370_19898# 0.31fF
C8888 a_25398_67214# ctopp 3.59fF
C8889 a_36717_47375# a_12981_62313# 0.40fF
C8890 vcm_commonmode a_9135_27239# 10.35fF
C8891 a_34251_52263# a_35438_57174# 0.38fF
C8892 a_7289_70767# a_2689_65103# 0.38fF
C8893 a_39222_48169# a_40458_70226# 0.38fF
C8894 a_20286_19898# a_20378_19532# 0.32fF
C8895 a_4891_47388# VDD 10.28fF
C8896 vcm_commonmode a_42466_8488# 0.86fF
C8897 a_33864_28111# a_12895_13967# 0.41fF
C8898 a_21382_11500# a_21382_10496# 1.00fF
C8899 a_11619_56615# a_1586_18695# 0.75fF
C8900 a_7461_27247# a_3301_26703# 0.30fF
C8901 a_25306_14878# a_25398_14512# 0.32fF
C8902 a_28011_41855# VDD 1.05fF
C8903 a_41370_69222# a_41462_69222# 0.32fF
C8904 a_41261_28335# a_42466_66210# 0.38fF
C8905 a_47486_18528# a_47486_17524# 1.00fF
C8906 a_2004_42453# a_2007_20149# 0.84fF
C8907 ctopn a_25744_7638# 2.62fF
C8908 a_5915_35943# a_3339_30503# 0.44fF
C8909 a_2295_17429# VDD 0.43fF
C8910 a_25971_52263# a_30418_72234# 0.34fF
C8911 a_42718_27497# a_44474_16520# 0.38fF
C8912 a_19374_55166# a_20378_55166# 0.97fF
C8913 a_42374_24918# VDD 0.36fF
C8914 a_2840_53511# a_3228_54171# 0.76fF
C8915 a_4903_31849# VDD 2.51fF
C8916 a_41427_52263# a_41462_62194# 0.38fF
C8917 a_23395_32463# a_27417_32509# 0.73fF
C8918 a_5179_47919# a_5345_47919# 0.66fF
C8919 a_1778_42631# VDD 0.76fF
C8920 vcm_commonmode a_30418_67214# 0.87fF
C8921 a_38557_32143# a_12727_67753# 0.40fF
C8922 a_37446_20536# VDD 0.51fF
C8923 a_48398_22910# a_48490_22544# 0.32fF
C8924 a_26402_63198# VDD 0.57fF
C8925 a_37446_10496# a_38450_10496# 0.97fF
C8926 a_23736_7638# a_23390_21540# 0.38fF
C8927 a_28756_7638# a_10515_23975# 0.41fF
C8928 a_39362_65206# a_39454_65206# 0.32fF
C8929 a_48490_14512# a_48490_13508# 1.00fF
C8930 vcm_commonmode a_44382_20902# 0.31fF
C8931 a_25300_39655# VDD 1.43fF
C8932 vcm_commonmode a_33338_63198# 0.31fF
C8933 a_28524_47919# VDD 0.80fF
C8934 a_20378_59182# VDD 0.51fF
C8935 vcm_commonmode a_27406_9492# 0.87fF
C8936 a_10515_23975# a_16362_22544# 19.89fF
C8937 a_30326_23914# a_30418_23548# 0.32fF
C8938 a_42709_29199# a_12895_13967# 0.40fF
C8939 a_13643_28327# a_14926_31849# 0.68fF
C8940 a_6831_63303# a_6467_55527# 0.83fF
C8941 a_23390_11500# a_24394_11500# 0.97fF
C8942 vcm_commonmode a_43470_16520# 0.87fF
C8943 a_24394_64202# ctopp 3.59fF
C8944 ctopn a_29414_13508# 3.59fF
C8945 a_2411_26133# a_2339_38129# 0.66fF
C8946 a_28547_51175# VDD 9.70fF
C8947 a_27314_66210# a_27406_66210# 0.32fF
C8948 vcm_commonmode a_27314_59182# 0.31fF
C8949 a_2292_17179# a_5179_10927# 0.52fF
C8950 vcm_commonmode a_12546_22351# 6.31fF
C8951 a_15548_30761# a_14361_29967# 0.36fF
C8952 a_2787_30503# a_6459_30511# 0.38fF
C8953 a_37446_12504# VDD 0.51fF
C8954 a_41462_70226# a_41462_69222# 1.00fF
C8955 a_18611_52047# a_10975_66407# 0.45fF
C8956 a_43270_27791# a_45478_10496# 0.38fF
C8957 a_47486_18528# a_48490_18528# 0.97fF
C8958 a_12899_10927# a_16746_17522# 0.41fF
C8959 vcm_commonmode a_36613_48169# 10.02fF
C8960 vcm_commonmode a_44382_12870# 0.31fF
C8961 a_27406_24552# a_28410_24552# 0.97fF
C8962 a_3339_32463# a_5363_30503# 1.33fF
C8963 a_23929_47381# VDD 0.57fF
C8964 a_39222_48169# a_12901_66959# 0.40fF
C8965 a_39362_19898# a_39454_19532# 0.32fF
C8966 a_32426_21540# VDD 0.51fF
C8967 vcm_commonmode a_35438_7484# 0.69fF
C8968 a_9503_26151# a_12895_13967# 0.41fF
C8969 a_24394_62194# a_25398_62194# 0.97fF
C8970 a_40458_11500# a_40458_10496# 1.00fF
C8971 a_1952_60431# a_2913_54991# 0.41fF
C8972 a_3452_70537# VDD 0.33fF
C8973 a_44382_14878# a_44474_14512# 0.32fF
C8974 vcm_commonmode a_39362_21906# 0.31fF
C8975 a_33430_69222# ctopp 3.59fF
C8976 a_14926_31849# a_23195_29967# 0.31fF
C8977 a_6372_38279# VDD 4.34fF
C8978 vcm_commonmode a_29414_64202# 0.87fF
C8979 a_1761_35407# a_33963_35507# 0.34fF
C8980 a_37446_17524# VDD 0.51fF
C8981 a_39299_48783# a_40050_48463# 2.20fF
C8982 a_41872_29423# a_43267_31055# 0.66fF
C8983 a_14287_51175# a_12901_66665# 0.40fF
C8984 a_4891_47388# a_23193_52245# 0.74fF
C8985 a_32951_27247# a_12877_14441# 0.41fF
C8986 a_23298_20902# a_23390_20536# 0.32fF
C8987 a_24394_60186# VDD 0.51fF
C8988 a_37446_55166# a_38450_55166# 0.97fF
C8989 a_1757_66415# VDD 0.62fF
C8990 vcm_commonmode a_44382_17890# 0.31fF
C8991 a_31422_65206# ctopp 3.59fF
C8992 a_14287_51175# a_6646_50639# 0.38fF
C8993 a_12899_3855# a_11902_27497# 0.40fF
C8994 a_29414_57174# a_30418_57174# 0.97fF
C8995 vcm_commonmode a_31330_60186# 0.31fF
C8996 a_32426_15516# a_33430_15516# 0.97fF
C8997 a_9503_26151# a_20378_11500# 0.38fF
C8998 a_5541_53609# VDD 0.40fF
C8999 a_30764_7638# a_30418_24552# 0.46fF
C9000 vcm_commonmode a_17366_19532# 1.82fF
C9001 a_11710_58487# a_11659_66567# 0.63fF
C9002 a_30418_71230# a_31422_71230# 0.97fF
C9003 vcm_commonmode a_38450_69222# 0.87fF
C9004 a_10515_22671# a_12901_58799# 23.69fF
C9005 a_49402_23914# a_49494_23548# 0.32fF
C9006 a_27752_7638# a_12899_10927# 0.41fF
C9007 a_29927_29199# a_34267_31599# 0.40fF
C9008 a_42466_11500# a_43470_11500# 0.97fF
C9009 a_46390_66210# a_46482_66210# 0.32fF
C9010 vcm_commonmode a_45478_22544# 0.87fF
C9011 vcm_commonmode m3_16264_21402# 3.21fF
C9012 a_27747_42359# VDD 0.63fF
C9013 vcm_commonmode a_36442_65206# 0.87fF
C9014 a_5682_69367# a_5254_67503# 1.78fF
C9015 a_39299_48783# a_12355_65103# 0.40fF
C9016 a_37919_28111# a_38450_9492# 0.38fF
C9017 a_12713_36483# a_21856_36513# 0.34fF
C9018 a_38450_18528# VDD 0.51fF
C9019 a_21290_72234# a_21382_72234# 0.32fF
C9020 a_43175_28335# a_12877_14441# 0.41fF
C9021 a_42709_29199# a_48490_15516# 0.38fF
C9022 a_18370_24552# VDD 0.61fF
C9023 vcm_commonmode a_21290_11866# 0.31fF
C9024 ctopn a_36442_8488# 3.40fF
C9025 a_46482_24552# a_47486_24552# 0.97fF
C9026 a_24740_7638# a_24394_22544# 0.38fF
C9027 a_9135_67503# VDD 0.41fF
C9028 a_2840_66103# a_6559_59879# 0.82fF
C9029 a_23298_12870# a_23390_12504# 0.32fF
C9030 vcm_commonmode a_45386_18894# 0.31fF
C9031 a_38450_66210# ctopp 3.59fF
C9032 vcm_commonmode a_25306_24918# 0.31fF
C9033 a_4443_46607# a_6559_22671# 1.70fF
C9034 a_19807_28111# a_18979_30287# 1.79fF
C9035 a_43267_31055# a_46482_69222# 0.38fF
C9036 a_18370_59182# a_18370_58178# 1.00fF
C9037 a_29414_55166# VDD 0.60fF
C9038 a_8583_33551# a_38115_52263# 0.61fF
C9039 a_43470_62194# a_44474_62194# 0.97fF
C9040 a_23447_28853# VDD 0.39fF
C9041 a_20378_57174# VDD 0.51fF
C9042 vcm_commonmode a_41462_14512# 0.87fF
C9043 a_5455_37039# VDD 0.41fF
C9044 vcm_commonmode a_20378_20536# 0.87fF
C9045 vcm_commonmode a_35346_55166# 0.30fF
C9046 a_47486_10496# VDD 0.51fF
C9047 a_29545_40193# VDD 1.32fF
C9048 vcm_commonmode a_27314_57174# 0.31fF
C9049 a_1761_35407# a_31959_34751# 0.42fF
C9050 a_31768_7638# a_31422_13508# 0.38fF
C9051 a_19720_7638# a_19374_14512# 0.38fF
C9052 a_42374_20902# a_42466_20536# 0.32fF
C9053 a_1643_59317# VDD 0.35fF
C9054 a_2411_26133# a_1591_38677# 0.34fF
C9055 a_19374_24552# m3_19276_24414# 2.81fF
C9056 a_31330_63198# a_31422_63198# 0.32fF
C9057 a_17507_52047# a_14831_50095# 1.14fF
C9058 a_22386_57174# a_22386_56170# 1.00fF
C9059 a_48490_57174# a_49494_57174# 0.97fF
C9060 vcm_commonmode a_46482_23548# 0.87fF
C9061 vcm_commonmode a_43470_66210# 0.87fF
C9062 a_18278_21906# a_18370_21540# 0.32fF
C9063 a_43269_29967# a_47486_15516# 0.38fF
C9064 a_34434_62194# VDD 0.51fF
C9065 vcm_commonmode a_20378_12504# 0.87fF
C9066 ctopn a_21382_9492# 3.58fF
C9067 a_13669_35253# VDD 5.20fF
C9068 ctopn a_37446_16520# 3.59fF
C9069 vcm_commonmode a_41370_62194# 0.31fF
C9070 vcm_commonmode a_32951_27247# 10.32fF
C9071 a_22015_28111# a_38067_47349# 0.61fF
C9072 a_42466_15516# VDD 0.51fF
C9073 a_25306_59182# a_25398_59182# 0.32fF
C9074 a_4149_20719# VDD 0.61fF
C9075 vcm_commonmode a_49402_15882# 0.30fF
C9076 a_42466_63198# ctopp 3.64fF
C9077 a_40458_71230# VDD 0.58fF
C9078 a_7000_65595# a_7039_65469# 0.46fF
C9079 a_31768_55394# a_31422_59182# 0.38fF
C9080 a_1689_10396# a_1929_12131# 0.63fF
C9081 a_4259_40847# VDD 0.62fF
C9082 a_12901_66959# a_16746_68220# 2.28fF
C9083 a_23298_17890# a_23390_17524# 0.32fF
C9084 a_40491_27247# a_43470_9492# 0.38fF
C9085 vcm_commonmode a_47394_71230# 0.31fF
C9086 a_43270_27791# a_12877_14441# 0.41fF
C9087 a_1761_27791# a_2235_30503# 1.22fF
C9088 a_36442_59182# ctopp 3.59fF
C9089 a_11067_47695# a_9731_22895# 0.35fF
C9090 a_29414_64202# a_29414_63198# 1.23fF
C9091 a_42374_12870# a_42466_12504# 0.32fF
C9092 a_22399_32143# VDD 0.57fF
C9093 vcm_commonmode a_20378_17524# 0.87fF
C9094 a_21663_42943# a_20897_42917# 0.32fF
C9095 a_14287_51175# a_18370_61190# 0.38fF
C9096 a_39299_48783# ctopp 2.63fF
C9097 a_15607_46805# a_4674_40277# 0.70fF
C9098 a_19374_13508# VDD 0.51fF
C9099 a_1761_44111# VDD 7.47fF
C9100 a_2021_17973# a_2411_19605# 0.83fF
C9101 a_8082_54599# VDD 0.35fF
C9102 a_21382_22544# a_21382_21540# 1.00fF
C9103 a_8491_27023# a_12899_10927# 0.41fF
C9104 a_30975_28023# VDD 0.33fF
C9105 vcm_commonmode a_26310_13874# 0.31fF
C9106 a_9135_27239# a_21382_24552# 0.46fF
C9107 a_28410_13508# a_29414_13508# 0.97fF
C9108 a_13835_36649# VDD 1.29fF
C9109 a_1761_22895# a_2021_17973# 0.33fF
C9110 vcm_commonmode a_47486_63198# 0.92fF
C9111 a_28547_51175# a_32426_64202# 0.38fF
C9112 a_5682_69367# a_8999_61493# 1.38fF
C9113 a_33430_68218# a_34434_68218# 0.97fF
C9114 vcm_commonmode a_43175_28335# 10.43fF
C9115 a_8583_33551# a_20267_30503# 0.44fF
C9116 a_1768_13103# a_1586_40455# 0.64fF
C9117 a_45478_56170# a_45478_55166# 1.00fF
C9118 a_41462_57174# a_41462_56170# 1.00fF
C9119 vcm_commonmode a_41462_59182# 0.87fF
C9120 a_3339_30503# a_15799_29941# 0.63fF
C9121 a_38499_42943# VDD 0.85fF
C9122 a_7841_12167# a_9765_32143# 0.40fF
C9123 a_37354_21906# a_37446_21540# 0.32fF
C9124 a_40458_60186# ctopp 3.59fF
C9125 a_18370_58178# a_18370_57174# 1.00fF
C9126 a_29760_7638# a_29414_23548# 0.38fF
C9127 a_43470_68218# VDD 0.51fF
C9128 a_1768_13103# a_3016_60949# 0.58fF
C9129 a_1954_61677# a_3295_54421# 0.39fF
C9130 vcm_commonmode a_21382_18528# 0.87fF
C9131 a_2099_59861# a_5346_33775# 1.85fF
C9132 a_43378_7850# VDD 0.62fF
C9133 a_25398_16520# a_25398_15516# 1.00fF
C9134 ctopn a_39454_22544# 3.58fF
C9135 a_12907_27023# a_24959_30503# 1.21fF
C9136 a_21187_29415# a_8491_41383# 2.56fF
C9137 a_2952_66139# a_2689_65103# 2.29fF
C9138 a_3339_43023# a_12357_37999# 2.34fF
C9139 a_10515_22671# a_16362_58178# 19.89fF
C9140 a_44382_59182# a_44474_59182# 0.32fF
C9141 a_32772_7638# a_32426_18528# 0.38fF
C9142 a_9599_57141# VDD 0.38fF
C9143 a_6008_69679# VDD 0.53fF
C9144 a_34251_52263# a_35438_65206# 0.38fF
C9145 a_42374_17890# a_42466_17524# 0.32fF
C9146 a_23390_72234# a_23390_71230# 1.00fF
C9147 a_29322_60186# a_29414_60186# 0.32fF
C9148 vcm_commonmode a_30418_10496# 0.87fF
C9149 a_9624_65301# VDD 1.03fF
C9150 a_48490_64202# a_48490_63198# 1.23fF
C9151 ctopn a_35438_14512# 3.59fF
C9152 a_1761_41935# a_3949_41935# 0.52fF
C9153 a_8123_56399# a_7265_56053# 1.18fF
C9154 a_42985_46831# a_12981_59343# 0.40fF
C9155 vcm_commonmode a_45478_60186# 0.87fF
C9156 a_18370_71230# ctopp 3.39fF
C9157 a_7841_12167# a_9955_20969# 1.08fF
C9158 a_29927_29199# a_18979_30287# 0.92fF
C9159 a_23901_44220# VDD 0.92fF
C9160 a_23395_52047# a_12983_63151# 0.40fF
C9161 a_24302_18894# a_24394_18528# 0.32fF
C9162 a_9135_27239# a_12899_11471# 0.41fF
C9163 a_40458_22544# a_40458_21540# 1.00fF
C9164 a_43470_56170# VDD 0.52fF
C9165 a_13669_39605# a_13837_39860# 0.44fF
C9166 a_47486_13508# a_48490_13508# 0.97fF
C9167 a_12621_36091# VDD 5.24fF
C9168 a_16746_67216# ctopp 1.68fF
C9169 a_26402_8488# VDD 0.58fF
C9170 a_29760_55394# a_12981_62313# 0.40fF
C9171 a_19374_68218# a_19374_67214# 1.00fF
C9172 vcm_commonmode a_17366_62194# 1.83fF
C9173 vcm_commonmode a_43270_27791# 10.47fF
C9174 a_31768_55394# a_31422_57174# 0.38fF
C9175 ctopn a_40458_23548# 3.40fF
C9176 a_7939_30503# a_3339_30503# 2.07fF
C9177 a_36717_47375# a_36442_70226# 0.38fF
C9178 vcm_commonmode a_33338_8854# 0.31fF
C9179 a_13349_37973# a_13909_38659# 0.46fF
C9180 a_1586_21959# VDD 10.50fF
C9181 vcm_commonmode a_25398_15516# 0.87fF
C9182 a_36442_57174# ctopp 3.58fF
C9183 a_33430_56170# a_34434_56170# 0.97fF
C9184 a_16362_71230# VDD 2.55fF
C9185 a_38557_32143# a_38450_66210# 0.38fF
C9186 a_1586_66567# a_5254_67503# 0.96fF
C9187 a_31768_7638# a_31422_7484# 0.34fF
C9188 a_1761_30511# a_13005_35823# 0.81fF
C9189 vcm_commonmode a_23390_71230# 0.86fF
C9190 a_36797_27497# a_37446_16520# 0.38fF
C9191 a_27752_7638# a_27406_14512# 0.38fF
C9192 a_42466_61190# VDD 0.51fF
C9193 a_1761_27791# a_1761_32143# 0.33fF
C9194 a_2959_47113# a_5190_59575# 1.07fF
C9195 vcm_commonmode a_35438_11500# 0.87fF
C9196 a_3339_32463# a_8423_39367# 1.05fF
C9197 a_26523_28111# ctopn 1.14fF
C9198 vcm_commonmode a_49402_61190# 0.30fF
C9199 a_36613_48169# a_37446_62194# 0.38fF
C9200 a_44474_16520# a_44474_15516# 1.00fF
C9201 vcm_commonmode a_39454_24552# 0.84fF
C9202 a_2292_43291# a_3983_45743# 0.31fF
C9203 a_29927_29199# a_37427_47893# 0.38fF
C9204 a_4842_45467# VDD 0.87fF
C9205 a_31768_55394# a_12727_67753# 0.40fF
C9206 vcm_commonmode a_21290_67214# 0.31fF
C9207 a_17366_70226# a_18370_70226# 0.97fF
C9208 a_29414_19532# a_29414_18528# 1.00fF
C9209 a_33338_10862# a_33430_10496# 0.32fF
C9210 a_46482_70226# VDD 0.51fF
C9211 a_25133_37571# VDD 3.24fF
C9212 a_21382_68218# ctopp 3.59fF
C9213 a_6459_30511# a_13390_29575# 0.45fF
C9214 a_8251_39367# VDD 0.34fF
C9215 vcm_commonmode a_41462_57174# 0.87fF
C9216 a_5915_30287# a_11143_31599# 0.38fF
C9217 a_22843_29415# a_12907_27023# 1.11fF
C9218 a_17682_50095# a_30005_48463# 0.36fF
C9219 a_27406_16520# VDD 0.51fF
C9220 a_21003_49007# VDD 0.45fF
C9221 a_12341_3311# a_12877_14441# 0.41fF
C9222 a_48398_60186# a_48490_60186# 0.32fF
C9223 vcm_commonmode a_18278_9858# 0.31fF
C9224 a_12907_27023# a_23395_32463# 0.32fF
C9225 a_19282_11866# a_19374_11500# 0.32fF
C9226 a_13353_30511# VDD 3.62fF
C9227 vcm_commonmode a_34342_16886# 0.31fF
C9228 a_1803_19087# a_12663_39783# 3.17fF
C9229 a_13576_42589# a_19967_41781# 0.86fF
C9230 a_21371_50959# VDD 11.52fF
C9231 a_24394_15516# a_24394_14512# 1.00fF
C9232 a_49494_7484# m3_49396_7346# 2.80fF
C9233 a_14926_31849# a_19626_31751# 0.54fF
C9234 a_26523_28111# a_8491_41383# 5.74fF
C9235 a_42188_43677# VDD 2.13fF
C9236 a_13183_52047# a_12355_65103# 0.41fF
C9237 a_43378_18894# a_43470_18528# 0.32fF
C9238 a_2847_18517# VDD 0.45fF
C9239 vcm_commonmode a_25971_52263# 10.02fF
C9240 a_32426_61190# a_33430_61190# 0.97fF
C9241 a_46482_55166# m3_46384_55078# 2.81fF
C9242 a_16362_60186# ctopp 1.35fF
C9243 a_23298_24918# a_23390_24552# 0.32fF
C9244 a_23567_35507# VDD 3.09fF
C9245 a_19374_7484# VDD 1.23fF
C9246 a_38450_68218# a_38450_67214# 1.00fF
C9247 a_4119_70741# a_6467_55527# 0.41fF
C9248 a_10515_63143# a_7841_12167# 0.50fF
C9249 a_11067_46823# a_7571_29199# 1.94fF
C9250 vcm_commonmode a_26402_68218# 0.87fF
C9251 a_25787_28327# a_12901_66959# 0.40fF
C9252 a_35438_58178# VDD 0.51fF
C9253 a_11053_62607# VDD 0.88fF
C9254 a_10680_52245# a_7050_53333# 1.76fF
C9255 a_20286_62194# a_20378_62194# 0.32fF
C9256 a_21382_56170# ctopp 3.40fF
C9257 a_49494_24552# m2_48260_24282# 0.60fF
C9258 a_32970_31145# a_30565_30199# 0.48fF
C9259 a_29269_40741# VDD 1.51fF
C9260 a_23390_69222# a_23390_68218# 1.00fF
C9261 vcm_commonmode a_20286_64202# 0.31fF
C9262 a_27236_50095# VDD 0.32fF
C9263 a_40458_72234# a_41462_72234# 0.97fF
C9264 a_35438_8488# a_36442_8488# 0.97fF
C9265 a_11574_22869# a_11130_22869# 0.80fF
C9266 ctopp m3_48392_55078# 0.35fF
C9267 a_34267_31599# VDD 0.40fF
C9268 a_25306_57174# a_25398_57174# 0.32fF
C9269 a_5179_74031# VDD 0.47fF
C9270 a_1770_14441# config_1_in[10] 0.60fF
C9271 a_28318_15882# a_28410_15516# 0.32fF
C9272 ctopn a_47486_21540# 3.58fF
C9273 a_2606_41079# a_3987_19623# 0.47fF
C9274 a_13183_52047# a_17366_67214# 0.38fF
C9275 a_36442_70226# a_37446_70226# 0.97fF
C9276 a_48490_19532# a_48490_18528# 1.00fF
C9277 a_13097_37455# a_14293_37455# 3.22fF
C9278 a_10515_23975# a_12895_13967# 0.93fF
C9279 a_7210_55081# a_8500_58799# 0.95fF
C9280 a_6773_27805# VDD 2.81fF
C9281 vcm_commonmode a_40458_13508# 0.87fF
C9282 a_47486_59182# a_47486_58178# 1.00fF
C9283 a_20378_61190# ctopp 3.59fF
C9284 ctopn a_24394_10496# 3.59fF
C9285 a_22386_69222# VDD 0.51fF
C9286 a_12473_36341# VDD 7.40fF
C9287 a_49494_9492# VDD 1.10fF
C9288 a_17366_16520# a_18370_16520# 0.97fF
C9289 vcm_commonmode a_26402_56170# 0.87fF
C9290 ctopn a_16746_23546# 1.42fF
C9291 a_4811_34855# a_3339_30503# 2.11fF
C9292 a_7987_15431# VDD 0.78fF
C9293 a_26310_71230# a_26402_71230# 0.32fF
C9294 vcm_commonmode a_29322_69222# 0.31fF
C9295 a_2959_47113# a_2952_46805# 0.35fF
C9296 a_49402_59182# VDD 0.31fF
C9297 a_34434_60186# a_34434_59182# 1.00fF
C9298 a_29414_22544# VDD 0.51fF
C9299 a_20378_65206# VDD 0.51fF
C9300 a_23390_63198# a_23390_62194# 1.00fF
C9301 a_38358_11866# a_38450_11500# 0.32fF
C9302 a_3949_41935# a_4578_40455# 0.47fF
C9303 a_43470_15516# a_43470_14512# 1.00fF
C9304 vcm_commonmode a_36350_22910# 0.31fF
C9305 a_24394_70226# ctopp 3.58fF
C9306 a_41462_58178# ctopp 3.59fF
C9307 a_10055_58791# a_16746_11498# 0.41fF
C9308 vcm_commonmode a_27314_65206# 0.31fF
C9309 a_36613_48169# a_12355_65103# 0.40fF
C9310 ctopn a_36629_27791# 2.62fF
C9311 a_17712_7638# a_17366_16520# 0.38fF
C9312 a_40675_27791# a_41462_16520# 0.38fF
C9313 a_28410_9492# a_28410_8488# 1.00fF
C9314 a_42374_24918# a_42466_24552# 0.32fF
C9315 a_24331_34239# VDD 0.88fF
C9316 ctopn a_19374_15516# 3.59fF
C9317 a_1803_19087# a_12473_42869# 0.97fF
C9318 vcm_commonmode a_25398_61190# 0.87fF
C9319 a_23390_67214# a_24394_67214# 0.97fF
C9320 vcm_commonmode a_12341_3311# 10.38fF
C9321 a_13183_52047# ctopp 2.36fF
C9322 a_25398_14512# VDD 0.51fF
C9323 a_41261_28335# a_42466_69222# 0.38fF
C9324 a_2872_44111# a_14985_51701# 0.65fF
C9325 a_20286_55166# VDD 0.35fF
C9326 a_16863_29415# a_41597_29967# 1.11fF
C9327 a_6515_62037# a_8491_57487# 0.43fF
C9328 a_39362_62194# a_39454_62194# 0.32fF
C9329 a_7755_26703# VDD 0.59fF
C9330 vcm_commonmode a_32334_14878# 0.31fF
C9331 ctopn a_29414_11500# 3.59fF
C9332 a_3972_25615# a_3355_25071# 0.40fF
C9333 a_38315_38053# VDD 0.82fF
C9334 a_42466_69222# a_42466_68218# 1.00fF
C9335 a_9914_68279# a_10010_68021# 0.53fF
C9336 ctopn a_33430_24552# 1.70fF
C9337 a_36328_49525# VDD 0.33fF
C9338 vcm_commonmode a_29414_70226# 0.87fF
C9339 a_6921_72943# a_2689_65103# 0.64fF
C9340 a_32426_8488# a_32426_7484# 1.00fF
C9341 a_30418_23548# VDD 0.52fF
C9342 a_42709_29199# a_48490_20536# 0.38fF
C9343 a_27406_66210# VDD 0.51fF
C9344 vcm_commonmode a_12985_16367# 6.31fF
C9345 a_44382_57174# a_44474_57174# 0.32fF
C9346 a_1761_52815# a_5915_35943# 0.83fF
C9347 a_47394_15882# a_47486_15516# 0.32fF
C9348 vcm_commonmode a_37354_23914# 0.31fF
C9349 a_7571_29199# a_18500_47491# 0.60fF
C9350 a_7755_11471# VDD 0.34fF
C9351 vcm_commonmode a_34342_66210# 0.31fF
C9352 a_25398_58178# a_26402_58178# 0.97fF
C9353 a_12869_2741# a_4443_46607# 0.91fF
C9354 a_39454_19532# VDD 0.51fF
C9355 a_32951_27247# a_12899_11471# 0.41fF
C9356 a_49494_21540# m3_49396_21402# 2.78fF
C9357 a_20378_9492# a_21382_9492# 0.97fF
C9358 a_29414_55166# m3_29316_55078# 2.81fF
C9359 a_21382_13508# a_21382_12504# 1.00fF
C9360 vcm_commonmode a_46390_19898# 0.31fF
C9361 a_30418_67214# ctopp 3.59fF
C9362 a_1761_44111# a_12663_40871# 0.67fF
C9363 a_36442_16520# a_37446_16520# 0.97fF
C9364 a_1768_16367# a_1761_35407# 0.99fF
C9365 a_45386_71230# a_45478_71230# 0.32fF
C9366 a_42709_29199# a_48490_12504# 0.38fF
C9367 a_2419_48783# VDD 6.70fF
C9368 vcm_commonmode a_47486_8488# 0.86fF
C9369 a_4758_45369# a_10503_52828# 2.83fF
C9370 a_40675_27791# a_12985_19087# 0.41fF
C9371 a_42466_63198# a_42466_62194# 1.00fF
C9372 a_1823_65853# a_4674_57685# 0.48fF
C9373 a_21371_50959# a_34482_29941# 0.46fF
C9374 vcm_commonmode a_18370_58178# 0.88fF
C9375 a_23395_52047# a_27406_59182# 0.38fF
C9376 a_2292_17179# a_1591_9839# 0.34fF
C9377 a_32611_39141# VDD 0.94fF
C9378 a_1586_66567# a_9513_65301# 0.55fF
C9379 a_14287_51175# a_6095_44807# 1.99fF
C9380 a_12516_7093# a_12983_63151# 0.67fF
C9381 a_4031_50247# a_4127_50069# 0.36fF
C9382 a_47486_9492# a_47486_8488# 1.00fF
C9383 a_47394_24918# VDD 0.35fF
C9384 a_4339_64521# a_9240_53877# 0.36fF
C9385 a_43269_29967# a_47486_20536# 0.38fF
C9386 a_35601_27497# a_11067_21583# 0.41fF
C9387 a_27535_30503# a_28757_27247# 0.47fF
C9388 a_13357_32143# VDD 2.42fF
C9389 a_33008_28853# a_28305_28879# 0.33fF
C9390 a_12899_2767# a_12899_3855# 3.61fF
C9391 a_47486_58178# a_47486_57174# 1.00fF
C9392 a_42466_67214# a_43470_67214# 0.97fF
C9393 a_16362_15516# a_12877_14441# 1.27fF
C9394 a_36613_48169# ctopp 2.62fF
C9395 a_3339_30503# a_12161_31849# 0.40fF
C9396 a_3983_12015# VDD 0.74fF
C9397 vcm_commonmode a_35438_67214# 0.87fF
C9398 a_1586_9991# a_2292_17179# 0.55fF
C9399 a_42466_20536# VDD 0.51fF
C9400 a_7755_74581# a_7921_74581# 0.42fF
C9401 a_11067_21583# a_12985_7663# 24.20fF
C9402 a_42709_29199# a_48490_17524# 0.38fF
C9403 a_43175_28335# a_12899_11471# 0.41fF
C9404 a_31422_63198# VDD 0.57fF
C9405 a_18703_29199# a_43269_29967# 0.32fF
C9406 a_49402_57174# VDD 0.31fF
C9407 vcm_commonmode a_16746_13506# 5.36fF
C9408 a_7571_26151# a_7841_12167# 0.78fF
C9409 a_24302_13874# a_24394_13508# 0.32fF
C9410 vcm_commonmode a_49402_20902# 0.30fF
C9411 a_11067_66191# a_9179_22351# 0.48fF
C9412 a_33727_39913# VDD 0.67fF
C9413 a_29322_68218# a_29414_68218# 0.32fF
C9414 a_28756_55394# a_28410_64202# 0.38fF
C9415 vcm_commonmode a_38358_63198# 0.31fF
C9416 a_22015_28111# a_13643_28327# 2.04fF
C9417 a_11067_66191# a_12757_9295# 0.33fF
C9418 a_12947_71576# a_16746_71232# 2.24fF
C9419 a_43269_29967# a_47486_12504# 0.38fF
C9420 a_25398_59182# VDD 0.51fF
C9421 a_28410_7484# a_29414_7484# 0.97fF
C9422 vcm_commonmode a_32426_9492# 0.87fF
C9423 a_7039_65469# VDD 0.50fF
C9424 a_15607_46805# a_25321_29673# 0.46fF
C9425 vcm_commonmode a_48490_16520# 0.87fF
C9426 a_29414_64202# ctopp 3.59fF
C9427 ctopn a_34434_13508# 3.59fF
C9428 vcm_commonmode a_32334_59182# 0.31fF
C9429 a_12985_19087# a_16362_9492# 1.27fF
C9430 a_4443_46607# a_2021_22325# 0.99fF
C9431 a_42466_12504# VDD 0.51fF
C9432 a_20897_42917# VDD 1.40fF
C9433 a_9503_26151# a_20378_10496# 0.38fF
C9434 a_7925_72399# a_9183_72007# 0.33fF
C9435 a_7377_18012# a_8015_20175# 0.58fF
C9436 a_3484_61493# VDD 0.32fF
C9437 a_3295_62083# a_4298_58951# 0.47fF
C9438 a_39454_9492# a_40458_9492# 0.97fF
C9439 vcm_commonmode a_49402_12870# 0.30fF
C9440 a_22386_64202# a_23390_64202# 0.97fF
C9441 a_40458_13508# a_40458_12504# 1.00fF
C9442 a_8123_34319# VDD 0.65fF
C9443 a_2840_66103# a_10680_52245# 1.25fF
C9444 a_12263_4391# a_12899_3311# 8.83fF
C9445 a_6559_22671# a_7078_36103# 0.88fF
C9446 a_13643_28327# a_37557_32463# 1.13fF
C9447 a_22015_28111# a_34062_47607# 0.63fF
C9448 a_18979_30287# VDD 11.90fF
C9449 a_31768_7638# a_31422_11500# 0.38fF
C9450 a_37446_21540# VDD 0.51fF
C9451 vcm_commonmode a_40458_7484# 0.68fF
C9452 a_43269_29967# a_47486_17524# 0.38fF
C9453 a_19374_22544# a_20378_22544# 0.97fF
C9454 a_5213_70223# VDD 0.45fF
C9455 a_38867_38591# VDD 0.86fF
C9456 vcm_commonmode a_44382_21906# 0.31fF
C9457 a_38450_69222# ctopp 3.59fF
C9458 a_2004_42453# a_3019_13621# 0.38fF
C9459 a_31768_55394# a_31422_65206# 0.38fF
C9460 vcm_commonmode a_34434_64202# 0.87fF
C9461 a_1915_35015# a_1887_34863# 0.34fF
C9462 a_42466_17524# VDD 0.51fF
C9463 a_2847_49855# VDD 0.52fF
C9464 a_46390_72234# a_46482_72234# 0.32fF
C9465 a_19374_72234# a_19374_71230# 1.00fF
C9466 a_43270_27791# a_45478_15516# 0.38fF
C9467 a_29414_60186# VDD 0.51fF
C9468 vcm_commonmode a_21290_10862# 0.31fF
C9469 a_12869_2741# a_12985_25615# 0.66fF
C9470 a_7773_63927# a_6467_55527# 0.86fF
C9471 vcm_commonmode a_49402_17890# 0.30fF
C9472 a_36442_65206# ctopp 3.59fF
C9473 a_12641_43124# a_12473_41781# 0.65fF
C9474 a_30418_67214# a_30418_66210# 1.00fF
C9475 vcm_commonmode a_36350_60186# 0.31fF
C9476 a_1950_59887# a_4148_60547# 0.61fF
C9477 a_41427_52263# a_12981_59343# 0.40fF
C9478 a_15607_46805# a_20267_30503# 0.73fF
C9479 a_6559_22671# a_6727_47607# 0.44fF
C9480 a_43362_28879# a_47486_68218# 0.38fF
C9481 a_16955_52047# a_12983_63151# 0.40fF
C9482 a_12907_56399# a_12727_67753# 0.36fF
C9483 a_4758_45369# a_4191_33449# 1.57fF
C9484 a_43270_27791# a_12899_11471# 0.41fF
C9485 a_4339_64521# a_4891_47388# 1.13fF
C9486 a_12889_39889# a_13669_39605# 1.25fF
C9487 a_26402_65206# a_26402_64202# 1.00fF
C9488 a_43378_13874# a_43470_13508# 0.32fF
C9489 vcm_commonmode a_22386_19532# 0.87fF
C9490 a_48398_68218# a_48490_68218# 0.32fF
C9491 a_17599_52263# a_12981_62313# 0.40fF
C9492 a_23395_52047# a_27406_57174# 0.38fF
C9493 a_2339_38129# a_5671_21495# 0.37fF
C9494 a_19807_28111# a_18703_29199# 1.37fF
C9495 a_37427_47893# VDD 0.94fF
C9496 a_28547_51175# a_32426_70226# 0.38fF
C9497 vcm_commonmode a_43470_69222# 0.87fF
C9498 a_1591_56623# VDD 1.02fF
C9499 a_47486_7484# a_48490_7484# 0.97fF
C9500 a_20378_23548# a_20378_22544# 1.00fF
C9501 a_2787_32679# a_2235_30503# 0.56fF
C9502 vcm_commonmode a_16362_15516# 4.47fF
C9503 a_29322_56170# a_29414_56170# 0.32fF
C9504 a_8459_71285# VDD 0.41fF
C9505 a_1761_52815# a_12713_36483# 1.07fF
C9506 a_40050_48463# a_45478_60186# 0.38fF
C9507 a_19374_11500# VDD 0.51fF
C9508 vcm_commonmode a_41462_65206# 0.87fF
C9509 a_34780_56398# a_34434_66210# 0.38fF
C9510 a_31422_69222# a_32426_69222# 0.97fF
C9511 a_39673_28111# a_40458_9492# 0.38fF
C9512 a_12473_37429# a_1761_34319# 1.11fF
C9513 a_8295_47388# a_3339_32463# 0.54fF
C9514 a_43470_18528# VDD 0.51fF
C9515 a_18611_52047# a_23390_72234# 0.34fF
C9516 a_26402_61190# a_26402_60186# 1.00fF
C9517 a_23390_24552# VDD 0.60fF
C9518 vcm_commonmode a_26310_11866# 0.31fF
C9519 ctopn a_41462_8488# 3.40fF
C9520 a_41462_64202# a_42466_64202# 0.97fF
C9521 a_1987_33402# VDD 0.51fF
C9522 a_43470_66210# ctopp 3.59fF
C9523 a_1950_59887# a_1586_51335# 0.73fF
C9524 a_25787_28327# a_33430_62194# 0.38fF
C9525 vcm_commonmode a_30326_24918# 0.31fF
C9526 a_43362_28879# a_47486_56170# 0.38fF
C9527 a_18151_52263# a_12727_67753# 0.40fF
C9528 a_38450_22544# a_39454_22544# 0.97fF
C9529 a_25269_27791# VDD 0.90fF
C9530 a_25398_57174# VDD 0.51fF
C9531 vcm_commonmode a_46482_14512# 0.87fF
C9532 a_29414_65206# a_30418_65206# 0.97fF
C9533 vcm_commonmode a_25398_20536# 0.87fF
C9534 vcm_commonmode a_40366_55166# 0.30fF
C9535 a_25398_17524# a_25398_16520# 1.00fF
C9536 vcm_commonmode a_32334_57174# 0.31fF
C9537 a_4119_70741# a_2952_66139# 1.05fF
C9538 a_4758_45369# a_12447_29199# 0.50fF
C9539 a_6559_59663# VDD 5.76fF
C9540 a_7571_29199# a_9955_20969# 0.71fF
C9541 a_20378_23548# a_21382_23548# 0.97fF
C9542 VDD dummypin[13] 0.95fF
C9543 a_29414_56170# a_29414_55166# 1.00fF
C9544 a_9637_30511# VDD 0.83fF
C9545 a_29175_28335# a_26748_7638# 0.94fF
C9546 a_14287_51175# VDD 15.15fF
C9547 a_49494_67214# a_49494_66210# 1.00fF
C9548 a_17366_66210# a_18370_66210# 0.97fF
C9549 a_8583_33551# m2_48260_54946# 0.43fF
C9550 a_42466_7484# m3_42368_7346# 2.80fF
C9551 a_16510_8760# a_9529_28335# 0.31fF
C9552 a_1761_49007# a_2021_17973# 7.18fF
C9553 a_29913_43457# VDD 1.37fF
C9554 vcm_commonmode a_48490_66210# 0.87fF
C9555 a_30573_52271# VDD 0.35fF
C9556 vcm_commonmode a_18611_52047# 10.02fF
C9557 a_39454_62194# VDD 0.51fF
C9558 a_1761_27791# a_4495_35925# 0.31fF
C9559 a_28318_61190# a_28410_61190# 0.32fF
C9560 a_39454_55166# m3_39356_55078# 2.81fF
C9561 vcm_commonmode a_25398_12504# 0.87fF
C9562 ctopn a_26402_9492# 3.58fF
C9563 a_10010_68021# VDD 0.42fF
C9564 a_45478_65206# a_45478_64202# 1.00fF
C9565 a_4351_67279# a_4482_57863# 0.88fF
C9566 ctopn a_42466_16520# 3.59fF
C9567 a_1689_10396# a_2411_26133# 0.72fF
C9568 a_9135_67503# a_9301_67503# 0.66fF
C9569 vcm_commonmode a_46390_62194# 0.31fF
C9570 a_13643_28327# a_22291_29415# 0.30fF
C9571 a_47486_15516# VDD 0.51fF
C9572 a_3031_47679# VDD 0.64fF
C9573 a_17366_71230# a_17366_70226# 1.00fF
C9574 vcm_commonmode a_17274_68218# 0.33fF
C9575 a_21371_52263# a_12901_66959# 0.40fF
C9576 a_29414_19532# a_30418_19532# 0.97fF
C9577 a_35601_27497# a_35438_13508# 0.38fF
C9578 a_39454_23548# a_39454_22544# 1.00fF
C9579 a_11067_67279# a_16362_19532# 19.89fF
C9580 a_47486_63198# ctopp 3.63fF
C9581 a_17507_52047# a_25015_48437# 0.71fF
C9582 a_16510_8760# a_12985_19087# 1.08fF
C9583 a_48398_56170# a_48490_56170# 0.32fF
C9584 a_45478_71230# VDD 0.58fF
C9585 a_1761_52815# a_15968_36061# 0.38fF
C9586 a_33430_66210# a_33430_65206# 1.00fF
C9587 a_34434_14512# a_35438_14512# 0.97fF
C9588 vcm_commonmode a_20378_21540# 0.87fF
C9589 a_13097_40719# VDD 2.29fF
C9590 VDD config_2_in[4] 1.16fF
C9591 a_27535_30503# a_20359_29199# 1.69fF
C9592 a_4127_50069# VDD 0.46fF
C9593 a_36613_48169# a_38557_32143# 0.36fF
C9594 a_45478_61190# a_45478_60186# 1.00fF
C9595 a_31330_8854# a_31422_8488# 0.32fF
C9596 a_41462_59182# ctopp 3.59fF
C9597 a_7841_22895# a_7187_23439# 0.38fF
C9598 a_26505_31599# VDD 0.78fF
C9599 vcm_commonmode a_25398_17524# 0.87fF
C9600 a_2004_42453# a_2411_26133# 0.71fF
C9601 a_7921_74581# VDD 0.67fF
C9602 a_42985_46831# a_8583_33551# 0.41fF
C9603 a_28757_27247# a_31691_32143# 0.35fF
C9604 a_34482_29941# a_18979_30287# 1.15fF
C9605 a_1586_40455# a_1761_22895# 0.43fF
C9606 a_24394_13508# VDD 0.51fF
C9607 a_18627_44581# VDD 0.79fF
C9608 a_32334_70226# a_32426_70226# 0.32fF
C9609 a_31422_62194# a_31422_61190# 1.00fF
C9610 a_22386_10496# a_22386_9492# 1.00fF
C9611 vcm_commonmode a_31330_13874# 0.31fF
C9612 a_48490_65206# a_49494_65206# 0.97fF
C9613 a_2283_15797# a_2873_13879# 0.31fF
C9614 a_44474_17524# a_44474_16520# 1.00fF
C9615 vcm_commonmode a_17274_56170# 0.33fF
C9616 a_43267_31055# a_46482_58178# 0.38fF
C9617 a_10515_22671# a_9989_46831# 1.08fF
C9618 a_31422_20536# a_31422_19532# 1.00fF
C9619 a_1586_18695# a_2143_15271# 1.87fF
C9620 a_29760_7638# a_29414_14512# 0.38fF
C9621 a_39454_23548# a_40458_23548# 0.97fF
C9622 a_8453_64757# VDD 0.60fF
C9623 a_2787_32679# a_1761_32143# 0.34fF
C9624 a_10899_28879# VDD 1.21fF
C9625 a_11067_67279# a_8295_47388# 0.66fF
C9626 a_12899_2767# a_9503_26151# 0.63fF
C9627 a_3143_22364# a_3325_18543# 1.11fF
C9628 a_46482_72234# VDD 1.35fF
C9629 vcm_commonmode a_46482_59182# 0.87fF
C9630 a_36442_66210# a_37446_66210# 0.97fF
C9631 ctopn a_16746_19530# 1.68fF
C9632 a_25971_52263# a_12355_65103# 0.40fF
C9633 a_36629_27791# a_36442_16520# 0.38fF
C9634 a_12341_3311# a_12899_11471# 0.41fF
C9635 a_7311_60975# VDD 0.32fF
C9636 a_12641_37684# a_12381_35836# 0.53fF
C9637 a_47394_61190# a_47486_61190# 0.32fF
C9638 a_45478_60186# ctopp 3.59fF
C9639 a_32951_27247# a_33430_23548# 0.36fF
C9640 a_48490_68218# VDD 0.54fF
C9641 vcm_commonmode a_26402_18528# 0.87fF
C9642 a_48398_7850# VDD 0.62fF
C9643 vcm_commonmode a_16746_61192# 5.36fF
C9644 a_19282_67214# a_19374_67214# 0.32fF
C9645 ctopn a_44474_22544# 3.58fF
C9646 a_2012_33927# a_2223_28617# 0.65fF
C9647 a_7695_31573# a_7281_29423# 0.38fF
C9648 a_34482_29941# a_37427_47893# 0.59fF
C9649 a_4191_33449# a_12447_29199# 1.12fF
C9650 a_38557_32143# a_38450_69222# 0.38fF
C9651 a_36442_71230# a_36442_70226# 1.00fF
C9652 a_48490_19532# a_49494_19532# 0.97fF
C9653 a_12341_3311# a_22386_13508# 0.38fF
C9654 a_17366_62194# ctopp 3.43fF
C9655 a_19780_38341# VDD 1.50fF
C9656 a_11067_67279# a_17712_7638# 0.40fF
C9657 a_32795_29967# a_26523_29199# 0.34fF
C9658 a_16101_31029# a_15799_29941# 0.49fF
C9659 a_1586_9991# a_3327_9308# 0.48fF
C9660 a_19675_49525# VDD 0.39fF
C9661 vcm_commonmode a_20286_70226# 0.31fF
C9662 a_32426_20536# a_33430_20536# 0.97fF
C9663 a_37354_58178# vcm_commonmode 0.31fF
C9664 vcm_commonmode a_35438_10496# 0.87fF
C9665 a_9135_27239# a_12985_7663# 0.41fF
C9666 a_3339_32463# a_1915_35015# 0.36fF
C9667 a_21382_63198# a_22386_63198# 0.97fF
C9668 a_8197_31599# VDD 1.73fF
C9669 ctopn a_40458_14512# 3.59fF
C9670 a_2317_28892# a_3325_18543# 0.65fF
C9671 a_1768_16367# a_1823_65853# 0.61fF
C9672 a_23390_71230# ctopp 3.40fF
C9673 ctopn a_19374_20536# 3.59fF
C9674 a_2012_33927# a_3301_26703# 0.90fF
C9675 a_30788_28487# a_19626_31751# 0.30fF
C9676 a_2847_12863# VDD 0.51fF
C9677 a_33727_44265# VDD 0.66fF
C9678 a_21290_58178# a_21382_58178# 0.32fF
C9679 a_2939_52245# VDD 0.39fF
C9680 a_16746_61192# a_16362_61190# 2.28fF
C9681 a_41462_10496# a_41462_9492# 1.00fF
C9682 a_40675_27791# VDD 6.51fF
C9683 a_22386_55166# m3_22288_55078# 2.81fF
C9684 a_48490_56170# VDD 0.56fF
C9685 a_6515_62037# a_7479_54439# 0.33fF
C9686 a_2021_17973# a_27359_43985# 0.33fF
C9687 a_31422_8488# VDD 0.58fF
C9688 vcm_commonmode a_22386_62194# 0.87fF
C9689 a_32334_16886# a_32426_16520# 0.32fF
C9690 ctopn a_45478_23548# 3.40fF
C9691 a_1643_57685# VDD 0.37fF
C9692 vcm_commonmode a_38358_8854# 0.31fF
C9693 m3_26304_7346# VDD 0.33fF
C9694 a_23736_7638# a_23390_16520# 0.38fF
C9695 a_49402_65206# VDD 0.31fF
C9696 vcm_commonmode a_30418_15516# 0.87fF
C9697 ctopn a_19374_12504# 3.59fF
C9698 a_43267_31055# a_13643_28327# 0.48fF
C9699 a_41462_57174# ctopp 3.58fF
C9700 a_18611_52047# a_23390_59182# 0.38fF
C9701 a_16043_38825# VDD 0.51fF
C9702 a_13349_37973# VDD 2.83fF
C9703 a_25744_7638# a_25398_9492# 0.38fF
C9704 a_8491_27023# a_18370_9492# 0.38fF
C9705 ctopn a_29760_7638# 2.62fF
C9706 vcm_commonmode a_28410_71230# 0.86fF
C9707 a_30418_21540# a_30418_20536# 1.00fF
C9708 a_5671_21495# a_10394_19605# 0.76fF
C9709 a_47486_61190# VDD 0.51fF
C9710 a_12907_27023# a_17712_7638# 1.51fF
C9711 a_18979_30287# a_36904_28879# 0.35fF
C9712 a_17366_55166# a_18370_55166# 0.97fF
C9713 vcm_commonmode a_40458_11500# 0.87fF
C9714 a_17366_24552# a_17366_23548# 1.00fF
C9715 a_35601_27497# a_12546_22351# 0.41fF
C9716 a_19374_67214# VDD 0.51fF
C9717 a_32426_12504# a_33430_12504# 0.97fF
C9718 a_38358_67214# a_38450_67214# 0.32fF
C9719 vcm_commonmode a_44474_24552# 0.84fF
C9720 a_25971_52263# ctopp 2.62fF
C9721 a_7862_34025# a_25263_29981# 0.63fF
C9722 a_22399_32143# a_23395_32463# 0.34fF
C9723 vcm_commonmode a_26310_67214# 0.31fF
C9724 a_2775_46025# a_28881_52271# 0.61fF
C9725 a_15599_28585# VDD 0.48fF
C9726 a_26402_68218# ctopp 3.59fF
C9727 ctopn a_19374_17524# 3.59fF
C9728 a_16362_9492# VDD 2.47fF
C9729 a_16265_39868# VDD 1.02fF
C9730 a_18151_52263# a_24394_64202# 0.38fF
C9731 a_2292_17179# a_5805_15279# 0.61fF
C9732 a_35601_27497# a_35438_7484# 0.34fF
C9733 vcm_commonmode a_46482_57174# 0.87fF
C9734 a_32426_16520# VDD 0.51fF
C9735 a_12901_58799# VDD 6.95fF
C9736 a_24302_7850# a_24394_7484# 0.32fF
C9737 vcm_commonmode a_23298_9858# 0.31fF
C9738 a_40458_63198# a_41462_63198# 0.97fF
C9739 vcm_commonmode a_39362_16886# 0.31fF
C9740 a_25269_27791# a_24740_7638# 0.36fF
C9741 a_27406_21540# a_28410_21540# 0.97fF
C9742 a_35346_9858# a_35438_9492# 0.32fF
C9743 a_18278_64202# a_18370_64202# 0.32fF
C9744 a_24394_7484# VDD 1.24fF
C9745 a_45478_58178# a_46482_58178# 0.97fF
C9746 vcm_commonmode a_31422_68218# 0.87fF
C9747 a_34434_59182# a_35438_59182# 0.97fF
C9748 a_25744_7638# a_12985_19087# 0.41fF
C9749 a_18370_64202# VDD 0.52fF
C9750 a_12355_15055# a_7187_23439# 0.95fF
C9751 a_41967_31375# a_11067_21583# 0.41fF
C9752 a_26402_56170# ctopp 3.40fF
C9753 a_18731_38825# VDD 0.62fF
C9754 ctopn a_20378_18528# 3.59fF
C9755 a_23395_52047# a_27406_65206# 0.38fF
C9756 vcm_commonmode a_25306_64202# 0.31fF
C9757 a_32426_17524# a_33430_17524# 0.97fF
C9758 a_26662_48981# VDD 1.01fF
C9759 a_49494_21540# a_49494_20536# 1.00fF
C9760 a_19374_60186# a_20378_60186# 0.97fF
C9761 a_36442_24552# a_36442_23548# 1.00fF
C9762 a_27535_30503# a_28446_31375# 0.75fF
C9763 a_21382_12504# a_21382_11500# 1.00fF
C9764 a_40139_32143# VDD 0.38fF
C9765 ctopn a_16746_14510# 1.68fF
C9766 a_9314_69367# VDD 2.10fF
C9767 a_34780_56398# a_12981_59343# 0.40fF
C9768 a_7571_26151# a_7571_29199# 1.51fF
C9769 a_41872_29423# a_43470_68218# 0.38fF
C9770 a_7050_53333# VDD 6.18fF
C9771 a_5671_21495# a_5535_18012# 2.02fF
C9772 vcm_commonmode a_45478_13508# 0.87fF
C9773 a_25398_61190# ctopp 3.59fF
C9774 ctopn a_29414_10496# 3.59fF
C9775 a_27406_69222# VDD 0.51fF
C9776 a_4275_36201# VDD 0.39fF
C9777 a_34222_43439# a_2021_17973# 1.18fF
C9778 a_1761_44111# a_19410_43439# 0.95fF
C9779 a_12341_3311# a_22386_7484# 0.34fF
C9780 a_18611_52047# a_23390_57174# 0.38fF
C9781 vcm_commonmode a_31422_56170# 0.87fF
C9782 a_10791_15529# VDD 0.62fF
C9783 vcm_commonmode a_34342_69222# 0.31fF
C9784 a_28756_55394# a_28410_70226# 0.38fF
C9785 a_42985_46831# a_12516_7093# 0.40fF
C9786 a_24740_7638# a_24394_13508# 0.38fF
C9787 a_43378_7850# a_43470_7484# 0.32fF
C9788 a_34434_22544# VDD 0.51fF
C9789 a_6095_44807# a_1586_45431# 0.44fF
C9790 a_43270_27791# a_45478_20536# 0.38fF
C9791 a_25398_65206# VDD 0.51fF
C9792 a_2840_66103# a_6095_44807# 0.43fF
C9793 a_41427_52263# a_41462_60186# 0.38fF
C9794 vcm_commonmode a_41370_22910# 0.31fF
C9795 a_29414_70226# ctopp 3.58fF
C9796 a_10531_31055# a_14625_30761# 0.39fF
C9797 a_1761_49007# a_37939_43455# 0.73fF
C9798 vcm_commonmode a_32334_65206# 0.31fF
C9799 a_25971_52263# a_30418_66210# 0.38fF
C9800 a_27314_69222# a_27406_69222# 0.32fF
C9801 a_33430_18528# a_33430_17524# 1.00fF
C9802 a_46482_21540# a_47486_21540# 0.97fF
C9803 a_8569_24527# VDD 0.84fF
C9804 vcm_commonmode a_16746_11498# 5.36fF
C9805 a_33864_28111# a_11067_21583# 0.41fF
C9806 a_7111_22351# a_5839_22351# 0.40fF
C9807 a_37354_64202# a_37446_64202# 0.32fF
C9808 ctopn a_24394_15516# 3.59fF
C9809 a_21371_50959# a_25419_50959# 3.81fF
C9810 a_1761_6031# VDD 0.54fF
C9811 a_9599_57141# a_9135_56623# 0.30fF
C9812 vcm_commonmode a_30418_61190# 0.87fF
C9813 a_29760_55394# a_29414_62194# 0.38fF
C9814 a_41872_29423# a_43470_56170# 0.38fF
C9815 a_7939_30503# a_14926_31849# 2.46fF
C9816 a_30418_14512# VDD 0.51fF
C9817 a_43270_27791# a_45478_12504# 0.38fF
C9818 a_12901_58799# a_16746_58180# 2.28fF
C9819 a_11067_47695# a_4191_33449# 1.49fF
C9820 a_8015_20175# VDD 0.42fF
C9821 a_25306_55166# VDD 0.35fF
C9822 a_34342_22910# a_34434_22544# 0.32fF
C9823 a_43175_28335# a_46482_18528# 0.38fF
C9824 a_6816_19355# a_4792_20443# 0.36fF
C9825 a_23390_10496# a_24394_10496# 0.97fF
C9826 a_12947_56817# VDD 3.62fF
C9827 vcm_commonmode a_37354_14878# 0.31fF
C9828 ctopn a_34434_11500# 3.59fF
C9829 a_19919_38695# a_12663_39783# 0.63fF
C9830 a_25306_65206# a_25398_65206# 0.32fF
C9831 a_34434_14512# a_34434_13508# 1.00fF
C9832 a_21187_29415# a_19807_28111# 6.79fF
C9833 vcm_commonmode a_34434_70226# 0.87fF
C9834 a_8295_47388# a_1586_18695# 0.62fF
C9835 a_38450_60186# a_39454_60186# 0.97fF
C9836 a_35438_23548# VDD 0.52fF
C9837 a_18370_58178# ctopp 3.58fF
C9838 a_32951_27247# a_12985_7663# 0.41fF
C9839 a_32426_66210# VDD 0.51fF
C9840 a_40458_12504# a_40458_11500# 1.00fF
C9841 a_38076_31573# VDD 0.32fF
C9842 a_1761_43567# a_3759_39991# 0.62fF
C9843 vcm_commonmode a_42374_23914# 0.31fF
C9844 a_35438_7484# m3_35340_7346# 2.80fF
C9845 vcm_commonmode a_39362_66210# 0.31fF
C9846 a_5682_69367# a_3024_67191# 0.35fF
C9847 a_27406_70226# a_27406_69222# 1.00fF
C9848 a_33430_18528# a_34434_18528# 0.97fF
C9849 a_44474_19532# VDD 0.51fF
C9850 a_2411_19605# a_4241_18543# 0.62fF
C9851 a_43270_27791# a_45478_17524# 0.38fF
C9852 a_20267_30503# a_30565_30199# 1.49fF
C9853 a_3339_43023# a_27535_30503# 0.32fF
C9854 a_6646_54135# VDD 0.74fF
C9855 a_42709_29199# a_11067_21583# 0.40fF
C9856 a_1959_68053# VDD 0.49fF
C9857 a_16510_8760# VDD 6.14fF
C9858 a_35438_67214# ctopp 3.59fF
C9859 a_5831_39189# a_1761_40847# 0.80fF
C9860 a_19720_55394# a_12901_66959# 0.40fF
C9861 a_6224_73095# a_5024_67885# 0.33fF
C9862 a_25306_19898# a_25398_19532# 0.32fF
C9863 a_16362_58178# VDD 2.48fF
C9864 a_8583_33551# a_1761_22895# 0.82fF
C9865 a_26402_11500# a_26402_10496# 1.00fF
C9866 vcm_commonmode a_23390_58178# 0.87fF
C9867 a_30326_14878# a_30418_14512# 0.32fF
C9868 a_42188_37149# VDD 2.45fF
C9869 a_49876_41198# VDD 4.78fF
C9870 a_46390_69222# a_46482_69222# 0.32fF
C9871 a_12621_36091# a_12549_35836# 0.37fF
C9872 a_27869_50095# VDD 4.02fF
C9873 a_33430_72234# a_34434_72234# 0.97fF
C9874 a_2511_60431# VDD 0.43fF
C9875 a_5363_30503# a_13357_32143# 0.68fF
C9876 a_24394_55166# a_25398_55166# 0.97fF
C9877 a_42709_29199# a_48490_21540# 0.38fF
C9878 a_43175_28335# a_12985_7663# 0.41fF
C9879 a_9503_26151# a_11067_21583# 0.41fF
C9880 vcm_commonmode a_16362_17524# 4.47fF
C9881 a_13067_38517# a_13909_41923# 3.94fF
C9882 a_28547_51175# a_2959_47113# 0.87fF
C9883 a_18370_15516# a_19374_15516# 0.97fF
C9884 vcm_commonmode a_40458_67214# 0.87fF
C9885 a_31768_7638# a_31422_10496# 0.38fF
C9886 a_47486_20536# VDD 0.51fF
C9887 a_1768_16367# a_1778_42631# 0.88fF
C9888 a_36442_63198# VDD 0.57fF
C9889 a_4685_37583# a_5915_30287# 0.95fF
C9890 a_42466_10496# a_43470_10496# 0.97fF
C9891 a_33864_28111# a_34434_24552# 0.43fF
C9892 a_9319_69141# VDD 0.48fF
C9893 a_44382_65206# a_44474_65206# 0.32fF
C9894 vcm_commonmode a_43378_63198# 0.31fF
C9895 a_27869_50095# a_26514_47375# 0.31fF
C9896 a_18703_29199# VDD 10.83fF
C9897 a_30418_59182# VDD 0.51fF
C9898 vcm_commonmode a_37446_9492# 0.87fF
C9899 m3_16264_69134# VDD 0.34fF
C9900 a_35346_23914# a_35438_23548# 0.32fF
C9901 a_12869_2741# a_12349_25847# 1.43fF
C9902 a_28410_11500# a_29414_11500# 0.97fF
C9903 a_34434_64202# ctopp 3.59fF
C9904 ctopn a_39454_13508# 3.59fF
C9905 a_39454_72234# VDD 1.23fF
C9906 vcm_commonmode a_37354_59182# 0.31fF
C9907 a_41261_28335# a_12727_58255# 0.40fF
C9908 a_32334_66210# a_32426_66210# 0.32fF
C9909 vcm_commonmode a_17366_22544# 1.82fF
C9910 a_33798_31145# a_32970_31145# 0.32fF
C9911 vcm_commonmode m3_16264_59094# 3.21fF
C9912 a_47486_12504# VDD 0.51fF
C9913 a_29483_42943# VDD 0.82fF
C9914 a_46482_70226# a_46482_69222# 1.00fF
C9915 a_18611_52047# a_12355_65103# 0.44fF
C9916 a_2099_59861# a_2411_26133# 0.70fF
C9917 a_14983_51157# a_17682_50095# 0.33fF
C9918 vcm_commonmode a_44474_72234# 0.69fF
C9919 a_12355_15055# a_8566_39215# 3.02fF
C9920 a_4891_47388# a_8295_47388# 0.76fF
C9921 a_1768_13103# a_1586_9991# 1.51fF
C9922 a_43269_29967# a_47486_21540# 0.38fF
C9923 a_32426_24552# a_33430_24552# 0.97fF
C9924 a_19743_34743# VDD 0.61fF
C9925 vcm_commonmode a_17274_18894# 0.33fF
C9926 ctopn a_12727_15529# 3.23fF
C9927 a_42985_46831# a_48490_63198# 0.42fF
C9928 a_4811_34855# a_14926_31849# 0.36fF
C9929 a_19807_28111# a_26523_28111# 0.85fF
C9930 a_8117_12559# VDD 0.75fF
C9931 a_3339_43023# inn_analog 2.70fF
C9932 a_34780_56398# a_34434_69222# 0.38fF
C9933 a_44382_19898# a_44474_19532# 0.32fF
C9934 a_42466_21540# VDD 0.51fF
C9935 vcm_commonmode a_45478_7484# 0.69fF
C9936 a_28756_7638# a_28410_18528# 0.38fF
C9937 a_4674_40277# a_5547_31599# 0.43fF
C9938 a_29414_62194# a_30418_62194# 0.97fF
C9939 a_45478_11500# a_45478_10496# 1.00fF
C9940 a_7637_69679# VDD 0.46fF
C9941 a_49402_14878# a_49494_14512# 0.32fF
C9942 a_4227_37887# VDD 0.56fF
C9943 vcm_commonmode a_49402_21906# 0.30fF
C9944 a_43470_69222# ctopp 3.59fF
C9945 a_19374_10496# VDD 0.51fF
C9946 a_19245_39747# VDD 0.80fF
C9947 vcm_commonmode a_39454_64202# 0.87fF
C9948 a_24740_7638# a_24394_7484# 0.35fF
C9949 a_1586_9991# a_4812_13879# 0.53fF
C9950 a_12473_36341# a_31959_34751# 0.33fF
C9951 a_47486_17524# VDD 0.51fF
C9952 a_1586_45431# VDD 6.54fF
C9953 a_42985_46831# a_48490_72234# 0.35fF
C9954 a_28318_20902# a_28410_20536# 0.32fF
C9955 a_9503_26151# a_20378_15516# 0.38fF
C9956 a_34434_60186# VDD 0.51fF
C9957 a_42466_55166# a_43470_55166# 0.97fF
C9958 a_5991_21263# VDD 0.37fF
C9959 vcm_commonmode a_26310_10862# 0.31fF
C9960 a_43270_27791# a_12985_7663# 0.41fF
C9961 a_7187_23439# a_8933_22583# 0.36fF
C9962 a_2840_66103# VDD 17.89fF
C9963 a_11067_46823# a_28757_27247# 0.55fF
C9964 a_2787_32679# a_4495_35925# 0.36fF
C9965 a_17274_63198# a_17366_63198# 0.32fF
C9966 a_6515_62037# a_6559_59879# 0.65fF
C9967 a_41462_65206# ctopp 3.59fF
C9968 a_28817_29111# a_29175_28335# 0.30fF
C9969 a_12357_37999# a_26417_40193# 0.51fF
C9970 a_34434_57174# a_35438_57174# 0.97fF
C9971 a_1643_72917# VDD 0.37fF
C9972 vcm_commonmode a_41370_60186# 0.31fF
C9973 a_37446_15516# a_38450_15516# 0.97fF
C9974 vcm_commonmode a_18370_23548# 0.88fF
C9975 a_11803_55311# a_12755_53030# 0.53fF
C9976 a_25321_29673# a_25263_29981# 0.47fF
C9977 a_13005_43983# VDD 1.46fF
C9978 a_35601_27497# a_35438_11500# 0.38fF
C9979 a_16746_58180# a_16362_58178# 2.28fF
C9980 a_3295_62083# VDD 6.21fF
C9981 a_20267_30503# a_26523_29199# 1.07fF
C9982 vcm_commonmode a_27406_19532# 0.87fF
C9983 a_37446_58178# a_37446_59182# 1.00fF
C9984 a_25787_28327# a_12869_2741# 0.49fF
C9985 a_11803_55311# a_12355_15055# 1.09fF
C9986 a_4811_34855# a_9367_29397# 0.82fF
C9987 a_21187_29415# a_29927_29199# 1.91fF
C9988 a_13643_28327# a_12907_27023# 7.94fF
C9989 a_35438_71230# a_36442_71230# 0.97fF
C9990 vcm_commonmode a_48490_69222# 0.87fF
C9991 m3_16264_16382# VDD 0.35fF
C9992 a_47486_11500# a_48490_11500# 0.97fF
C9993 vcm_commonmode a_21290_15882# 0.31fF
C9994 a_19720_55394# a_19374_59182# 0.38fF
C9995 a_49750_39288# VDD 0.40fF
C9996 a_19374_72234# m3_19276_72146# 2.80fF
C9997 a_13353_30511# a_18162_31055# 0.73fF
C9998 a_24394_11500# VDD 0.51fF
C9999 a_4960_40847# VDD 0.92fF
C10000 vcm_commonmode a_46482_65206# 0.87fF
C10001 a_12713_36483# a_12381_35836# 0.97fF
C10002 a_29055_49525# a_27869_50095# 0.60fF
C10003 a_48490_18528# VDD 0.54fF
C10004 vcm_commonmode a_19282_71230# 0.31fF
C10005 a_28410_24552# VDD 0.60fF
C10006 vcm_commonmode a_31330_11866# 0.31fF
C10007 ctopn a_46482_8488# 3.40fF
C10008 a_1586_21959# a_2143_15271# 0.72fF
C10009 a_12355_15055# a_12981_62313# 23.96fF
C10010 a_28318_12870# a_28410_12504# 0.32fF
C10011 a_3417_33231# VDD 1.09fF
C10012 a_48490_66210# ctopp 3.43fF
C10013 vcm_commonmode a_35346_24918# 0.31fF
C10014 a_18611_52047# ctopp 2.62fF
C10015 vcm_commonmode a_16362_67214# 4.47fF
C10016 a_41967_31375# a_42466_8488# 0.38fF
C10017 a_23390_59182# a_23390_58178# 1.00fF
C10018 a_38450_55166# VDD 0.60fF
C10019 a_48490_62194# a_49494_62194# 0.97fF
C10020 a_30418_57174# VDD 0.51fF
C10021 a_7841_12167# a_9083_13879# 0.51fF
C10022 vcm_commonmode a_30418_20536# 0.87fF
C10023 vcm_commonmode a_45386_55166# 0.30fF
C10024 a_5259_39367# VDD 0.58fF
C10025 a_19374_68218# a_20378_68218# 0.97fF
C10026 vcm_commonmode a_19374_63198# 0.92fF
C10027 a_16955_52047# a_20378_64202# 0.38fF
C10028 vcm_commonmode a_37354_57174# 0.31fF
C10029 a_17682_50095# a_28108_48463# 0.81fF
C10030 a_11067_23759# a_12947_8725# 0.30fF
C10031 a_47394_20902# a_47486_20536# 0.32fF
C10032 a_14287_51175# a_5363_30503# 0.81fF
C10033 a_23736_7638# a_12877_16911# 0.41fF
C10034 a_36350_63198# a_36442_63198# 0.32fF
C10035 a_27406_57174# a_27406_56170# 1.00fF
C10036 a_30412_42589# VDD 2.22fF
C10037 a_12341_3311# a_22386_11500# 0.38fF
C10038 a_26748_7638# a_26402_9492# 0.38fF
C10039 a_10975_66407# a_9484_11989# 0.63fF
C10040 a_12755_51562# VDD 1.19fF
C10041 a_2843_71829# a_2747_72007# 0.45fF
C10042 a_23298_21906# a_23390_21540# 0.32fF
C10043 a_44474_62194# VDD 0.51fF
C10044 a_25744_7638# VDD 6.49fF
C10045 vcm_commonmode a_30418_12504# 0.87fF
C10046 ctopn a_31422_9492# 3.58fF
C10047 a_4351_67279# a_10957_57711# 0.37fF
C10048 ctopn a_47486_16520# 3.58fF
C10049 a_1761_25071# a_2411_26133# 1.33fF
C10050 vcm_commonmode a_3339_43023# 2.52fF
C10051 a_34482_29941# a_18703_29199# 0.56fF
C10052 a_4191_33449# a_18539_47617# 0.33fF
C10053 vcm_commonmode a_22294_68218# 0.31fF
C10054 a_30326_59182# a_30418_59182# 0.32fF
C10055 a_37919_28111# a_38450_19532# 0.38fF
C10056 a_18979_30287# a_23395_32463# 0.47fF
C10057 a_10515_63143# a_12341_3311# 1.49fF
C10058 a_41967_31375# a_12546_22351# 0.41fF
C10059 a_1761_50639# a_12473_37429# 1.07fF
C10060 vcm_commonmode a_25398_21540# 0.87fF
C10061 a_11067_67279# a_11619_3303# 1.14fF
C10062 a_1761_50639# a_20713_40193# 0.62fF
C10063 a_3413_10389# VDD 0.63fF
C10064 a_19743_41271# VDD 0.61fF
C10065 a_18611_52047# a_23390_65206# 0.38fF
C10066 a_28318_17890# a_28410_17524# 0.32fF
C10067 a_14831_50095# VDD 5.15fF
C10068 a_39362_72234# a_39454_72234# 0.32fF
C10069 a_36797_27497# a_12727_15529# 0.41fF
C10070 a_5363_30503# a_26505_31599# 0.42fF
C10071 a_31422_55166# a_32426_55166# 0.97fF
C10072 a_46482_59182# ctopp 3.59fF
C10073 a_1586_36727# a_1591_38677# 0.72fF
C10074 a_34434_64202# a_34434_63198# 1.23fF
C10075 a_47394_12870# a_47486_12504# 0.32fF
C10076 vcm_commonmode a_30418_17524# 0.87fF
C10077 a_23395_52047# a_12981_59343# 0.40fF
C10078 vcm_commonmode a_17366_60186# 1.83fF
C10079 a_5682_69367# a_9828_56311# 0.31fF
C10080 a_9307_30663# a_8197_31599# 0.42fF
C10081 a_29927_29199# a_26523_28111# 0.98fF
C10082 a_29414_13508# VDD 0.51fF
C10083 a_37446_58178# a_37446_57174# 1.00fF
C10084 a_27183_44581# VDD 0.88fF
C10085 a_39389_52271# a_39454_68218# 0.38fF
C10086 a_2012_33927# a_2473_34293# 0.32fF
C10087 a_1757_19631# VDD 0.62fF
C10088 a_5179_74031# a_5345_74031# 0.68fF
C10089 a_6831_63303# a_7387_46831# 0.43fF
C10090 a_26402_22544# a_26402_21540# 1.00fF
C10091 a_2315_24540# VDD 2.62fF
C10092 vcm_commonmode a_36350_13874# 0.31fF
C10093 a_16746_61192# ctopp 1.68fF
C10094 a_33430_13508# a_34434_13508# 0.97fF
C10095 a_1761_30511# VDD 7.38fF
C10096 a_5831_39189# a_8540_42167# 0.30fF
C10097 a_38450_68218# a_39454_68218# 0.97fF
C10098 vcm_commonmode a_22294_56170# 0.31fF
C10099 a_19720_55394# a_19374_57174# 0.38fF
C10100 a_19333_48463# VDD 0.38fF
C10101 a_41427_52263# a_12516_7093# 0.40fF
C10102 a_18151_52263# a_24394_70226# 0.38fF
C10103 a_32951_27247# a_33430_14512# 0.38fF
C10104 a_8583_33551# a_12447_29199# 1.29fF
C10105 a_12341_3311# a_12985_7663# 0.45fF
C10106 a_49876_41198# a_50198_39208# 0.60fF
C10107 a_19967_41781# a_18127_35797# 0.30fF
C10108 a_46482_57174# a_46482_56170# 1.00fF
C10109 a_19374_56170# a_20378_56170# 0.97fF
C10110 a_11067_67279# a_11145_60431# 0.45fF
C10111 a_36613_48169# a_37446_60186# 0.38fF
C10112 ctopn a_21382_19532# 3.59fF
C10113 a_1761_47919# a_12725_44527# 0.82fF
C10114 a_21371_52263# a_26402_66210# 0.38fF
C10115 ctopn a_19720_7638# 2.62fF
C10116 a_19946_51157# VDD 0.79fF
C10117 a_1586_69367# a_1591_71317# 0.80fF
C10118 a_42374_21906# a_42466_21540# 0.32fF
C10119 a_35601_27497# a_12985_16367# 0.41fF
C10120 a_12907_27023# a_11619_3303# 0.37fF
C10121 a_26523_28111# a_28817_29111# 0.65fF
C10122 a_49494_20536# m3_49396_20398# 2.78fF
C10123 a_23390_58178# a_23390_57174# 1.00fF
C10124 a_33864_28111# a_12546_22351# 0.41fF
C10125 a_6559_22671# a_4495_35925# 0.65fF
C10126 vcm_commonmode a_31422_18528# 0.87fF
C10127 vcm_commonmode a_21290_61190# 0.31fF
C10128 a_21371_50959# a_25398_62194# 0.38fF
C10129 a_7987_15431# a_7959_15279# 0.38fF
C10130 a_30418_16520# a_30418_15516# 1.00fF
C10131 a_39389_52271# a_39454_56170# 0.38fF
C10132 a_1689_10396# a_2292_17179# 1.12fF
C10133 a_3339_43023# a_3162_43023# 0.35fF
C10134 a_49402_59182# a_49494_59182# 0.32fF
C10135 a_1768_13103# config_2_in[6] 0.64fF
C10136 a_40491_27247# a_43470_19532# 0.38fF
C10137 a_19282_10862# a_19374_10496# 0.32fF
C10138 a_22386_62194# ctopp 3.59fF
C10139 a_18370_70226# VDD 0.52fF
C10140 a_30127_38053# VDD 0.93fF
C10141 vcm_commonmode a_22386_55166# 0.84fF
C10142 VDD result_out[8] 0.76fF
C10143 a_47394_17890# a_47486_17524# 0.32fF
C10144 vcm_commonmode a_12257_56623# 6.21fF
C10145 a_20359_29199# a_11067_46823# 2.46fF
C10146 a_2899_16367# VDD 0.42fF
C10147 a_2686_70223# a_2689_65103# 0.33fF
C10148 vcm_commonmode a_25306_70226# 0.31fF
C10149 a_42374_58178# vcm_commonmode 0.31fF
C10150 a_5363_30503# a_8197_31599# 0.40fF
C10151 a_34342_60186# a_34434_60186# 0.32fF
C10152 vcm_commonmode a_40458_10496# 0.87fF
C10153 a_1803_19087# a_2012_33927# 0.35fF
C10154 ctopn a_45478_14512# 3.59fF
C10155 a_17222_27247# a_15681_27497# 0.66fF
C10156 a_28410_71230# ctopp 3.40fF
C10157 ctopn a_24394_20536# 3.59fF
C10158 a_28410_7484# m3_28312_7346# 2.80fF
C10159 a_2787_30503# a_8753_31055# 0.60fF
C10160 a_1591_43029# VDD 0.59fF
C10161 a_29322_18894# a_29414_18528# 0.32fF
C10162 a_14293_37455# a_13576_37149# 2.47fF
C10163 a_2872_44111# a_19531_49007# 0.41fF
C10164 a_2021_22325# config_1_in[13] 0.59fF
C10165 a_45478_22544# a_45478_21540# 1.00fF
C10166 a_2021_22325# a_5441_27791# 0.42fF
C10167 a_18370_61190# a_19374_61190# 0.97fF
C10168 a_11711_27247# VDD 0.32fF
C10169 a_42709_29199# a_12546_22351# 0.40fF
C10170 a_36442_8488# VDD 0.58fF
C10171 vcm_commonmode a_27406_62194# 0.87fF
C10172 a_24394_68218# a_24394_67214# 1.00fF
C10173 a_11067_21583# a_12727_13353# 0.30fF
C10174 a_7467_57863# VDD 0.55fF
C10175 vcm_commonmode a_43378_8854# 0.31fF
C10176 m3_41364_7346# VDD 0.42fF
C10177 a_36629_27791# a_12985_19087# 0.41fF
C10178 vcm_commonmode a_35438_15516# 0.87fF
C10179 ctopn a_24394_12504# 3.59fF
C10180 a_17599_52263# a_12907_27023# 1.06fF
C10181 a_38450_56170# a_39454_56170# 0.97fF
C10182 a_46482_57174# ctopp 3.58fF
C10183 a_43362_28879# a_10515_22671# 0.40fF
C10184 a_16362_17524# a_12899_11471# 1.27fF
C10185 ctopn a_40491_27247# 2.63fF
C10186 a_17493_50639# VDD 0.92fF
C10187 vcm_commonmode a_33430_71230# 0.86fF
C10188 a_25971_52263# a_31768_55394# 0.31fF
C10189 a_29760_55394# a_28547_51175# 0.40fF
C10190 a_20286_55166# a_20378_55166# 0.32fF
C10191 a_21382_8488# a_22386_8488# 0.97fF
C10192 vcm_commonmode a_45478_11500# 0.87fF
C10193 a_9503_26151# a_12546_22351# 0.41fF
C10194 a_3339_43023# a_6816_19355# 1.13fF
C10195 a_24394_67214# VDD 0.51fF
C10196 a_10515_32143# VDD 0.40fF
C10197 a_6831_63303# a_6835_46823# 2.01fF
C10198 a_21371_50959# a_2959_47113# 0.42fF
C10199 a_13183_52047# a_17366_61190# 0.38fF
C10200 a_49494_16520# a_49494_15516# 1.00fF
C10201 ctopn a_19374_21540# 3.59fF
C10202 a_22386_70226# a_23390_70226# 0.97fF
C10203 vcm_commonmode a_31330_67214# 0.31fF
C10204 a_24740_7638# a_24394_11500# 0.38fF
C10205 a_34434_19532# a_34434_18528# 1.00fF
C10206 a_13909_37571# a_13097_37455# 0.48fF
C10207 a_39454_58178# a_40458_58178# 0.97fF
C10208 a_38358_10862# a_38450_10496# 0.32fF
C10209 a_29175_28335# VDD 6.75fF
C10210 a_31422_68218# ctopp 3.59fF
C10211 ctopn a_24394_17524# 3.59fF
C10212 a_21382_9492# VDD 0.51fF
C10213 a_27267_39605# VDD 0.43fF
C10214 a_37446_16520# VDD 0.51fF
C10215 a_20378_60186# a_20378_59182# 1.00fF
C10216 vcm_commonmode a_28318_9858# 0.31fF
C10217 m3_26304_72146# VDD 0.33fF
C10218 a_10515_23975# a_11067_21583# 24.00fF
C10219 a_5831_39189# a_1761_34319# 0.40fF
C10220 a_24302_11866# a_24394_11500# 0.32fF
C10221 vcm_commonmode a_44382_16886# 0.31fF
C10222 a_12473_41781# a_13909_41923# 1.14fF
C10223 a_32426_72234# VDD 1.25fF
C10224 a_34251_52263# a_12727_58255# 0.40fF
C10225 a_29414_15516# a_29414_14512# 1.00fF
C10226 a_1761_49007# a_27359_43985# 0.64fF
C10227 a_48398_18894# a_48490_18528# 0.32fF
C10228 a_5691_36727# a_4811_34855# 0.35fF
C10229 vcm_commonmode a_37446_72234# 0.69fF
C10230 a_37446_61190# a_38450_61190# 0.97fF
C10231 a_6467_55527# a_7107_58487# 0.38fF
C10232 a_3355_25071# VDD 0.83fF
C10233 a_28318_24918# a_28410_24552# 0.32fF
C10234 a_13107_34789# VDD 0.93fF
C10235 a_29414_7484# VDD 1.60fF
C10236 a_13005_43983# a_12663_40871# 0.58fF
C10237 a_43470_68218# a_43470_67214# 1.00fF
C10238 a_39299_48783# a_44474_63198# 0.42fF
C10239 a_16955_52047# a_4758_45369# 0.43fF
C10240 a_2216_28309# a_3325_29967# 0.40fF
C10241 a_25971_52263# a_30418_69222# 0.38fF
C10242 vcm_commonmode a_36442_68218# 0.87fF
C10243 a_23390_64202# VDD 0.51fF
C10244 a_25306_62194# a_25398_62194# 0.32fF
C10245 a_31422_56170# ctopp 3.40fF
C10246 a_7155_55509# a_9424_60949# 0.67fF
C10247 ctopn a_25398_18528# 3.59fF
C10248 vcm_commonmode a_30326_64202# 0.31fF
C10249 a_28410_69222# a_28410_68218# 1.00fF
C10250 a_21187_29415# VDD 8.19fF
C10251 a_18370_8488# a_18370_7484# 1.00fF
C10252 a_40458_8488# a_41462_8488# 0.97fF
C10253 a_38358_55166# a_38450_55166# 0.32fF
C10254 vcm_commonmode a_16746_10494# 5.36fF
C10255 a_1923_59583# VDD 6.23fF
C10256 a_30326_57174# a_30418_57174# 0.32fF
C10257 a_33338_15882# a_33430_15516# 0.32fF
C10258 a_12381_43957# VDD 9.27fF
C10259 vcm_commonmode a_10975_66407# 6.22fF
C10260 a_41462_70226# a_42466_70226# 0.97fF
C10261 a_39673_28111# a_12877_16911# 0.41fF
C10262 a_9485_62613# VDD 0.58fF
C10263 a_12447_29199# a_38210_30199# 0.43fF
C10264 a_18307_27791# VDD 0.34fF
C10265 a_30418_61190# ctopp 3.59fF
C10266 ctopn a_34434_10496# 3.59fF
C10267 a_32426_69222# VDD 0.51fF
C10268 a_17863_36595# VDD 1.61fF
C10269 vcm_commonmode a_18278_19898# 0.31fF
C10270 a_21371_52263# a_12869_2741# 6.91fF
C10271 a_29760_55394# a_29414_55166# 0.46fF
C10272 a_2021_17973# a_13716_43047# 1.34fF
C10273 a_2191_68565# a_2099_64757# 0.76fF
C10274 a_22386_16520# a_23390_16520# 0.97fF
C10275 vcm_commonmode a_36442_56170# 0.87fF
C10276 a_31330_71230# a_31422_71230# 0.32fF
C10277 vcm_commonmode a_39362_69222# 0.31fF
C10278 a_7519_59575# a_4298_58951# 0.59fF
C10279 a_39454_60186# a_39454_59182# 1.00fF
C10280 a_39454_22544# VDD 0.51fF
C10281 vcm_commonmode a_19374_8488# 0.86fF
C10282 a_9503_26151# a_20378_20536# 0.38fF
C10283 a_30418_65206# VDD 0.51fF
C10284 a_29927_29199# a_35815_31751# 0.53fF
C10285 a_49494_24552# m3_49396_24414# 2.81fF
C10286 a_28410_63198# a_28410_62194# 1.00fF
C10287 a_43378_11866# a_43470_11500# 0.32fF
C10288 a_7987_64213# a_6515_62037# 0.38fF
C10289 a_48490_15516# a_48490_14512# 1.00fF
C10290 a_51936_39932# VDD 0.36fF
C10291 vcm_commonmode a_46390_22910# 0.31fF
C10292 a_34434_70226# ctopp 3.58fF
C10293 vcm_commonmode m3_16264_20398# 3.21fF
C10294 a_32887_42405# VDD 0.93fF
C10295 vcm_commonmode a_37354_65206# 0.31fF
C10296 a_2292_17179# a_7571_16917# 0.35fF
C10297 a_8583_33551# a_1761_49007# 0.44fF
C10298 a_33430_9492# a_33430_8488# 1.00fF
C10299 a_19282_24918# VDD 0.36fF
C10300 a_47394_24918# a_47486_24552# 0.32fF
C10301 a_3339_32463# a_5915_30287# 0.44fF
C10302 a_11521_66567# a_11521_58951# 0.47fF
C10303 ctopn a_29414_15516# 3.59fF
C10304 a_28410_67214# a_29414_67214# 0.97fF
C10305 vcm_commonmode a_35438_61190# 0.87fF
C10306 a_7000_43541# a_3339_32463# 0.92fF
C10307 a_35438_14512# VDD 0.51fF
C10308 a_10699_69679# a_10865_69679# 0.72fF
C10309 a_9503_26151# a_20378_12504# 0.38fF
C10310 a_9872_20175# VDD 0.31fF
C10311 a_30326_55166# VDD 0.35fF
C10312 a_1643_63125# VDD 0.36fF
C10313 a_44382_62194# a_44474_62194# 0.32fF
C10314 a_20747_27765# VDD 1.08fF
C10315 vcm_commonmode a_42374_14878# 0.31fF
C10316 ctopn a_39454_11500# 3.59fF
C10317 a_18127_35797# a_1761_27791# 0.64fF
C10318 vcm_commonmode a_21290_20902# 0.31fF
C10319 a_31280_40517# VDD 1.90fF
C10320 a_47486_69222# a_47486_68218# 1.00fF
C10321 a_9989_46831# VDD 1.85fF
C10322 a_43362_28879# a_12901_66665# 0.40fF
C10323 vcm_commonmode a_39454_70226# 0.87fF
C10324 a_2163_59585# VDD 0.47fF
C10325 a_37446_8488# a_37446_7484# 1.00fF
C10326 a_40458_23548# VDD 0.52fF
C10327 a_23390_58178# ctopp 3.59fF
C10328 a_43270_27791# a_45478_21540# 0.38fF
C10329 a_37446_66210# VDD 0.51fF
C10330 VDD config_1_in[15] 1.16fF
C10331 vcm_commonmode a_20378_16520# 0.87fF
C10332 a_17507_52047# a_17682_50095# 0.51fF
C10333 a_37551_42333# a_19967_41781# 0.38fF
C10334 a_49402_57174# a_49494_57174# 0.32fF
C10335 vcm_commonmode a_47394_23914# 0.31fF
C10336 a_1761_49007# a_34222_43439# 0.35fF
C10337 a_20743_43493# VDD 0.82fF
C10338 vcm_commonmode a_44382_66210# 0.31fF
C10339 a_30418_58178# a_31422_58178# 0.97fF
C10340 a_49494_19532# VDD 1.13fF
C10341 a_2686_70223# a_2843_71829# 0.50fF
C10342 a_9503_26151# a_20378_17524# 0.38fF
C10343 a_25398_9492# a_26402_9492# 0.97fF
C10344 a_28589_27247# VDD 0.41fF
C10345 vcm_commonmode a_21290_12870# 0.31fF
C10346 a_26402_13508# a_26402_12504# 1.00fF
C10347 a_35647_35877# VDD 0.96fF
C10348 a_40458_67214# ctopp 3.59fF
C10349 a_13390_29575# a_9529_28335# 0.38fF
C10350 a_12357_37999# a_13067_38517# 1.02fF
C10351 a_41462_16520# a_42466_16520# 0.97fF
C10352 a_4811_34855# a_30788_28487# 1.03fF
C10353 a_26523_28111# VDD 8.79fF
C10354 a_11067_13095# a_7078_36103# 0.30fF
C10355 a_2099_59861# a_4674_40277# 0.67fF
C10356 a_8933_22583# a_10275_21495# 0.34fF
C10357 a_47486_63198# a_47486_62194# 1.00fF
C10358 a_3247_10389# a_3413_10389# 0.42fF
C10359 a_12801_38517# a_23415_41263# 0.31fF
C10360 vcm_commonmode a_28410_58178# 0.87fF
C10361 a_41872_29423# a_12901_58799# 0.40fF
C10362 vcm_commonmode a_16362_21540# 4.47fF
C10363 a_1689_10396# a_3327_9308# 0.42fF
C10364 a_19720_55394# a_19374_65206# 0.38fF
C10365 a_12901_66959# a_16362_68218# 1.15fF
C10366 a_36821_50095# VDD 0.63fF
C10367 a_4339_64521# a_7050_53333# 0.31fF
C10368 a_2787_30503# VDD 13.39fF
C10369 vcm_commonmode a_21290_17890# 0.31fF
C10370 a_18053_28879# a_20747_27765# 0.34fF
C10371 a_2021_17973# a_2339_38129# 0.50fF
C10372 a_2451_72373# VDD 5.64fF
C10373 a_12983_63151# a_16746_66212# 2.28fF
C10374 a_16955_52047# a_12981_59343# 0.40fF
C10375 a_47486_67214# a_48490_67214# 0.97fF
C10376 vcm_commonmode a_10055_58791# 6.29fF
C10377 a_17488_48731# a_4674_40277# 0.39fF
C10378 a_4443_46607# a_10407_47607# 0.37fF
C10379 vcm_commonmode a_45478_67214# 0.87fF
C10380 a_34251_52263# a_35438_68218# 0.38fF
C10381 a_10680_54171# VDD 0.58fF
C10382 a_1586_69367# a_1923_73087# 0.35fF
C10383 a_2411_19605# a_1586_9991# 0.33fF
C10384 a_41462_63198# VDD 0.57fF
C10385 a_10515_22671# a_16362_57174# 1.15fF
C10386 a_29322_13874# a_29414_13508# 0.32fF
C10387 a_18811_36965# VDD 0.86fF
C10388 a_20881_28111# a_15681_27497# 0.35fF
C10389 a_3339_43023# a_12970_34191# 0.32fF
C10390 a_1761_22895# a_13716_43047# 1.59fF
C10391 a_14258_44527# a_1803_20719# 0.85fF
C10392 a_43267_31055# a_12355_15055# 0.40fF
C10393 vcm_commonmode a_48398_63198# 0.31fF
C10394 a_34342_68218# a_34434_68218# 0.32fF
C10395 a_43362_28879# a_43269_29967# 0.43fF
C10396 a_21187_29415# a_34482_29941# 0.56fF
C10397 a_7387_48469# VDD 0.46fF
C10398 a_16955_52047# a_20378_70226# 0.38fF
C10399 a_34780_56398# a_12516_7093# 0.40fF
C10400 a_4891_47388# a_2595_47653# 0.31fF
C10401 a_1591_19631# a_1757_19631# 0.69fF
C10402 a_35438_59182# VDD 0.51fF
C10403 a_33430_7484# a_34434_7484# 0.97fF
C10404 a_11308_22057# VDD 0.44fF
C10405 vcm_commonmode a_42466_9492# 0.87fF
C10406 a_12981_62313# a_16362_62194# 1.15fF
C10407 a_39454_64202# ctopp 3.59fF
C10408 ctopn a_44474_13508# 3.59fF
C10409 a_16955_52047# a_30525_49551# 0.39fF
C10410 a_43378_72234# VDD 0.61fF
C10411 vcm_commonmode a_42374_59182# 0.31fF
C10412 a_25787_28327# a_33430_60186# 0.38fF
C10413 vcm_commonmode a_22386_22544# 0.87fF
C10414 a_17599_52263# a_22386_66210# 0.38fF
C10415 a_17366_69222# a_18370_69222# 0.97fF
C10416 a_35601_27497# a_35438_10496# 0.38fF
C10417 a_26397_51183# a_27869_50095# 1.07fF
C10418 a_16362_72234# a_17366_72234# 0.97fF
C10419 a_2419_48783# a_8295_47388# 0.44fF
C10420 a_26748_7638# a_12727_15529# 0.41fF
C10421 a_31768_7638# a_31422_15516# 0.38fF
C10422 a_9135_27239# a_12727_13353# 0.41fF
C10423 a_9215_61127# VDD 0.54fF
C10424 a_3339_43023# a_11067_46823# 0.32fF
C10425 a_44474_9492# a_45478_9492# 0.97fF
C10426 a_11619_56615# a_9989_46831# 0.59fF
C10427 a_23736_7638# a_12895_13967# 0.41fF
C10428 a_3339_32463# a_5915_35943# 0.48fF
C10429 a_27406_64202# a_28410_64202# 0.97fF
C10430 a_45478_13508# a_45478_12504# 1.00fF
C10431 vcm_commonmode a_22294_18894# 0.31fF
C10432 a_11067_63143# a_12024_30199# 0.64fF
C10433 a_12355_65103# a_3339_43023# 0.66fF
C10434 a_17507_52047# a_21382_62194# 0.38fF
C10435 a_34251_52263# a_35438_56170# 0.38fF
C10436 a_18703_29199# a_24959_30503# 7.52fF
C10437 a_4215_51157# a_2872_44111# 1.08fF
C10438 a_47486_21540# VDD 0.51fF
C10439 a_24394_22544# a_25398_22544# 0.97fF
C10440 a_39727_27765# VDD 0.64fF
C10441 a_10239_57167# VDD 0.51fF
C10442 vcm_commonmode a_18370_14512# 0.88fF
C10443 a_7387_69929# VDD 0.52fF
C10444 a_7749_37903# VDD 0.70fF
C10445 a_48490_69222# ctopp 3.43fF
C10446 a_1761_46287# a_1761_44111# 1.77fF
C10447 a_24394_10496# VDD 0.51fF
C10448 vcm_commonmode a_44474_64202# 0.87fF
C10449 a_1586_40455# a_2606_41079# 0.50fF
C10450 a_25971_52263# a_12907_56399# 2.22fF
C10451 a_39454_60186# VDD 0.51fF
C10452 a_16746_23546# VDD 33.42fF
C10453 vcm_commonmode a_31330_10862# 0.31fF
C10454 a_30440_31573# VDD 0.53fF
C10455 a_46482_65206# ctopp 3.59fF
C10456 a_5254_67503# a_8999_61493# 1.30fF
C10457 vcm_commonmode a_46390_60186# 0.31fF
C10458 a_35438_67214# a_35438_66210# 1.00fF
C10459 vcm_commonmode a_23390_23548# 0.87fF
C10460 a_21382_7484# m3_21284_7346# 2.80fF
C10461 a_15607_46805# a_12447_29199# 2.40fF
C10462 a_26267_43983# VDD 0.35fF
C10463 vcm_commonmode a_20378_66210# 0.87fF
C10464 a_12473_37429# a_13576_37149# 0.97fF
C10465 a_19502_51157# a_19946_51157# 0.72fF
C10466 a_36629_27791# VDD 6.49fF
C10467 a_9135_27239# a_10515_23975# 0.41fF
C10468 a_31422_65206# a_31422_64202# 1.00fF
C10469 a_48398_13874# a_48490_13508# 0.32fF
C10470 vcm_commonmode a_32426_19532# 0.87fF
C10471 a_16362_67214# ctopp 1.35fF
C10472 vcm_commonmode a_18278_62194# 0.31fF
C10473 a_40050_48463# a_12257_56623# 0.40fF
C10474 a_19374_15516# VDD 0.51fF
C10475 a_25398_23548# a_25398_22544# 1.00fF
C10476 a_41967_31375# a_12985_16367# 0.41fF
C10477 a_18127_35797# a_13669_38517# 0.54fF
C10478 a_1768_16367# a_1591_56623# 0.52fF
C10479 a_7803_55509# a_8491_57487# 1.18fF
C10480 a_1895_30138# VDD 0.53fF
C10481 vcm_commonmode a_26310_15882# 0.31fF
C10482 a_19374_63198# ctopp 3.64fF
C10483 a_16955_52047# a_32227_48169# 0.75fF
C10484 a_34342_56170# a_34434_56170# 0.32fF
C10485 a_17366_71230# VDD 0.64fF
C10486 a_39222_48169# a_10515_22671# 0.40fF
C10487 a_19374_66210# a_19374_65206# 1.00fF
C10488 a_1768_13103# config_1_in[5] 0.43fF
C10489 a_20378_14512# a_21382_14512# 0.97fF
C10490 a_11067_67279# a_28756_7638# 0.41fF
C10491 a_22386_72234# m3_22288_72146# 2.80fF
C10492 a_29414_11500# VDD 0.51fF
C10493 a_15931_39859# VDD 0.71fF
C10494 a_36442_69222# a_37446_69222# 0.97fF
C10495 a_12341_3311# a_22386_10496# 0.38fF
C10496 vcm_commonmode a_24302_71230# 0.31fF
C10497 a_26402_72234# a_27406_72234# 0.97fF
C10498 a_31422_61190# a_31422_60186# 1.00fF
C10499 a_17274_8854# a_17366_8488# 0.32fF
C10500 a_33430_24552# VDD 0.60fF
C10501 vcm_commonmode a_36350_11866# 0.31fF
C10502 a_46482_64202# a_47486_64202# 0.97fF
C10503 a_2099_59861# a_14298_32143# 0.63fF
C10504 a_12516_7093# a_11067_47695# 9.72fF
C10505 vcm_commonmode a_40366_24918# 0.31fF
C10506 a_23395_52047# a_8583_33551# 0.31fF
C10507 a_4811_34855# a_23736_7638# 0.49fF
C10508 a_13357_32143# a_14646_29423# 0.56fF
C10509 a_34482_29941# a_26523_28111# 0.45fF
C10510 a_18278_70226# a_18370_70226# 0.32fF
C10511 a_4215_51157# a_9668_51451# 0.59fF
C10512 a_43470_55166# VDD 0.60fF
C10513 a_43470_22544# a_44474_22544# 0.97fF
C10514 a_17366_62194# a_17366_61190# 1.00fF
C10515 a_35438_57174# VDD 0.51fF
C10516 VDD result_out[1] 0.73fF
C10517 a_34434_65206# a_35438_65206# 0.97fF
C10518 vcm_commonmode a_35438_20536# 0.87fF
C10519 vcm_commonmode a_24394_63198# 0.92fF
C10520 a_30418_17524# a_30418_16520# 1.00fF
C10521 vcm_commonmode a_42374_57174# 0.31fF
C10522 a_2606_41079# a_1761_49007# 1.72fF
C10523 a_21169_49007# VDD 0.33fF
C10524 a_4891_47388# a_23487_50095# 0.37fF
C10525 a_17366_20536# a_17366_19532# 1.00fF
C10526 a_25398_23548# a_26402_23548# 0.97fF
C10527 a_21371_50959# a_29147_50069# 0.43fF
C10528 a_9179_22351# a_8935_27791# 1.17fF
C10529 a_1761_41935# a_18127_35797# 3.10fF
C10530 a_25398_72234# VDD 1.59fF
C10531 a_22386_66210# a_23390_66210# 0.97fF
C10532 a_28756_55394# a_12727_58255# 0.40fF
C10533 vcm_commonmode a_18370_59182# 0.88fF
C10534 a_4351_67279# a_11067_67279# 4.10fF
C10535 ctopn a_32772_7638# 2.66fF
C10536 a_12473_37429# a_12381_35836# 0.42fF
C10537 a_2686_70223# a_4119_70741# 0.46fF
C10538 vcm_commonmode a_30418_72234# 0.69fF
C10539 a_33864_28111# a_12985_16367# 0.41fF
C10540 a_49494_62194# VDD 1.10fF
C10541 a_33338_61190# a_33430_61190# 0.32fF
C10542 a_1761_25615# VDD 0.38fF
C10543 a_12659_54965# VDD 1.44fF
C10544 vcm_commonmode a_35438_12504# 0.87fF
C10545 a_17366_60186# ctopp 3.43fF
C10546 ctopn a_36442_9492# 3.58fF
C10547 a_20378_68218# VDD 0.51fF
C10548 a_1768_13103# a_1591_54447# 0.64fF
C10549 a_12381_43957# a_12663_40871# 1.77fF
C10550 a_20286_7850# VDD 0.62fF
C10551 a_39222_48169# a_40458_63198# 0.42fF
C10552 a_7155_55509# a_7803_55509# 0.79fF
C10553 ctopn a_16746_22542# 1.67fF
C10554 a_2292_43291# a_4563_32900# 0.78fF
C10555 a_21371_52263# a_26402_69222# 0.38fF
C10556 vcm_commonmode a_27314_68218# 0.31fF
C10557 a_22386_71230# a_22386_70226# 1.00fF
C10558 a_34434_19532# a_35438_19532# 0.97fF
C10559 a_8583_33551# a_34222_43439# 2.21fF
C10560 a_39673_28111# a_40458_19532# 0.38fF
C10561 a_44474_23548# a_44474_22544# 1.00fF
C10562 a_29760_7638# a_12985_19087# 0.41fF
C10563 a_10975_65327# a_11141_65327# 0.72fF
C10564 a_2840_66103# a_4339_64521# 3.18fF
C10565 a_38450_66210# a_38450_65206# 1.00fF
C10566 a_3327_9308# a_9227_12015# 0.55fF
C10567 a_39454_14512# a_40458_14512# 0.97fF
C10568 vcm_commonmode a_30418_21540# 0.87fF
C10569 ctopn a_16362_18528# 1.35fF
C10570 vcm_commonmode a_48490_58178# 0.87fF
C10571 a_41427_52263# a_41462_72234# 0.34fF
C10572 a_18370_20536# a_19374_20536# 0.97fF
C10573 a_36350_8854# a_36442_8488# 0.32fF
C10574 a_49494_24552# VDD 1.18fF
C10575 a_22291_29415# a_4811_34855# 0.40fF
C10576 a_35815_31751# VDD 3.07fF
C10577 vcm_commonmode a_35438_17524# 0.87fF
C10578 vcm_commonmode a_22386_60186# 0.87fF
C10579 a_7939_30503# a_11155_30663# 0.41fF
C10580 a_34434_13508# VDD 0.51fF
C10581 a_21095_47919# a_21261_47919# 0.39fF
C10582 a_35217_44509# VDD 0.78fF
C10583 a_37354_70226# a_37446_70226# 0.32fF
C10584 a_6743_19881# VDD 1.14fF
C10585 a_6559_59663# a_8295_47388# 0.61fF
C10586 a_1586_51335# a_9707_51325# 0.43fF
C10587 a_43269_29967# a_12727_15529# 0.41fF
C10588 a_42709_29199# a_12985_16367# 0.40fF
C10589 a_36442_62194# a_36442_61190# 1.00fF
C10590 a_27406_10496# a_27406_9492# 1.00fF
C10591 a_20378_56170# VDD 0.52fF
C10592 vcm_commonmode a_41370_13874# 0.31fF
C10593 a_8199_58229# a_7479_54439# 1.34fF
C10594 a_4351_67279# a_12907_27023# 0.52fF
C10595 a_12641_36596# VDD 2.45fF
C10596 a_21371_50959# a_25398_55166# 0.47fF
C10597 a_18278_16886# a_18370_16520# 0.32fF
C10598 a_49494_17524# a_49494_16520# 1.00fF
C10599 a_18611_52047# a_12899_3855# 4.59fF
C10600 vcm_commonmode a_27314_56170# 0.31fF
C10601 ctopn a_17366_23548# 0.37fF
C10602 a_9275_15253# VDD 0.86fF
C10603 a_25015_48437# VDD 1.02fF
C10604 a_36442_20536# a_36442_19532# 1.00fF
C10605 a_44474_23548# a_45478_23548# 0.97fF
C10606 a_12257_56623# ctopp 2.99fF
C10607 a_41462_66210# a_42466_66210# 0.97fF
C10608 ctopn a_26402_19532# 3.59fF
C10609 a_8753_31055# a_10531_31055# 0.52fF
C10610 a_4674_40277# a_2787_32679# 1.33fF
C10611 a_2007_10901# VDD 0.40fF
C10612 a_40050_48463# a_10975_66407# 0.40fF
C10613 ctopn a_37919_28111# 2.62fF
C10614 a_24849_51183# VDD 0.65fF
C10615 a_32951_27247# a_12727_13353# 0.41fF
C10616 a_9503_26151# a_12985_16367# 0.41fF
C10617 a_19374_61190# VDD 0.51fF
C10618 a_7571_29199# a_9179_22351# 0.36fF
C10619 a_4298_58951# a_7749_55535# 0.85fF
C10620 a_11803_55311# a_12725_44527# 1.65fF
C10621 a_18370_12504# a_19374_12504# 0.97fF
C10622 vcm_commonmode a_36442_18528# 0.87fF
C10623 a_13390_29575# a_14273_27791# 0.53fF
C10624 a_24302_67214# a_24394_67214# 0.32fF
C10625 vcm_commonmode a_26310_61190# 0.31fF
C10626 vcm_commonmode a_16362_24552# 1.87fF
C10627 a_41462_71230# a_41462_70226# 1.00fF
C10628 a_3143_66972# a_4351_67279# 0.49fF
C10629 a_1586_51335# a_5612_52520# 0.81fF
C10630 a_9424_60949# a_9526_61751# 0.50fF
C10631 a_7169_56311# VDD 0.32fF
C10632 a_27406_62194# ctopp 3.59fF
C10633 a_1761_40847# a_1761_39215# 1.91fF
C10634 a_23390_70226# VDD 0.51fF
C10635 a_36579_38007# VDD 0.64fF
C10636 a_40458_58178# VDD 0.51fF
C10637 vcm_commonmode a_27406_55166# 0.84fF
C10638 vcm_commonmode a_18370_57174# 0.88fF
C10639 a_36551_49007# VDD 0.38fF
C10640 a_39222_48169# a_12901_66665# 0.40fF
C10641 vcm_commonmode a_30326_70226# 0.31fF
C10642 a_37446_20536# a_38450_20536# 0.97fF
C10643 vcm_commonmode a_45478_10496# 0.87fF
C10644 a_26402_63198# a_27406_63198# 0.97fF
C10645 a_16270_72234# VDD 0.74fF
C10646 a_10975_66407# a_12355_65103# 24.99fF
C10647 a_33430_71230# ctopp 3.40fF
C10648 ctopn a_29414_20536# 3.59fF
C10649 a_33694_30761# a_32970_31145# 0.32fF
C10650 a_15548_30761# a_23747_31055# 0.31fF
C10651 a_20881_28111# a_23626_31573# 0.43fF
C10652 a_10055_58791# a_16746_12502# 2.28fF
C10653 a_24740_7638# a_24394_10496# 0.38fF
C10654 a_14287_51175# a_14646_29423# 2.41fF
C10655 a_26310_58178# a_26402_58178# 0.32fF
C10656 a_42709_29199# a_48490_16520# 0.38fF
C10657 a_43175_28335# a_12727_13353# 0.41fF
C10658 a_46482_10496# a_46482_9492# 1.00fF
C10659 a_21290_9858# a_21382_9492# 0.32fF
C10660 a_32951_27247# a_10515_23975# 0.40fF
C10661 a_14675_35831# VDD 0.62fF
C10662 a_2539_42106# a_2411_26133# 0.68fF
C10663 a_41462_8488# VDD 0.58fF
C10664 vcm_commonmode a_32426_62194# 0.87fF
C10665 a_37354_16886# a_37446_16520# 0.32fF
C10666 a_5039_42167# a_17488_48731# 1.01fF
C10667 a_12047_57685# VDD 0.45fF
C10668 a_20378_59182# a_21382_59182# 0.97fF
C10669 a_11763_21237# VDD 0.51fF
C10670 vcm_commonmode a_48398_8854# 0.31fF
C10671 a_39673_28111# a_12895_13967# 0.41fF
C10672 a_6831_63303# a_6382_61127# 0.56fF
C10673 a_13390_29575# VDD 2.31fF
C10674 vcm_commonmode a_40458_15516# 0.87fF
C10675 ctopn a_29414_12504# 3.59fF
C10676 vcm_commonmode a_19282_58178# 0.31fF
C10677 a_36717_47375# a_12901_58799# 0.40fF
C10678 a_30875_39095# VDD 0.63fF
C10679 a_12935_31287# a_6459_30511# 0.33fF
C10680 a_35033_42044# VDD 0.92fF
C10681 a_18370_17524# a_19374_17524# 0.97fF
C10682 a_1761_31055# a_32327_35839# 1.53fF
C10683 a_10055_58791# a_12899_11471# 0.70fF
C10684 a_23271_50943# VDD 0.52fF
C10685 vcm_commonmode a_38450_71230# 0.86fF
C10686 a_32334_72234# a_32426_72234# 0.32fF
C10687 a_1923_54591# a_1683_52271# 0.57fF
C10688 a_35438_21540# a_35438_20536# 1.00fF
C10689 a_3295_62083# a_4674_57685# 0.36fF
C10690 a_22386_24552# a_22386_23548# 1.00fF
C10691 a_29414_67214# VDD 0.51fF
C10692 a_37446_12504# a_38450_12504# 0.97fF
C10693 a_9529_28335# a_12985_25615# 1.02fF
C10694 a_12357_37999# a_12473_41781# 2.09fF
C10695 a_43378_67214# a_43470_67214# 0.32fF
C10696 ctopn a_24394_21540# 3.59fF
C10697 a_3983_12879# VDD 0.42fF
C10698 vcm_commonmode a_36350_67214# 0.31fF
C10699 a_31768_55394# a_31422_68218# 0.38fF
C10700 a_7755_74581# a_8575_74853# 0.35fF
C10701 a_43269_29967# a_47486_16520# 0.38fF
C10702 a_7295_44647# a_17651_30485# 0.37fF
C10703 a_8453_51727# a_9668_51451# 0.69fF
C10704 vcm_commonmode a_17366_13508# 1.82fF
C10705 a_43175_28335# a_10515_23975# 0.41fF
C10706 a_2216_28309# VDD 5.88fF
C10707 a_36442_68218# ctopp 3.59fF
C10708 ctopn a_29414_17524# 3.59fF
C10709 a_26402_9492# VDD 0.51fF
C10710 a_36708_39655# VDD 1.80fF
C10711 a_39389_52271# a_12355_15055# 0.40fF
C10712 a_22015_28111# a_20635_29415# 0.45fF
C10713 a_19807_28111# a_16863_29415# 0.82fF
C10714 a_42466_16520# VDD 0.51fF
C10715 a_43267_31055# a_46482_71230# 0.38fF
C10716 a_12947_71576# a_12901_66665# 23.41fF
C10717 a_23395_52047# a_12516_7093# 0.40fF
C10718 a_29322_7850# a_29414_7484# 0.32fF
C10719 vcm_commonmode a_33338_9858# 0.31fF
C10720 m3_41364_72146# VDD 0.42fF
C10721 a_34482_29941# a_35815_31751# 0.61fF
C10722 a_3339_32463# a_7939_30503# 1.01fF
C10723 a_41462_24552# m3_41364_24414# 2.81fF
C10724 a_45478_63198# a_46482_63198# 0.97fF
C10725 a_33641_29967# VDD 3.28fF
C10726 vcm_commonmode a_49402_16886# 0.30fF
C10727 a_3949_41935# a_4314_40821# 1.58fF
C10728 a_36350_72234# VDD 0.62fF
C10729 a_29760_55394# a_29414_60186# 0.38fF
C10730 a_22595_43177# VDD 0.62fF
C10731 a_14287_51175# a_18370_66210# 0.38fF
C10732 a_40050_48463# a_45478_67214# 0.38fF
C10733 a_19374_18528# a_19374_17524# 1.00fF
C10734 a_1761_37039# a_13005_35823# 2.44fF
C10735 a_7841_12167# a_9367_29397# 0.96fF
C10736 a_43270_27791# a_12727_13353# 0.41fF
C10737 a_32426_21540# a_33430_21540# 0.97fF
C10738 a_3938_61493# VDD 0.60fF
C10739 a_40366_9858# a_40458_9492# 0.32fF
C10740 a_10472_26159# VDD 2.22fF
C10741 a_23298_64202# a_23390_64202# 0.32fF
C10742 a_10975_66407# ctopp 3.23fF
C10743 a_34434_7484# VDD 1.37fF
C10744 a_31768_55394# a_31422_56170# 0.38fF
C10745 a_1929_10651# VDD 4.32fF
C10746 a_33802_47375# VDD 0.32fF
C10747 vcm_commonmode a_41462_68218# 0.87fF
C10748 a_39454_59182# a_40458_59182# 0.97fF
C10749 a_6467_55527# a_13925_51727# 0.56fF
C10750 a_1770_14441# a_1689_10396# 0.33fF
C10751 a_8491_27023# a_18370_19532# 0.38fF
C10752 a_25744_7638# a_25398_19532# 0.38fF
C10753 a_20286_22910# a_20378_22544# 0.32fF
C10754 a_28410_64202# VDD 0.51fF
C10755 a_37919_28111# a_36797_27497# 0.30fF
C10756 a_36442_56170# ctopp 3.40fF
C10757 a_6598_69653# VDD 0.53fF
C10758 a_6095_44807# a_6515_62037# 0.75fF
C10759 a_20378_14512# a_20378_13508# 1.00fF
C10760 ctopn a_30418_18528# 3.59fF
C10761 a_15683_40767# VDD 1.05fF
C10762 vcm_commonmode a_35346_64202# 0.31fF
C10763 a_37446_17524# a_38450_17524# 0.97fF
C10764 a_5915_30287# a_4903_31849# 0.34fF
C10765 a_13005_35823# a_1761_32143# 2.80fF
C10766 a_24394_60186# a_25398_60186# 0.97fF
C10767 a_8105_21263# VDD 0.54fF
C10768 a_31768_7638# a_31422_20536# 0.38fF
C10769 a_41462_24552# a_41462_23548# 1.00fF
C10770 a_8307_66415# VDD 0.33fF
C10771 a_26402_12504# a_26402_11500# 1.00fF
C10772 a_13183_52047# a_22989_48437# 0.34fF
C10773 a_12641_43124# a_12641_42036# 3.09fF
C10774 a_9707_73807# VDD 0.38fF
C10775 a_6559_22671# a_4674_40277# 0.31fF
C10776 a_11803_55311# a_12727_67753# 1.07fF
C10777 a_19374_18528# a_20378_18528# 0.97fF
C10778 a_16746_19530# VDD 33.20fF
C10779 a_6224_73095# a_6327_72917# 0.64fF
C10780 a_1770_14441# a_2004_42453# 0.39fF
C10781 vcm_commonmode inn_analog 0.59fF
C10782 a_35438_61190# ctopp 3.59fF
C10783 ctopn a_39454_10496# 3.59fF
C10784 a_43270_27791# a_10515_23975# 0.41fF
C10785 a_13867_39958# a_13669_39605# 0.30fF
C10786 a_37446_69222# VDD 0.51fF
C10787 a_1923_59583# a_9319_62613# 0.34fF
C10788 a_4812_13879# a_5345_10927# 0.60fF
C10789 vcm_commonmode a_23298_19898# 0.31fF
C10790 a_38557_32143# a_12257_56623# 0.40fF
C10791 vcm_commonmode a_41462_56170# 0.87fF
C10792 a_1761_34319# a_35602_34191# 0.31fF
C10793 vcm_commonmode a_44382_69222# 0.31fF
C10794 a_31768_7638# a_31422_12504# 0.38fF
C10795 a_3714_58345# VDD 2.41fF
C10796 a_48398_7850# a_48490_7484# 0.32fF
C10797 a_44474_22544# VDD 0.51fF
C10798 vcm_commonmode a_24394_8488# 0.86fF
C10799 a_35438_65206# VDD 0.51fF
C10800 a_9319_62613# a_9485_62613# 0.47fF
C10801 a_26063_30511# VDD 0.36fF
C10802 vcm_commonmode a_12877_14441# 6.31fF
C10803 a_10515_63143# a_3339_43023# 1.14fF
C10804 a_9063_71553# VDD 0.43fF
C10805 a_25787_28327# a_10515_22671# 0.40fF
C10806 a_39454_70226# ctopp 3.58fF
C10807 vcm_commonmode a_42374_65206# 0.31fF
C10808 a_32334_69222# a_32426_69222# 0.32fF
C10809 a_1950_59887# a_10975_65327# 0.56fF
C10810 a_38450_18528# a_38450_17524# 1.00fF
C10811 a_19720_55394# a_28756_55394# 0.43fF
C10812 a_18611_52047# a_18151_52263# 0.40fF
C10813 a_8491_57487# a_11303_53511# 0.61fF
C10814 a_12447_29199# a_28841_29575# 1.72fF
C10815 a_12641_37684# a_13669_35253# 0.96fF
C10816 a_24302_24918# VDD 0.36fF
C10817 a_42374_64202# a_42466_64202# 0.32fF
C10818 ctopn a_34434_15516# 3.59fF
C10819 vcm_commonmode a_40458_61190# 0.87fF
C10820 a_9307_30663# a_2787_30503# 0.34fF
C10821 a_4811_34855# a_27797_29423# 0.67fF
C10822 a_13643_28327# a_18979_30287# 2.13fF
C10823 a_40458_14512# VDD 0.51fF
C10824 a_4259_45199# VDD 0.39fF
C10825 a_19374_20536# VDD 0.51fF
C10826 a_34342_55166# VDD 0.36fF
C10827 a_31768_7638# a_31422_17524# 0.38fF
C10828 a_39362_22910# a_39454_22544# 0.32fF
C10829 a_5274_62313# VDD 0.54fF
C10830 a_6372_38279# a_5915_30287# 1.40fF
C10831 a_12907_27023# a_15799_29941# 0.58fF
C10832 a_13669_39605# a_13669_38517# 0.31fF
C10833 a_28410_10496# a_29414_10496# 0.97fF
C10834 vcm_commonmode a_47394_14878# 0.31fF
C10835 ctopn a_44474_11500# 3.59fF
C10836 a_1761_40847# a_1799_29556# 0.31fF
C10837 a_30326_65206# a_30418_65206# 0.32fF
C10838 a_39454_14512# a_39454_13508# 1.00fF
C10839 vcm_commonmode a_26310_20902# 0.31fF
C10840 a_7803_55509# a_7479_54439# 0.58fF
C10841 a_2235_30503# a_24768_27247# 0.70fF
C10842 a_3339_43023# a_3607_34639# 0.35fF
C10843 a_52778_39198# VDD 1.01fF
C10844 a_11067_67279# a_7939_30503# 0.42fF
C10845 vcm_commonmode a_44474_70226# 0.87fF
C10846 a_7519_59575# VDD 1.14fF
C10847 a_43470_60186# a_44474_60186# 0.97fF
C10848 a_8295_47388# a_7050_53333# 0.32fF
C10849 a_45478_23548# VDD 0.52fF
C10850 a_28410_58178# ctopp 3.59fF
C10851 a_21290_23914# a_21382_23548# 0.32fF
C10852 a_9503_26151# a_20378_21540# 0.38fF
C10853 a_49494_24552# a_49494_23548# 1.00fF
C10854 a_42466_66210# VDD 0.51fF
C10855 VDD config_1_in[0] 0.90fF
C10856 a_45478_12504# a_45478_11500# 1.00fF
C10857 a_10531_31055# VDD 2.33fF
C10858 vcm_commonmode a_25398_16520# 0.87fF
C10859 a_18370_72234# VDD 1.42fF
C10860 a_18278_66210# a_18370_66210# 0.32fF
C10861 a_17507_52047# a_12727_58255# 0.40fF
C10862 a_19374_12504# VDD 0.51fF
C10863 a_1761_49007# a_13716_43047# 1.18fF
C10864 a_31648_43781# VDD 1.74fF
C10865 a_5682_69367# a_5024_67885# 0.38fF
C10866 vcm_commonmode a_49402_66210# 0.30fF
C10867 a_32426_70226# a_32426_69222# 1.00fF
C10868 a_38450_18528# a_39454_18528# 0.97fF
C10869 vcm_commonmode a_23390_72234# 0.69fF
C10870 a_6559_59879# a_11877_50645# 0.60fF
C10871 a_29760_7638# VDD 6.61fF
C10872 vcm_commonmode a_26310_12870# 0.31fF
C10873 a_4528_26159# a_7059_24135# 0.96fF
C10874 a_18370_24552# a_19374_24552# 0.97fF
C10875 a_11947_68279# VDD 0.54fF
C10876 a_2289_35113# VDD 0.39fF
C10877 a_45478_67214# ctopp 3.59fF
C10878 a_43362_28879# a_47486_55166# 0.55fF
C10879 a_23685_29111# a_9529_28335# 0.41fF
C10880 a_36717_47375# a_36442_63198# 0.42fF
C10881 a_11067_67279# a_11067_66191# 0.46fF
C10882 a_20635_29415# a_22291_29415# 0.80fF
C10883 a_16863_29415# a_29927_29199# 0.88fF
C10884 a_17599_52263# a_22386_69222# 0.38fF
C10885 a_2419_48783# a_9135_49557# 0.61fF
C10886 a_30326_19898# a_30418_19532# 0.32fF
C10887 a_9872_20969# VDD 0.41fF
C10888 vcm_commonmode a_17366_7484# 0.69fF
C10889 a_31422_11500# a_31422_10496# 1.00fF
C10890 a_11067_67279# a_12895_13967# 23.49fF
C10891 a_1761_52815# a_19594_35823# 0.32fF
C10892 vcm_commonmode a_33430_58178# 0.87fF
C10893 a_1923_59583# a_4339_64521# 0.83fF
C10894 a_35346_14878# a_35438_14512# 0.32fF
C10895 vcm_commonmode a_21290_21906# 0.31fF
C10896 a_14039_41271# VDD 0.62fF
C10897 VDD config_2_in[1] 1.24fF
C10898 a_12663_35431# a_13005_35823# 2.67fF
C10899 a_22843_29415# a_21187_29415# 0.57fF
C10900 a_19374_17524# VDD 0.51fF
C10901 a_7251_50069# VDD 0.88fF
C10902 a_4482_57863# a_10687_52553# 0.34fF
C10903 a_12341_3311# a_12727_13353# 0.41fF
C10904 a_5363_30503# a_2787_30503# 0.55fF
C10905 a_8583_33551# a_15607_46805# 0.31fF
C10906 a_29414_55166# a_30418_55166# 0.97fF
C10907 a_2787_32679# a_6883_37019# 0.49fF
C10908 vcm_commonmode a_26310_17890# 0.31fF
C10909 a_20378_57174# a_21382_57174# 0.97fF
C10910 a_8575_74853# VDD 4.32fF
C10911 a_23390_15516# a_24394_15516# 0.97fF
C10912 a_24959_30503# a_26523_28111# 0.35fF
C10913 a_16707_44535# VDD 0.61fF
C10914 a_6559_22671# a_5671_21495# 0.82fF
C10915 a_3339_43023# a_4446_40553# 0.64fF
C10916 VDD config_2_in[9] 0.81fF
C10917 a_2327_54135# VDD 0.44fF
C10918 a_46482_63198# VDD 0.57fF
C10919 a_47486_10496# a_48490_10496# 0.97fF
C10920 a_2419_55687# VDD 1.12fF
C10921 a_49402_65206# a_49494_65206# 0.32fF
C10922 a_25447_36919# VDD 0.63fF
C10923 a_17507_52047# a_21382_55166# 0.46fF
C10924 a_12985_16367# a_12727_13353# 1.03fF
C10925 a_2467_48981# a_1761_49007# 0.44fF
C10926 a_4443_46607# VDD 16.34fF
C10927 a_21382_71230# a_22386_71230# 0.97fF
C10928 vcm_commonmode a_20378_69222# 0.87fF
C10929 a_40458_59182# VDD 0.51fF
C10930 vcm_commonmode a_47486_9492# 0.87fF
C10931 a_40366_23914# a_40458_23548# 0.32fF
C10932 a_6515_62037# VDD 3.76fF
C10933 a_20359_29199# a_41967_31375# 1.27fF
C10934 a_33430_11500# a_34434_11500# 0.97fF
C10935 a_11812_30511# VDD 0.35fF
C10936 a_44474_64202# ctopp 3.59fF
C10937 a_43362_28879# VDD 10.15fF
C10938 a_37354_66210# a_37446_66210# 0.32fF
C10939 vcm_commonmode a_47394_59182# 0.31fF
C10940 vcm_commonmode a_27406_22544# 0.87fF
C10941 a_2401_41941# VDD 0.32fF
C10942 vcm_commonmode a_18370_65206# 0.88fF
C10943 a_38557_32143# a_10975_66407# 0.40fF
C10944 a_8583_33551# a_77086_40693# 1.13fF
C10945 a_20378_18528# VDD 0.51fF
C10946 a_1923_54591# a_2163_54589# 0.32fF
C10947 a_12641_37684# a_12621_36091# 0.51fF
C10948 ctopn a_18370_8488# 3.39fF
C10949 a_37446_24552# a_38450_24552# 0.97fF
C10950 a_12341_3311# a_10515_23975# 0.46fF
C10951 a_49402_68218# VDD 0.31fF
C10952 a_2840_66103# a_2959_47113# 1.26fF
C10953 vcm_commonmode a_27314_18894# 0.31fF
C10954 a_20378_66210# ctopp 3.59fF
C10955 vcm_commonmode a_16362_61190# 4.47fF
C10956 a_5639_15279# a_5805_15279# 0.39fF
C10957 a_18703_29199# a_38067_47349# 0.52fF
C10958 a_16746_14510# VDD 33.20fF
C10959 a_7644_46805# VDD 0.97fF
C10960 a_49402_19898# a_49494_19532# 0.32fF
C10961 a_6467_55527# a_37534_51701# 0.46fF
C10962 a_6372_38279# a_5915_35943# 0.33fF
C10963 a_34434_62194# a_35438_62194# 0.97fF
C10964 vcm_commonmode a_23390_14512# 0.87fF
C10965 a_21479_38053# VDD 0.91fF
C10966 vcm_commonmode a_18278_55166# 0.31fF
C10967 a_29414_10496# VDD 0.51fF
C10968 a_2787_32679# a_3987_19623# 1.84fF
C10969 a_75111_40050# VDD 0.53fF
C10970 vcm_commonmode a_49494_64202# 0.91fF
C10971 a_20195_49793# VDD 0.47fF
C10972 a_25787_28327# a_12901_66665# 0.40fF
C10973 a_35601_27497# a_35438_15516# 0.38fF
C10974 a_10515_23975# a_12985_16367# 0.97fF
C10975 a_33338_20902# a_33430_20536# 0.32fF
C10976 a_44474_60186# VDD 0.51fF
C10977 a_1586_51335# a_8491_57487# 0.48fF
C10978 vcm_commonmode a_36350_10862# 0.31fF
C10979 a_22294_63198# a_22386_63198# 0.32fF
C10980 a_2223_28617# a_3143_22364# 0.43fF
C10981 a_14273_27791# a_12985_25615# 0.82fF
C10982 a_39454_57174# a_40458_57174# 0.97fF
C10983 a_1823_72381# VDD 3.02fF
C10984 a_1768_16367# a_2840_66103# 0.40fF
C10985 a_42466_15516# a_43470_15516# 0.97fF
C10986 vcm_commonmode a_28410_23548# 0.87fF
C10987 vcm_commonmode a_25398_66210# 0.87fF
C10988 a_2099_59861# a_1586_36727# 1.65fF
C10989 a_4311_52245# VDD 0.37fF
C10990 a_16746_62196# VDD 33.19fF
C10991 a_12447_29199# a_26523_29199# 0.31fF
C10992 a_16362_9492# a_16746_9490# 2.28fF
C10993 a_49402_56170# VDD 0.31fF
C10994 vcm_commonmode a_37446_19532# 0.87fF
C10995 a_42466_58178# a_42466_59182# 1.00fF
C10996 ctopn a_19374_16520# 3.59fF
C10997 vcm_commonmode a_23298_62194# 0.31fF
C10998 a_2235_30503# a_6243_30662# 0.32fF
C10999 a_27535_30503# a_7295_44647# 4.23fF
C11000 a_22843_29415# a_26523_28111# 0.90fF
C11001 a_24394_15516# VDD 0.51fF
C11002 a_40458_71230# a_41462_71230# 0.97fF
C11003 a_2124_57979# VDD 0.65fF
C11004 a_12901_58799# a_16746_59184# 0.41fF
C11005 a_19720_7638# a_12985_19087# 0.41fF
C11006 a_4903_29975# VDD 0.35fF
C11007 vcm_commonmode a_31330_15882# 0.31fF
C11008 a_24394_63198# ctopp 3.64fF
C11009 a_3949_41935# a_7244_39189# 1.15fF
C11010 a_22386_71230# VDD 0.58fF
C11011 a_29760_55394# a_12901_58799# 0.40fF
C11012 a_18045_39105# VDD 1.55fF
C11013 a_25398_72234# m3_25300_72146# 2.80fF
C11014 a_34434_11500# VDD 0.51fF
C11015 a_22632_41831# VDD 1.73fF
C11016 vcm_commonmode a_29322_71230# 0.31fF
C11017 a_5535_18012# a_6738_19783# 0.45fF
C11018 a_1761_39215# a_1761_34319# 0.48fF
C11019 a_38450_24552# VDD 0.60fF
C11020 vcm_commonmode a_41370_11866# 0.31fF
C11021 a_18370_59182# ctopp 3.58fF
C11022 a_4339_64521# a_10680_54171# 0.53fF
C11023 a_37919_28111# a_38450_22544# 0.38fF
C11024 a_12907_27023# a_4811_34855# 1.12fF
C11025 a_20378_64202# a_20378_63198# 1.23fF
C11026 a_33338_12870# a_33430_12504# 0.32fF
C11027 a_1987_31812# VDD 0.70fF
C11028 a_2317_28892# a_2223_28617# 0.95fF
C11029 vcm_commonmode a_45386_24918# 0.31fF
C11030 a_25787_28327# a_10680_52245# 0.38fF
C11031 a_3339_30503# a_15548_30761# 0.58fF
C11032 a_23395_52047# a_27406_68218# 0.38fF
C11033 a_28410_59182# a_28410_58178# 1.00fF
C11034 a_8295_47388# a_1586_45431# 0.41fF
C11035 a_49494_55166# VDD 1.25fF
C11036 a_12985_25615# VDD 0.88fF
C11037 a_40458_57174# VDD 0.51fF
C11038 a_19374_13508# a_20378_13508# 0.97fF
C11039 a_35033_37692# VDD 0.86fF
C11040 vcm_commonmode a_40458_20536# 0.87fF
C11041 a_1689_10396# a_2021_17973# 2.25fF
C11042 a_15871_39913# VDD 0.63fF
C11043 a_24394_68218# a_25398_68218# 0.97fF
C11044 a_28547_51175# a_12355_15055# 0.40fF
C11045 vcm_commonmode a_29414_63198# 0.92fF
C11046 vcm_commonmode a_47394_57174# 0.31fF
C11047 a_41261_28335# a_42466_71230# 0.38fF
C11048 a_16955_52047# a_12516_7093# 0.40fF
C11049 a_12341_3311# a_22386_15516# 0.38fF
C11050 a_16362_59182# VDD 2.48fF
C11051 a_36442_56170# a_36442_55166# 1.00fF
C11052 a_34434_24552# m3_34336_24702# 2.45fF
C11053 a_41370_63198# a_41462_63198# 0.32fF
C11054 a_30203_31055# VDD 0.32fF
C11055 a_15459_41781# a_12641_42036# 2.27fF
C11056 a_48490_58178# ctopp 3.43fF
C11057 a_32426_57174# a_32426_56170# 1.00fF
C11058 a_29322_72234# VDD 0.63fF
C11059 a_21371_50959# a_25398_60186# 0.38fF
C11060 vcm_commonmode a_23390_59182# 0.87fF
C11061 a_7815_42453# VDD 0.67fF
C11062 a_41427_52263# a_41462_67214# 0.38fF
C11063 a_28547_51175# a_31659_31751# 3.85fF
C11064 a_28318_21906# a_28410_21540# 0.32fF
C11065 a_12641_37684# a_12473_36341# 0.30fF
C11066 vcm_commonmode a_40458_12504# 0.87fF
C11067 a_22386_60186# ctopp 3.59fF
C11068 ctopn a_41462_9492# 3.58fF
C11069 a_25398_68218# VDD 0.51fF
C11070 a_6559_22671# a_6883_37019# 0.43fF
C11071 a_29177_34753# VDD 1.23fF
C11072 a_2021_17973# a_2004_42453# 2.32fF
C11073 a_25306_7850# VDD 0.63fF
C11074 a_46390_58178# a_46482_58178# 0.32fF
C11075 a_12727_13353# a_16362_15516# 19.89fF
C11076 a_23395_52047# a_27406_56170# 0.38fF
C11077 ctopn a_21382_22544# 3.58fF
C11078 vcm_commonmode a_32334_68218# 0.31fF
C11079 a_4379_18756# a_4075_18543# 0.48fF
C11080 a_35346_59182# a_35438_59182# 0.32fF
C11081 a_40491_27247# a_12985_19087# 0.41fF
C11082 a_7571_29199# a_14926_31849# 0.95fF
C11083 a_15607_46805# a_38210_30199# 0.37fF
C11084 a_49494_23548# m3_49396_23410# 2.78fF
C11085 a_13143_29575# VDD 1.24fF
C11086 a_21387_38591# VDD 0.82fF
C11087 a_11067_63143# a_5595_33205# 0.59fF
C11088 vcm_commonmode a_35438_21540# 0.87fF
C11089 a_1586_21959# config_1_in[14] 0.33fF
C11090 a_8017_40847# VDD 0.35fF
C11091 a_33338_17890# a_33430_17524# 0.32fF
C11092 a_27535_30503# a_11067_46823# 0.42fF
C11093 a_20286_60186# a_20378_60186# 0.32fF
C11094 a_40491_27247# a_43470_22544# 0.38fF
C11095 a_39454_64202# a_39454_63198# 1.23fF
C11096 a_40581_31599# VDD 1.81fF
C11097 vcm_commonmode a_40458_17524# 0.87fF
C11098 ctopn a_17366_14512# 3.43fF
C11099 a_32167_29611# a_32772_7638# 0.48fF
C11100 a_10221_74031# VDD 0.66fF
C11101 vcm_commonmode a_27406_60186# 0.87fF
C11102 a_39454_13508# VDD 0.51fF
C11103 a_42466_58178# a_42466_57174# 1.00fF
C11104 a_34823_44535# VDD 0.57fF
C11105 a_31422_22544# a_31422_21540# 1.00fF
C11106 a_7773_63927# a_8491_57487# 0.57fF
C11107 a_25398_56170# VDD 0.52fF
C11108 vcm_commonmode a_46390_13874# 0.31fF
C11109 a_38450_13508# a_39454_13508# 0.97fF
C11110 a_13097_36367# VDD 4.27fF
C11111 a_24800_43041# a_12381_43957# 3.16fF
C11112 a_1761_25071# a_1586_36727# 0.45fF
C11113 a_43470_68218# a_44474_68218# 0.97fF
C11114 a_1768_16367# a_1761_30511# 0.36fF
C11115 vcm_commonmode a_32334_56170# 0.31fF
C11116 a_31768_55394# a_12257_56623# 0.40fF
C11117 ctopn a_22386_23548# 3.40fF
C11118 a_12727_15529# VDD 7.20fF
C11119 a_29847_48734# VDD 0.47fF
C11120 a_26748_7638# a_26402_19532# 0.38fF
C11121 a_2411_26133# a_3137_37589# 0.39fF
C11122 a_25787_28327# a_19807_28111# 2.13fF
C11123 a_24394_56170# a_25398_56170# 0.97fF
C11124 a_18370_57174# ctopp 3.57fF
C11125 a_21371_52263# a_10515_22671# 0.44fF
C11126 ctopn a_31422_19532# 3.59fF
C11127 a_2235_30503# a_6162_28487# 0.51fF
C11128 a_9414_10383# VDD 0.37fF
C11129 a_37307_51339# VDD 0.71fF
C11130 a_19374_72234# a_20378_72234# 0.97fF
C11131 a_43270_27791# a_45478_16520# 0.38fF
C11132 a_47394_21906# a_47486_21540# 0.32fF
C11133 a_24394_61190# VDD 0.51fF
C11134 vcm_commonmode a_17366_11500# 1.82fF
C11135 a_28410_58178# a_28410_57174# 1.00fF
C11136 a_1770_14441# a_2099_59861# 7.22fF
C11137 vcm_commonmode a_41462_18528# 0.87fF
C11138 a_41334_29575# a_39727_27765# 0.44fF
C11139 a_28841_29575# a_27752_7638# 0.59fF
C11140 a_16152_43677# a_12641_43124# 0.88fF
C11141 vcm_commonmode a_31330_61190# 0.31fF
C11142 a_35438_16520# a_35438_15516# 1.00fF
C11143 vcm_commonmode a_21382_24552# 0.84fF
C11144 a_4500_45289# VDD 0.76fF
C11145 a_1923_73087# a_9135_67503# 0.35fF
C11146 a_20378_19532# a_20378_18528# 1.00fF
C11147 a_1689_10396# a_2411_19605# 0.54fF
C11148 a_2775_46025# a_10687_52553# 0.33fF
C11149 a_19720_7638# a_19374_18528# 0.38fF
C11150 a_18979_30287# a_19626_31751# 0.51fF
C11151 a_29927_29199# a_31084_30485# 0.67fF
C11152 a_10515_63143# a_10055_58791# 0.60fF
C11153 a_24302_10862# a_24394_10496# 0.32fF
C11154 a_16362_57174# VDD 2.48fF
C11155 a_32426_62194# ctopp 3.59fF
C11156 a_32772_7638# a_32426_24552# 0.42fF
C11157 a_28410_70226# VDD 0.51fF
C11158 vcm_commonmode a_16746_20534# 5.36fF
C11159 vcm_commonmode a_32334_55166# 0.31fF
C11160 a_17711_40183# VDD 0.59fF
C11161 vcm_commonmode a_23390_57174# 0.87fF
C11162 a_16863_29415# VDD 9.15fF
C11163 vcm_commonmode a_35346_70226# 0.31fF
C11164 a_1761_27791# a_7281_29423# 0.38fF
C11165 a_39362_60186# a_39454_60186# 0.32fF
C11166 a_12727_58255# a_10515_22671# 0.49fF
C11167 a_16362_23548# a_16746_23546# 2.28fF
C11168 a_22015_28111# a_41842_27221# 0.52fF
C11169 vcm_commonmode a_16362_16520# 4.47fF
C11170 a_10873_27497# a_7369_24233# 0.54fF
C11171 a_5975_71829# VDD 0.37fF
C11172 a_38450_71230# ctopp 3.40fF
C11173 ctopn a_34434_20536# 3.59fF
C11174 a_2787_30503# a_18162_31055# 0.46fF
C11175 a_18662_43671# VDD 1.15fF
C11176 a_41261_28335# a_12983_63151# 0.40fF
C11177 a_34342_18894# a_34434_18528# 0.32fF
C11178 a_13123_38231# a_13005_35823# 1.99fF
C11179 a_4298_58951# a_7313_53047# 0.59fF
C11180 a_16362_21540# a_12985_7663# 1.27fF
C11181 a_1823_76181# a_5682_69367# 1.04fF
C11182 a_12907_27023# a_11902_27497# 0.96fF
C11183 a_23390_61190# a_24394_61190# 0.97fF
C11184 a_7749_55535# VDD 1.09fF
C11185 a_10055_58791# a_35601_27497# 0.41fF
C11186 vcm_commonmode a_16746_12502# 5.36fF
C11187 a_2125_68053# VDD 0.66fF
C11188 a_21859_35831# VDD 0.64fF
C11189 a_5085_23047# config_1_in[13] 0.39fF
C11190 a_41872_29423# a_43470_55166# 0.52fF
C11191 a_46482_8488# VDD 0.58fF
C11192 a_39299_48783# a_12981_62313# 0.40fF
C11193 vcm_commonmode a_37446_62194# 0.87fF
C11194 a_28547_51175# a_32426_63198# 0.42fF
C11195 a_29414_68218# a_29414_67214# 1.00fF
C11196 a_22015_28111# a_34221_47695# 0.44fF
C11197 a_14287_51175# a_18370_69222# 0.38fF
C11198 a_17366_58178# VDD 0.57fF
C11199 a_23685_29111# VDD 1.05fF
C11200 vcm_commonmode a_45478_15516# 0.87fF
C11201 ctopn a_34434_12504# 3.59fF
C11202 a_16955_52047# a_15607_46805# 0.43fF
C11203 a_43470_56170# a_44474_56170# 0.97fF
C11204 vcm_commonmode a_24302_58178# 0.31fF
C11205 a_4674_40277# a_2021_22325# 0.45fF
C11206 a_13107_41317# VDD 0.94fF
C11207 a_12713_36483# a_13669_35253# 3.88fF
C11208 a_27869_50095# a_29147_50069# 0.32fF
C11209 a_34780_56398# a_34434_72234# 0.34fF
C11210 vcm_commonmode a_43470_71230# 0.86fF
C11211 a_24740_7638# a_24394_15516# 0.38fF
C11212 a_25306_55166# a_25398_55166# 0.32fF
C11213 a_26402_8488# a_27406_8488# 0.97fF
C11214 a_34434_67214# VDD 0.51fF
C11215 vcm_commonmode a_12899_11471# 6.31fF
C11216 a_19282_15882# a_19374_15516# 0.32fF
C11217 ctopn a_29414_21540# 3.59fF
C11218 a_43267_31055# a_12727_67753# 0.40fF
C11219 a_27406_70226# a_28410_70226# 0.97fF
C11220 vcm_commonmode a_41370_67214# 0.31fF
C11221 a_39454_19532# a_39454_18528# 1.00fF
C11222 a_43378_10862# a_43470_10496# 0.32fF
C11223 vcm_commonmode a_22386_13508# 0.87fF
C11224 a_9485_69141# VDD 0.66fF
C11225 a_41462_68218# ctopp 3.59fF
C11226 ctopn a_34434_17524# 3.59fF
C11227 a_1591_29973# a_1895_30138# 0.39fF
C11228 a_31422_9492# VDD 0.51fF
C11229 a_47486_16520# VDD 0.51fF
C11230 a_3983_48469# VDD 0.44fF
C11231 a_21371_50959# a_4351_67279# 0.40fF
C11232 a_17274_71230# a_17366_71230# 0.32fF
C11233 ctopn a_39223_32463# 2.62fF
C11234 a_25398_60186# a_25398_59182# 1.00fF
C11235 vcm_commonmode a_38358_9858# 0.31fF
C11236 a_34482_29941# a_40581_31599# 1.00fF
C11237 a_29322_11866# a_29414_11500# 0.32fF
C11238 a_39222_48169# VDD 7.32fF
C11239 a_34434_15516# a_34434_14512# 1.00fF
C11240 a_4429_14191# a_1929_10651# 0.40fF
C11241 vcm_commonmode a_18278_22910# 0.31fF
C11242 vcm_commonmode m3_16264_58090# 3.21fF
C11243 a_2235_30503# a_9529_28335# 2.09fF
C11244 a_31768_55394# a_10975_66407# 0.40fF
C11245 a_13835_36649# a_12713_36483# 0.43fF
C11246 a_5135_50069# VDD 0.90fF
C11247 vcm_commonmode a_40050_48463# 10.13fF
C11248 a_42466_61190# a_43470_61190# 0.97fF
C11249 a_19374_9492# a_19374_8488# 1.00fF
C11250 a_33338_24918# a_33430_24552# 0.33fF
C11251 a_21948_34973# VDD 1.45fF
C11252 a_12263_4391# a_9731_22895# 1.49fF
C11253 a_39454_7484# VDD 1.23fF
C11254 a_2021_22325# a_6607_42167# 1.43fF
C11255 a_48490_68218# a_48490_67214# 1.00fF
C11256 a_23395_52047# a_6467_55527# 0.34fF
C11257 a_42985_46831# a_12901_66959# 0.40fF
C11258 vcm_commonmode a_46482_68218# 0.87fF
C11259 a_1770_14441# a_1761_25071# 0.70fF
C11260 a_33430_64202# VDD 0.51fF
C11261 a_30326_62194# a_30418_62194# 0.32fF
C11262 a_25787_28327# a_29927_29199# 8.54fF
C11263 a_26433_39631# a_30115_38695# 0.36fF
C11264 a_41462_56170# ctopp 3.40fF
C11265 ctopn a_35438_18528# 3.59fF
C11266 a_20839_41001# VDD 0.57fF
C11267 a_33430_69222# a_33430_68218# 1.00fF
C11268 vcm_commonmode a_40366_64202# 0.31fF
C11269 a_8569_49007# VDD 1.04fF
C11270 a_21371_52263# a_12901_66665# 0.40fF
C11271 a_43378_55166# a_43470_55166# 0.32fF
C11272 a_45478_8488# a_46482_8488# 0.97fF
C11273 a_23390_8488# a_23390_7484# 1.00fF
C11274 a_17927_31573# VDD 0.52fF
C11275 a_35346_57174# a_35438_57174# 0.32fF
C11276 a_2124_73211# VDD 0.58fF
C11277 a_1950_59887# a_9577_60437# 0.43fF
C11278 a_38358_15882# a_38450_15516# 0.32fF
C11279 vcm_commonmode a_19282_23914# 0.31fF
C11280 vcm_commonmode a_12355_65103# 6.25fF
C11281 a_46482_70226# a_47486_70226# 0.97fF
C11282 a_4891_47388# a_4563_32900# 0.47fF
C11283 a_21382_19532# VDD 0.51fF
C11284 a_7217_53047# VDD 0.68fF
C11285 a_19720_7638# VDD 6.42fF
C11286 a_40458_61190# ctopp 3.59fF
C11287 ctopn a_44474_10496# 3.59fF
C11288 a_42466_69222# VDD 0.51fF
C11289 a_33727_36649# VDD 0.66fF
C11290 vcm_commonmode a_28318_19898# 0.31fF
C11291 a_25787_28327# a_33430_55166# 0.42fF
C11292 a_1803_20719# a_6269_43567# 0.51fF
C11293 a_27406_16520# a_28410_16520# 0.97fF
C11294 a_25787_28327# a_28817_29111# 0.38fF
C11295 vcm_commonmode a_46482_56170# 0.87fF
C11296 a_4811_34855# a_4903_31849# 0.95fF
C11297 a_13643_28327# a_18703_29199# 0.54fF
C11298 a_6435_47893# VDD 0.51fF
C11299 a_36350_71230# a_36442_71230# 0.32fF
C11300 vcm_commonmode a_49402_69222# 0.30fF
C11301 a_44474_60186# a_44474_59182# 1.00fF
C11302 a_49494_22544# VDD 1.10fF
C11303 vcm_commonmode a_29414_8488# 0.86fF
C11304 a_35601_27497# a_35438_20536# 0.38fF
C11305 a_27752_7638# a_27406_18528# 0.38fF
C11306 a_40458_65206# VDD 0.51fF
C11307 a_33430_63198# a_33430_62194# 1.00fF
C11308 a_48398_11866# a_48490_11500# 0.32fF
C11309 a_1586_51335# a_7479_54439# 0.65fF
C11310 a_12947_71576# VDD 4.33fF
C11311 a_17599_52263# a_12901_58799# 0.40fF
C11312 a_44474_70226# ctopp 3.58fF
C11313 a_5098_41641# VDD 1.03fF
C11314 vcm_commonmode a_47394_65206# 0.31fF
C11315 a_25306_72234# a_25398_72234# 0.32fF
C11316 a_24740_7638# a_12727_15529# 0.41fF
C11317 a_6559_22671# a_7369_24233# 0.39fF
C11318 a_38450_9492# a_38450_8488# 1.00fF
C11319 a_29322_24918# VDD 0.36fF
C11320 a_31768_7638# a_31422_21540# 0.38fF
C11321 a_20359_29199# a_3339_30503# 0.48fF
C11322 ctopn a_39454_15516# 3.59fF
C11323 vcm_commonmode a_45478_61190# 0.87fF
C11324 a_33430_67214# a_34434_67214# 0.97fF
C11325 a_18151_52263# a_3339_43023# 0.55fF
C11326 a_21371_52263# a_10680_52245# 0.77fF
C11327 a_45478_14512# VDD 0.51fF
C11328 vcm_commonmode a_17366_67214# 1.83fF
C11329 a_18611_52047# a_23390_68218# 0.38fF
C11330 a_35601_27497# a_35438_12504# 0.38fF
C11331 a_2411_26133# a_3972_25615# 0.60fF
C11332 a_24394_20536# VDD 0.51fF
C11333 a_39362_55166# VDD 0.35fF
C11334 a_4314_40821# a_4495_35925# 0.55fF
C11335 a_49402_62194# a_49494_62194# 0.32fF
C11336 vcm_commonmode a_31330_20902# 0.31fF
C11337 a_11067_13095# a_6752_29941# 0.39fF
C11338 a_7078_36103# VDD 1.10fF
C11339 a_20286_68218# a_20378_68218# 0.32fF
C11340 a_21371_50959# a_12355_15055# 0.40fF
C11341 vcm_commonmode a_20286_63198# 0.31fF
C11342 vcm_commonmode a_49494_70226# 0.90fF
C11343 a_1950_59887# a_8958_65961# 0.52fF
C11344 a_38557_32143# a_38450_71230# 0.38fF
C11345 a_19374_7484# a_20378_7484# 0.97fF
C11346 a_42466_8488# a_42466_7484# 1.00fF
C11347 a_33430_58178# ctopp 3.59fF
C11348 a_47486_66210# VDD 0.51fF
C11349 a_27406_24552# m3_27308_24414# 2.81fF
C11350 vcm_commonmode a_30418_16520# 0.87fF
C11351 ctopn a_16362_13508# 1.35fF
C11352 a_22294_72234# VDD 0.62fF
C11353 a_17507_52047# a_21382_60186# 0.38fF
C11354 a_23395_32463# a_33641_29967# 1.05fF
C11355 a_24394_12504# VDD 0.51fF
C11356 a_36613_48169# a_37446_67214# 0.38fF
C11357 a_35438_58178# a_36442_58178# 0.97fF
C11358 a_25517_37455# a_12473_36341# 0.90fF
C11359 a_12683_51329# VDD 0.52fF
C11360 a_35601_27497# a_35438_17524# 0.38fF
C11361 a_1823_76181# a_1586_66567# 0.54fF
C11362 a_30418_9492# a_31422_9492# 0.97fF
C11363 a_40491_27247# VDD 6.31fF
C11364 vcm_commonmode a_31330_12870# 0.31fF
C11365 a_16746_68220# VDD 33.19fF
C11366 a_31422_13508# a_31422_12504# 1.00fF
C11367 a_16928_35303# VDD 1.63fF
C11368 a_46482_16520# a_47486_16520# 0.97fF
C11369 vcm_commonmode ctopp 97.05fF
C11370 a_18611_52047# a_23390_56170# 0.38fF
C11371 a_12907_56399# a_12257_56623# 0.35fF
C11372 a_6727_47607# VDD 0.59fF
C11373 a_19374_21540# VDD 0.51fF
C11374 vcm_commonmode a_22386_7484# 0.69fF
C11375 a_4758_45369# a_19576_51701# 0.31fF
C11376 a_12341_3311# a_22386_20536# 0.38fF
C11377 a_51714_39886# a_51936_39932# 0.53fF
C11378 a_23736_7638# a_11067_21583# 0.41fF
C11379 vcm_commonmode a_26310_21906# 0.31fF
C11380 a_20378_69222# ctopp 3.59fF
C11381 a_2606_41079# a_2339_38129# 0.36fF
C11382 a_23415_41263# VDD 1.46fF
C11383 vcm_commonmode a_16746_64204# 5.37fF
C11384 vcm_commonmode a_44382_58178# 0.31fF
C11385 a_24394_17524# VDD 0.51fF
C11386 a_17682_50095# VDD 4.05fF
C11387 a_49402_24918# a_49494_24552# 0.32fF
C11388 vcm_commonmode a_31330_17890# 0.31fF
C11389 a_18370_65206# ctopp 3.58fF
C11390 a_1803_19087# a_13909_41923# 2.10fF
C11391 a_21382_67214# a_21382_66210# 1.00fF
C11392 vcm_commonmode a_18278_60186# 0.31fF
C11393 a_25263_44535# VDD 0.60fF
C11394 a_12341_3311# a_22386_12504# 0.38fF
C11395 a_8295_47388# a_9989_46831# 0.53fF
C11396 a_5179_74031# a_1923_73087# 0.31fF
C11397 a_16362_61190# ctopp 1.35fF
C11398 a_17366_65206# a_17366_64202# 1.00fF
C11399 a_34342_13874# a_34434_13508# 0.32fF
C11400 a_32971_35281# VDD 1.95fF
C11401 a_13183_52047# a_12981_62313# 0.40fF
C11402 a_39362_68218# a_39454_68218# 0.32fF
C11403 a_18151_52263# a_12257_56623# 0.40fF
C11404 a_2830_15431# VDD 0.38fF
C11405 vcm_commonmode a_25398_69222# 0.87fF
C11406 a_2419_48783# a_11711_50645# 0.52fF
C11407 a_14287_51175# a_5915_30287# 0.51fF
C11408 a_45478_59182# VDD 0.51fF
C11409 a_38450_7484# a_39454_7484# 0.97fF
C11410 a_32772_7638# a_12985_19087# 0.41fF
C11411 a_16362_65206# VDD 2.48fF
C11412 a_31084_30485# VDD 0.96fF
C11413 a_21371_52263# a_19807_28111# 0.32fF
C11414 a_6773_27805# a_7461_27247# 0.76fF
C11415 a_20286_56170# a_20378_56170# 0.32fF
C11416 a_19720_55394# a_10515_22671# 0.40fF
C11417 vcm_commonmode a_32426_22544# 0.87fF
C11418 a_3949_41935# VDD 4.04fF
C11419 a_22386_69222# a_23390_69222# 0.97fF
C11420 vcm_commonmode a_23390_65206# 0.87fF
C11421 a_2411_18517# a_10239_16367# 0.35fF
C11422 a_25398_18528# VDD 0.51fF
C11423 a_12341_3311# a_22386_17524# 0.38fF
C11424 a_17366_61190# a_17366_60186# 1.00fF
C11425 ctopn a_23390_8488# 3.40fF
C11426 a_32426_64202# a_33430_64202# 0.97fF
C11427 a_5346_33775# VDD 0.77fF
C11428 vcm_commonmode a_32334_18894# 0.31fF
C11429 a_25398_66210# ctopp 3.59fF
C11430 a_17311_46833# VDD 0.42fF
C11431 a_29414_22544# a_30418_22544# 0.97fF
C11432 a_30023_41959# a_30757_37455# 0.77fF
C11433 a_7571_29199# a_17358_31069# 0.43fF
C11434 a_6467_55527# a_7829_60431# 0.44fF
C11435 a_12899_3311# VDD 7.98fF
C11436 vcm_commonmode a_28410_14512# 0.87fF
C11437 a_20378_65206# a_21382_65206# 0.97fF
C11438 vcm_commonmode a_23298_55166# 0.30fF
C11439 a_34434_10496# VDD 0.51fF
C11440 a_12899_11471# a_16362_16520# 19.89fF
C11441 a_2011_34837# a_2235_30503# 0.99fF
C11442 a_49494_60186# VDD 1.14fF
C11443 a_2775_46025# a_1923_54591# 0.45fF
C11444 vcm_commonmode a_41370_10862# 0.31fF
C11445 a_20378_56170# a_20378_55166# 1.00fF
C11446 a_1768_13103# config_2_in[12] 0.79fF
C11447 a_39244_41953# a_38011_42035# 0.78fF
C11448 a_1761_43567# a_33856_40743# 0.45fF
C11449 a_6913_72399# VDD 0.58fF
C11450 a_3024_67191# a_8994_63927# 0.38fF
C11451 a_40458_67214# a_40458_66210# 1.00fF
C11452 a_7803_55509# a_7987_64213# 0.66fF
C11453 vcm_commonmode a_33430_23548# 0.87fF
C11454 a_11711_12559# VDD 0.45fF
C11455 vcm_commonmode a_30418_66210# 0.87fF
C11456 a_34251_52263# a_12983_63151# 0.40fF
C11457 VDD dummypin[0] 0.64fF
C11458 a_24683_51183# a_24849_51183# 0.66fF
C11459 a_21382_62194# VDD 0.51fF
C11460 a_12355_15055# a_2419_48783# 0.61fF
C11461 a_19282_61190# a_19374_61190# 0.32fF
C11462 a_12349_25847# VDD 2.61fF
C11463 a_36442_65206# a_36442_64202# 1.00fF
C11464 a_14735_35805# VDD 1.49fF
C11465 vcm_commonmode a_42466_19532# 0.87fF
C11466 ctopn a_24394_16520# 3.59fF
C11467 a_39389_52271# a_39454_55166# 0.46fF
C11468 a_2787_30503# a_17712_7638# 0.39fF
C11469 a_36613_48169# a_12981_62313# 0.40fF
C11470 vcm_commonmode a_28318_62194# 0.31fF
C11471 a_28756_55394# a_28410_63198# 0.42fF
C11472 a_29414_15516# VDD 0.51fF
C11473 a_20378_19532# a_21382_19532# 0.97fF
C11474 a_4503_21523# VDD 0.47fF
C11475 a_37919_28111# a_12985_19087# 0.41fF
C11476 a_30418_23548# a_30418_22544# 1.00fF
C11477 a_24893_37429# a_25091_37782# 0.30fF
C11478 a_3295_62083# a_1952_60431# 0.62fF
C11479 a_11395_62037# a_11299_62215# 0.36fF
C11480 vcm_commonmode a_36350_15882# 0.31fF
C11481 a_29414_63198# ctopp 3.64fF
C11482 a_39362_56170# a_39454_56170# 0.32fF
C11483 a_27406_71230# VDD 0.58fF
C11484 a_24394_66210# a_24394_65206# 1.00fF
C11485 a_25398_14512# a_26402_14512# 0.97fF
C11486 a_24413_39087# VDD 1.18fF
C11487 a_11067_66191# a_1586_21959# 1.33fF
C11488 a_28410_72234# m3_28312_72146# 2.80fF
C11489 a_39454_11500# VDD 0.51fF
C11490 a_12907_56399# a_10975_66407# 4.82fF
C11491 a_41462_69222# a_42466_69222# 0.97fF
C11492 ctopn a_42718_27497# 2.63fF
C11493 a_10239_16911# VDD 0.41fF
C11494 vcm_commonmode a_34342_71230# 0.31fF
C11495 a_12546_22351# a_2411_18517# 0.56fF
C11496 a_36442_61190# a_36442_60186# 1.00fF
C11497 a_22294_8854# a_22386_8488# 0.32fF
C11498 a_43470_24552# VDD 0.60fF
C11499 vcm_commonmode a_46390_11866# 0.31fF
C11500 a_23390_59182# ctopp 3.59fF
C11501 a_39673_28111# a_40458_22544# 0.38fF
C11502 a_14354_32117# VDD 1.25fF
C11503 a_1761_52815# a_12251_39069# 0.36fF
C11504 a_2847_44629# VDD 0.37fF
C11505 a_23298_70226# a_23390_70226# 0.32fF
C11506 a_39389_52271# a_12727_67753# 0.40fF
C11507 a_40366_58178# a_40458_58178# 0.32fF
C11508 a_48490_22544# a_49494_22544# 0.97fF
C11509 a_22386_62194# a_22386_61190# 1.00fF
C11510 a_1683_27399# VDD 0.52fF
C11511 a_45478_57174# VDD 0.51fF
C11512 a_7210_55081# a_8453_51727# 0.35fF
C11513 a_39454_65206# a_40458_65206# 0.97fF
C11514 a_4351_67279# a_6559_59663# 1.56fF
C11515 a_1591_36501# VDD 0.44fF
C11516 vcm_commonmode a_45478_20536# 0.87fF
C11517 a_15193_44005# a_12621_44099# 0.46fF
C11518 a_14258_44527# a_22632_42919# 0.56fF
C11519 a_1761_25071# a_2021_17973# 1.13fF
C11520 a_3339_43023# a_1761_34319# 6.82fF
C11521 a_1761_47919# a_13909_41923# 3.46fF
C11522 a_22448_39429# VDD 1.65fF
C11523 vcm_commonmode a_34434_63198# 0.92fF
C11524 a_35438_17524# a_35438_16520# 1.00fF
C11525 a_32135_49007# VDD 0.33fF
C11526 a_22386_20536# a_22386_19532# 1.00fF
C11527 a_2007_20149# VDD 0.84fF
C11528 a_24740_7638# a_24394_20536# 0.38fF
C11529 a_30418_23548# a_31422_23548# 0.97fF
C11530 a_1823_63677# a_2775_46025# 1.41fF
C11531 a_10055_58791# a_41967_31375# 0.41fF
C11532 a_28817_29111# a_37919_28111# 0.52fF
C11533 a_4960_40847# a_5490_41365# 0.78fF
C11534 a_12641_42036# a_13909_41923# 1.31fF
C11535 a_25787_28327# VDD 13.65fF
C11536 vcm_commonmode a_28410_59182# 0.87fF
C11537 a_27406_66210# a_28410_66210# 0.97fF
C11538 a_30788_28487# a_32823_29397# 0.37fF
C11539 a_15959_42943# VDD 0.96fF
C11540 a_18151_52263# a_10975_66407# 0.49fF
C11541 a_17599_52263# a_2840_66103# 0.32fF
C11542 vcm_commonmode a_38557_32143# 10.02fF
C11543 a_5190_59575# a_10687_52553# 0.57fF
C11544 a_4792_20443# a_5825_20495# 0.79fF
C11545 a_1799_29556# a_2473_34293# 2.44fF
C11546 a_38358_61190# a_38450_61190# 0.32fF
C11547 vcm_commonmode a_45478_12504# 0.87fF
C11548 a_27406_60186# ctopp 3.59fF
C11549 ctopn a_46482_9492# 3.58fF
C11550 a_30418_68218# VDD 0.51fF
C11551 a_2235_30503# VDD 11.16fF
C11552 a_1768_16367# a_1761_25615# 0.42fF
C11553 a_30326_7850# VDD 0.62fF
C11554 a_16955_52047# a_6467_55527# 1.25fF
C11555 ctopn a_26402_22544# 3.58fF
C11556 a_11067_46823# a_7295_44647# 0.52fF
C11557 a_27406_71230# a_27406_70226# 1.00fF
C11558 a_41427_52263# a_12901_66959# 0.40fF
C11559 vcm_commonmode a_37354_68218# 0.31fF
C11560 a_41967_31375# a_42466_9492# 0.38fF
C11561 a_39454_19532# a_40458_19532# 0.97fF
C11562 a_24740_7638# a_24394_12504# 0.38fF
C11563 a_49494_23548# a_49494_22544# 1.00fF
C11564 a_43470_66210# a_43470_65206# 1.00fF
C11565 a_44474_14512# a_45478_14512# 0.97fF
C11566 vcm_commonmode a_40458_21540# 0.87fF
C11567 a_11619_56615# a_12349_25847# 0.71fF
C11568 a_11179_9981# VDD 0.49fF
C11569 a_19720_55394# a_12901_66665# 0.40fF
C11570 a_44474_72234# a_45478_72234# 0.97fF
C11571 a_23390_20536# a_24394_20536# 0.97fF
C11572 a_35601_27497# a_12877_14441# 0.41fF
C11573 a_41370_8854# a_41462_8488# 0.32fF
C11574 vcm_commonmode a_17366_10496# 1.82fF
C11575 a_2847_66389# VDD 0.35fF
C11576 vcm_commonmode a_45478_17524# 0.87fF
C11577 ctopn a_22386_14512# 3.59fF
C11578 a_10873_27497# a_17222_27247# 0.60fF
C11579 vcm_commonmode a_32426_60186# 0.87fF
C11580 a_44474_13508# VDD 0.51fF
C11581 a_12549_44212# VDD 3.42fF
C11582 a_42374_70226# a_42466_70226# 0.32fF
C11583 a_8295_47388# a_21169_49007# 0.58fF
C11584 a_2872_44111# a_18335_50645# 0.34fF
C11585 a_40675_27791# a_12877_16911# 0.41fF
C11586 a_24740_7638# a_24394_17524# 0.38fF
C11587 a_6831_63303# a_4298_58951# 0.56fF
C11588 a_41462_62194# a_41462_61190# 1.00fF
C11589 a_1586_51335# a_6559_59879# 0.53fF
C11590 a_32426_10496# a_32426_9492# 1.00fF
C11591 a_30418_56170# VDD 0.52fF
C11592 a_10055_58791# a_33864_28111# 0.41fF
C11593 a_20623_36595# VDD 2.12fF
C11594 a_3668_56311# a_6138_54599# 0.42fF
C11595 a_3339_43023# a_3339_30503# 1.07fF
C11596 a_23298_16886# a_23390_16520# 0.32fF
C11597 vcm_commonmode a_37354_56170# 0.31fF
C11598 ctopn a_27406_23548# 3.40fF
C11599 a_8123_14741# VDD 0.47fF
C11600 a_41462_20536# a_41462_19532# 1.00fF
C11601 vcm_commonmode a_20286_8854# 0.31fF
C11602 a_22015_28111# a_32823_29397# 0.62fF
C11603 a_17222_27247# a_19889_27497# 0.95fF
C11604 a_13909_41923# a_23789_39100# 1.34fF
C11605 a_23390_57174# ctopp 3.58fF
C11606 a_1757_71317# VDD 0.61fF
C11607 a_46482_66210# a_47486_66210# 0.97fF
C11608 ctopn a_36442_19532# 3.59fF
C11609 a_2235_30503# a_18053_28879# 0.57fF
C11610 a_30052_32117# a_30565_30199# 0.60fF
C11611 vcm_commonmode m3_16264_19394# 3.21fF
C11612 a_34699_42035# VDD 1.62fF
C11613 a_40050_48463# a_12355_65103# 0.40fF
C11614 a_10975_66407# a_9642_10357# 0.30fF
C11615 a_21382_21540# a_21382_20536# 1.00fF
C11616 a_9503_26151# a_20378_16520# 0.38fF
C11617 a_29414_61190# VDD 0.51fF
C11618 a_12907_27023# a_10964_25615# 0.70fF
C11619 vcm_commonmode a_22386_11500# 0.87fF
C11620 a_39673_28111# a_11067_21583# 0.41fF
C11621 a_10391_67477# VDD 0.35fF
C11622 a_23390_12504# a_24394_12504# 0.97fF
C11623 a_38454_34191# VDD 0.48fF
C11624 vcm_commonmode a_46482_18528# 0.87fF
C11625 a_29322_67214# a_29414_67214# 0.32fF
C11626 vcm_commonmode a_36350_61190# 0.31fF
C11627 vcm_commonmode a_26402_24552# 0.84fF
C11628 a_19720_55394# a_19374_68218# 0.38fF
C11629 a_46482_71230# a_46482_70226# 1.00fF
C11630 a_3339_43023# a_13835_43177# 0.57fF
C11631 a_2124_63419# VDD 0.64fF
C11632 a_5490_41365# a_1761_30511# 0.48fF
C11633 a_10055_58791# a_42709_29199# 0.40fF
C11634 a_37446_62194# ctopp 3.59fF
C11635 a_33430_70226# VDD 0.51fF
C11636 a_1761_37039# VDD 8.10fF
C11637 vcm_commonmode a_36442_55166# 0.84fF
C11638 a_1761_25071# a_1761_22895# 9.74fF
C11639 a_1761_46287# a_12381_43957# 0.63fF
C11640 a_14287_51175# a_12355_15055# 1.44fF
C11641 vcm_commonmode a_28410_57174# 0.87fF
C11642 a_13809_48463# VDD 0.40fF
C11643 vcm_commonmode a_40366_70226# 0.31fF
C11644 a_34780_56398# a_34434_71230# 0.38fF
C11645 a_42466_20536# a_43470_20536# 0.97fF
C11646 VDD config_1_in[13] 2.49fF
C11647 a_20378_24552# m3_20280_24414# 2.81fF
C11648 a_31422_63198# a_32426_63198# 0.97fF
C11649 a_5441_27791# VDD 0.64fF
C11650 vcm_commonmode a_21290_16886# 0.31fF
C11651 a_31768_55394# a_27535_30503# 0.77fF
C11652 a_39223_32463# a_39454_23548# 0.38fF
C11653 a_8485_71855# VDD 0.52fF
C11654 a_40050_48463# a_45478_61190# 0.38fF
C11655 a_11710_58487# a_11053_62607# 0.56fF
C11656 a_43470_71230# ctopp 3.40fF
C11657 ctopn a_39454_20536# 3.59fF
C11658 a_25787_28327# a_33430_67214# 0.38fF
C11659 a_31330_58178# a_31422_58178# 0.32fF
C11660 a_29361_51727# VDD 3.45fF
C11661 a_18370_21540# a_19374_21540# 0.97fF
C11662 a_1803_19087# a_1683_31599# 0.33fF
C11663 a_26310_9858# a_26402_9492# 0.32fF
C11664 a_10055_58791# a_9503_26151# 0.41fF
C11665 a_1761_32143# VDD 7.53fF
C11666 vcm_commonmode a_42466_62194# 0.87fF
C11667 a_42374_16886# a_42466_16520# 0.32fF
C11668 vcm_commonmode a_35601_27497# 10.35fF
C11669 a_19720_55394# a_19374_56170# 0.38fF
C11670 a_7939_30503# a_13357_32143# 0.47fF
C11671 a_16863_29415# a_24959_30503# 1.18fF
C11672 a_1923_73087# a_10010_68021# 0.30fF
C11673 a_22386_58178# VDD 0.51fF
C11674 a_25398_59182# a_26402_59182# 0.97fF
C11675 a_8491_41383# a_14298_32143# 0.52fF
C11676 a_12663_39783# a_16043_38825# 0.49fF
C11677 a_6095_44807# a_8199_58229# 0.45fF
C11678 ctopn a_39454_12504# 3.59fF
C11679 a_25787_28327# a_34482_29941# 0.52fF
C11680 a_23736_7638# a_12546_22351# 0.41fF
C11681 a_13349_37973# a_12663_39783# 0.81fF
C11682 vcm_commonmode a_29322_58178# 0.31fF
C11683 vcm_commonmode a_12985_7663# 6.29fF
C11684 a_23390_17524# a_24394_17524# 0.97fF
C11685 vcm_commonmode a_48490_71230# 0.85fF
C11686 a_40458_21540# a_40458_20536# 1.00fF
C11687 a_11480_23957# VDD 0.41fF
C11688 a_27406_24552# a_27406_23548# 1.00fF
C11689 a_9955_20969# a_6816_19355# 0.36fF
C11690 a_25744_7638# a_25398_22544# 0.38fF
C11691 a_8491_27023# a_18370_22544# 0.38fF
C11692 a_5531_22895# a_4798_23759# 0.51fF
C11693 a_39454_67214# VDD 0.51fF
C11694 a_42466_12504# a_43470_12504# 0.97fF
C11695 a_7901_74281# VDD 0.67fF
C11696 a_48398_67214# a_48490_67214# 0.32fF
C11697 a_40050_48463# ctopp 2.63fF
C11698 ctopn a_34434_21540# 3.59fF
C11699 a_7862_34025# a_14625_30761# 0.37fF
C11700 a_5043_44085# VDD 0.35fF
C11701 vcm_commonmode a_46390_67214# 0.31fF
C11702 a_11067_67279# a_7841_12167# 0.37fF
C11703 a_7313_53047# VDD 0.43fF
C11704 a_1591_72943# a_1591_64239# 0.53fF
C11705 a_11067_13095# a_4674_40277# 1.08fF
C11706 a_29760_7638# a_29414_18528# 0.38fF
C11707 a_32772_7638# VDD 6.17fF
C11708 vcm_commonmode a_27406_13508# 0.87fF
C11709 a_16707_36919# VDD 0.62fF
C11710 a_46482_68218# ctopp 3.59fF
C11711 ctopn a_39454_17524# 3.59fF
C11712 a_36442_9492# VDD 0.51fF
C11713 a_4191_33449# a_17488_48731# 0.75fF
C11714 vcm_commonmode a_16746_69224# 5.36fF
C11715 a_34342_7850# a_34434_7484# 0.32fF
C11716 a_16746_22542# VDD 33.20fF
C11717 vcm_commonmode a_43378_9858# 0.31fF
C11718 a_10073_23439# a_10526_22057# 0.73fF
C11719 a_18979_30287# a_7939_30503# 0.88fF
C11720 a_15607_46805# a_32367_28309# 0.50fF
C11721 vcm_commonmode a_23298_22910# 0.31fF
C11722 a_1761_52815# a_1799_29556# 0.93fF
C11723 a_41167_42943# VDD 0.90fF
C11724 a_18278_69222# a_18370_69222# 0.32fF
C11725 a_24394_18528# a_24394_17524# 1.00fF
C11726 a_12473_37429# a_13669_35253# 0.41fF
C11727 a_17039_51157# a_4191_33449# 0.51fF
C11728 a_16362_18528# VDD 2.47fF
C11729 a_13183_52047# a_17366_72234# 0.34fF
C11730 a_37446_21540# a_38450_21540# 0.97fF
C11731 a_45386_9858# a_45478_9492# 0.32fF
C11732 a_6567_25615# VDD 0.39fF
C11733 a_28318_64202# a_28410_64202# 0.32fF
C11734 a_12355_65103# ctopp 3.23fF
C11735 a_44474_7484# VDD 1.25fF
C11736 a_7695_31573# a_8461_32937# 0.86fF
C11737 a_1929_12131# VDD 4.53fF
C11738 a_44474_59182# a_45478_59182# 0.97fF
C11739 a_25306_22910# a_25398_22544# 0.32fF
C11740 a_38450_64202# VDD 0.51fF
C11741 a_15607_46805# a_26523_29199# 0.44fF
C11742 vcm_commonmode a_19282_14878# 0.31fF
C11743 ctopn a_16362_11500# 1.35fF
C11744 a_46482_56170# ctopp 3.40fF
C11745 a_12355_65103# a_16746_64204# 2.28fF
C11746 a_25398_14512# a_25398_13508# 1.00fF
C11747 a_13557_37999# VDD 1.79fF
C11748 ctopn a_40458_18528# 3.59fF
C11749 vcm_commonmode a_45386_64202# 0.31fF
C11750 a_1586_66567# a_1591_66415# 0.81fF
C11751 a_42466_17524# a_43470_17524# 0.97fF
C11752 a_13097_36367# a_31959_34751# 0.56fF
C11753 a_22843_29415# a_16863_29415# 1.66fF
C11754 vcm_commonmode a_16746_70228# 5.36fF
C11755 a_11067_13095# a_6607_42167# 1.92fF
C11756 a_29414_60186# a_30418_60186# 0.97fF
C11757 a_17366_23548# VDD 0.58fF
C11758 vcm_commonmode a_77451_38925# 140.35fF
C11759 a_46482_24552# a_46482_23548# 1.00fF
C11760 a_31422_12504# a_31422_11500# 1.00fF
C11761 a_32319_31599# VDD 0.50fF
C11762 a_4351_67279# a_7050_53333# 0.70fF
C11763 a_12889_40977# a_13909_41923# 0.34fF
C11764 vcm_commonmode a_24302_23914# 0.31fF
C11765 a_23507_44265# VDD 0.61fF
C11766 a_18370_70226# a_18370_69222# 1.00fF
C11767 vcm_commonmode a_21290_66210# 0.31fF
C11768 a_28756_55394# a_12983_63151# 0.40fF
C11769 a_24394_18528# a_25398_18528# 0.97fF
C11770 a_26402_19532# VDD 0.51fF
C11771 a_9353_72399# a_9707_73807# 0.39fF
C11772 a_9424_60949# VDD 0.69fF
C11773 a_37919_28111# VDD 6.39fF
C11774 a_45478_61190# ctopp 3.59fF
C11775 a_16510_8760# a_12877_16911# 1.07fF
C11776 a_47486_69222# VDD 0.51fF
C11777 a_1923_59583# a_1952_60431# 0.34fF
C11778 a_12663_35431# VDD 9.20fF
C11779 vcm_commonmode a_33338_19898# 0.31fF
C11780 a_17366_67214# ctopp 3.43fF
C11781 a_34251_52263# a_35438_55166# 0.46fF
C11782 a_8583_33551# a_8461_32937# 0.97fF
C11783 a_18151_52263# a_24394_63198# 0.42fF
C11784 a_25971_52263# a_12981_62313# 0.40fF
C11785 a_9779_47919# VDD 0.41fF
C11786 a_37919_28111# a_38450_13508# 0.38fF
C11787 a_16362_19532# a_16746_19530# 2.28fF
C11788 a_6559_22671# a_4798_23759# 0.33fF
C11789 vcm_commonmode a_34434_8488# 0.86fF
C11790 a_6467_55527# a_2952_53333# 0.34fF
C11791 a_45478_65206# VDD 0.51fF
C11792 a_26433_39631# a_13669_38517# 0.39fF
C11793 a_17366_11500# a_17366_10496# 1.00fF
C11794 a_21290_14878# a_21382_14512# 0.32fF
C11795 a_14646_29423# a_13390_29575# 0.89fF
C11796 a_37354_69222# a_37446_69222# 0.32fF
C11797 a_43470_18528# a_43470_17524# 1.00fF
C11798 a_11877_50645# VDD 0.65fF
C11799 a_23395_52047# a_27406_72234# 0.34fF
C11800 a_16362_55166# a_17366_55166# 0.97fF
C11801 a_34342_24918# VDD 0.36fF
C11802 a_47394_64202# a_47486_64202# 0.32fF
C11803 a_11067_67279# a_11067_21583# 0.63fF
C11804 ctopn a_44474_15516# 3.59fF
C11805 vcm_commonmode a_22386_67214# 0.87fF
C11806 a_28547_51175# a_12727_67753# 0.40fF
C11807 a_29414_20536# VDD 0.51fF
C11808 a_44382_55166# VDD 0.35fF
C11809 a_44382_22910# a_44474_22544# 0.32fF
C11810 a_18370_63198# VDD 0.57fF
C11811 a_33430_10496# a_34434_10496# 0.97fF
C11812 a_5073_27247# VDD 0.52fF
C11813 a_43175_28335# a_46482_24552# 0.55fF
C11814 a_35346_65206# a_35438_65206# 0.32fF
C11815 a_44474_14512# a_44474_13508# 1.00fF
C11816 vcm_commonmode a_36350_20902# 0.31fF
C11817 vcm_commonmode a_25306_63198# 0.31fF
C11818 a_1586_45431# a_7000_43541# 0.95fF
C11819 a_8199_58229# VDD 1.98fF
C11820 a_48490_60186# a_49494_60186# 0.97fF
C11821 vcm_commonmode a_19374_9492# 0.87fF
C11822 a_35601_27497# a_35438_21540# 0.38fF
C11823 a_26310_23914# a_26402_23548# 0.32fF
C11824 a_18979_30287# a_4811_34855# 0.98fF
C11825 a_19374_11500# a_20378_11500# 0.97fF
C11826 a_16228_28335# VDD 1.92fF
C11827 vcm_commonmode a_35438_16520# 0.87fF
C11828 a_16746_64204# ctopp 1.68fF
C11829 ctopn a_21382_13508# 3.59fF
C11830 a_21371_52263# VDD 14.11fF
C11831 vcm_commonmode a_19282_59182# 0.31fF
C11832 a_23298_66210# a_23390_66210# 0.32fF
C11833 a_29414_12504# VDD 0.51fF
C11834 a_37446_70226# a_37446_69222# 1.00fF
C11835 a_13183_52047# a_17366_66210# 0.38fF
C11836 a_3325_69135# a_3693_68047# 0.31fF
C11837 a_43470_18528# a_44474_18528# 0.97fF
C11838 a_12473_37429# a_12621_36091# 0.90fF
C11839 a_5915_35943# a_16510_8760# 0.45fF
C11840 a_21267_52047# VDD 0.82fF
C11841 vcm_commonmode a_31768_55394# 10.01fF
C11842 a_2899_27023# VDD 0.41fF
C11843 a_12481_54447# VDD 0.49fF
C11844 a_47486_55166# m3_47388_55078# 2.81fF
C11845 vcm_commonmode a_36350_12870# 0.31fF
C11846 a_2840_66103# a_28881_52271# 0.53fF
C11847 a_23390_24552# a_24394_24552# 0.97fF
C11848 a_23507_35561# VDD 0.60fF
C11849 a_12549_44212# a_12663_40871# 0.31fF
C11850 a_34780_56398# a_12901_66959# 0.40fF
C11851 a_40491_27247# a_43470_13508# 0.38fF
C11852 a_35346_19898# a_35438_19532# 0.32fF
C11853 a_24394_21540# VDD 0.51fF
C11854 vcm_commonmode a_27406_7484# 0.69fF
C11855 a_18979_30287# a_27890_32459# 0.40fF
C11856 a_20378_62194# a_21382_62194# 0.97fF
C11857 a_36442_11500# a_36442_10496# 1.00fF
C11858 a_40366_14878# a_40458_14512# 0.32fF
C11859 vcm_commonmode a_31330_21906# 0.31fF
C11860 a_25398_69222# ctopp 3.59fF
C11861 ctopn a_12899_10927# 3.23fF
C11862 a_32611_41317# VDD 0.87fF
C11863 vcm_commonmode a_21382_64202# 0.87fF
C11864 vcm_commonmode a_49402_58178# 0.30fF
C11865 a_29414_17524# VDD 0.51fF
C11866 a_41427_52263# a_41261_28335# 3.30fF
C11867 a_1591_64239# a_1591_57711# 0.32fF
C11868 a_19282_20902# a_19374_20536# 0.32fF
C11869 a_1768_16367# config_2_in[1] 0.76fF
C11870 a_12727_58255# VDD 7.18fF
C11871 a_4339_64521# a_7217_53047# 0.72fF
C11872 a_38239_32375# VDD 0.51fF
C11873 vcm_commonmode a_36350_17890# 0.31fF
C11874 a_23390_65206# ctopp 3.59fF
C11875 a_11803_55311# a_4215_51157# 0.53fF
C11876 a_1761_43567# a_19629_39631# 1.44fF
C11877 a_25398_57174# a_26402_57174# 0.97fF
C11878 vcm_commonmode a_23298_60186# 0.31fF
C11879 a_28410_15516# a_29414_15516# 0.97fF
C11880 a_6467_55527# a_3295_54421# 1.22fF
C11881 a_1761_40847# config_2_in[7] 1.12fF
C11882 a_12447_29199# a_8273_42479# 0.30fF
C11883 a_2689_65103# a_6095_44807# 0.33fF
C11884 a_17682_50095# a_24959_30503# 0.53fF
C11885 a_1586_45431# a_7553_48469# 0.61fF
C11886 vcm_commonmode a_30418_69222# 0.87fF
C11887 a_26402_71230# a_27406_71230# 0.97fF
C11888 a_12341_3311# a_22386_21540# 0.38fF
C11889 a_45386_23914# a_45478_23548# 0.32fF
C11890 a_38450_11500# a_39454_11500# 0.97fF
C11891 a_38557_32143# a_11067_46823# 0.53fF
C11892 a_3949_41935# a_5363_30503# 0.38fF
C11893 a_42374_66210# a_42466_66210# 0.32fF
C11894 vcm_commonmode a_37446_22544# 0.87fF
C11895 a_8491_41383# a_20267_30503# 0.60fF
C11896 a_13576_42589# VDD 3.21fF
C11897 vcm_commonmode a_28410_65206# 0.87fF
C11898 a_38557_32143# a_12355_65103# 0.40fF
C11899 a_1586_18695# a_8289_14741# 0.33fF
C11900 a_2216_28309# a_1915_35015# 2.94fF
C11901 a_13576_37149# a_1761_31055# 4.44fF
C11902 a_30418_18528# VDD 0.51fF
C11903 a_18278_72234# a_18370_72234# 0.32fF
C11904 a_12985_7663# a_16746_20534# 0.41fF
C11905 a_1761_39215# a_33155_35839# 0.51fF
C11906 ctopn a_28410_8488# 3.40fF
C11907 a_39673_28111# a_12546_22351# 0.41fF
C11908 a_42466_24552# a_43470_24552# 0.97fF
C11909 a_19282_12870# a_19374_12504# 0.32fF
C11910 a_26267_34473# VDD 0.56fF
C11911 vcm_commonmode a_37354_18894# 0.31fF
C11912 a_30418_66210# ctopp 3.59fF
C11913 a_23395_52047# a_19576_51701# 2.29fF
C11914 a_7841_12167# a_1586_18695# 0.59fF
C11915 a_12357_37999# a_24893_37429# 1.97fF
C11916 vcm_commonmode a_17274_24918# 0.31fF
C11917 a_10515_32143# a_11711_32143# 0.48fF
C11918 a_4191_33449# a_2787_32679# 0.62fF
C11919 a_14287_51175# a_4811_34855# 0.46fF
C11920 a_3339_43023# a_1803_19087# 8.09fF
C11921 a_21382_55166# VDD 0.60fF
C11922 a_41967_31375# a_12877_14441# 0.41fF
C11923 a_39454_62194# a_40458_62194# 0.97fF
C11924 vcm_commonmode a_33430_14512# 0.87fF
C11925 a_28756_7638# a_28410_24552# 0.47fF
C11926 a_4578_40455# a_3305_38671# 0.66fF
C11927 a_39468_37479# VDD 1.90fF
C11928 vcm_commonmode a_28318_55166# 0.30fF
C11929 a_39454_10496# VDD 0.51fF
C11930 a_4351_67279# a_2840_66103# 2.39fF
C11931 a_2191_68565# a_1823_65853# 0.98fF
C11932 a_37919_28111# a_38450_7484# 0.34fF
C11933 vcm_commonmode a_19282_57174# 0.31fF
C11934 a_2595_47653# a_7387_48469# 0.60fF
C11935 a_25971_52263# a_30418_71230# 0.38fF
C11936 a_38358_20902# a_38450_20536# 0.32fF
C11937 a_3295_54421# a_1823_58773# 1.12fF
C11938 vcm_commonmode a_46390_10862# 0.31fF
C11939 a_27314_63198# a_27406_63198# 0.32fF
C11940 a_5179_10927# a_5345_10927# 0.72fF
C11941 a_18370_57174# a_18370_56170# 1.00fF
C11942 a_44474_57174# a_45478_57174# 0.97fF
C11943 a_41427_52263# a_41462_61190# 0.38fF
C11944 a_10975_66407# a_16362_66210# 19.89fF
C11945 a_47486_15516# a_48490_15516# 0.97fF
C11946 vcm_commonmode a_38450_23548# 0.87fF
C11947 a_7571_29199# a_3339_32463# 0.78fF
C11948 a_29760_55394# a_29414_67214# 0.38fF
C11949 vcm_commonmode a_35438_66210# 0.87fF
C11950 a_12473_37429# a_12473_36341# 1.95fF
C11951 a_8295_47388# a_4443_46607# 0.59fF
C11952 a_25744_7638# a_12877_16911# 0.41fF
C11953 a_35601_27497# a_12899_11471# 0.41fF
C11954 a_26402_62194# VDD 0.51fF
C11955 a_2411_26133# a_1683_33237# 0.34fF
C11956 a_7571_29199# a_7841_29673# 0.38fF
C11957 a_30418_55166# m3_30320_55078# 2.81fF
C11958 a_1923_54591# a_2163_56765# 0.76fF
C11959 a_2748_68565# VDD 0.33fF
C11960 vcm_commonmode a_47486_19532# 0.87fF
C11961 ctopn a_29414_16520# 3.59fF
C11962 a_4674_40277# a_4314_40821# 0.42fF
C11963 vcm_commonmode a_33338_62194# 0.31fF
C11964 a_11067_13095# a_6883_37019# 0.39fF
C11965 a_34434_15516# VDD 0.51fF
C11966 a_1923_73087# a_1959_68053# 0.34fF
C11967 a_45478_71230# a_46482_71230# 0.97fF
C11968 a_21290_59182# a_21382_59182# 0.32fF
C11969 a_11067_47695# a_17039_51157# 1.36fF
C11970 a_12166_21501# VDD 0.50fF
C11971 a_11067_13095# a_5039_42167# 0.65fF
C11972 a_40675_27791# a_12895_13967# 0.41fF
C11973 a_1823_76181# a_6098_73095# 0.32fF
C11974 vcm_commonmode a_41370_15882# 0.31fF
C11975 a_34434_63198# ctopp 3.64fF
C11976 a_32426_71230# VDD 0.58fF
C11977 config_2_in[2] config_2_in[1] 0.77fF
C11978 a_33764_38567# VDD 1.79fF
C11979 a_10506_29967# a_6459_30511# 0.87fF
C11980 a_31422_72234# m3_31324_72146# 2.80fF
C11981 a_44474_11500# VDD 0.51fF
C11982 a_35932_41953# VDD 1.36fF
C11983 a_19282_17890# a_19374_17524# 0.32fF
C11984 vcm_commonmode a_39362_71230# 0.31fF
C11985 a_4298_58951# a_6795_51157# 1.52fF
C11986 a_33864_28111# a_12877_14441# 0.41fF
C11987 a_28410_59182# ctopp 3.59fF
C11988 a_25398_64202# a_25398_63198# 1.23fF
C11989 a_38358_12870# a_38450_12504# 0.32fF
C11990 a_9484_11989# a_9642_10357# 0.58fF
C11991 a_10515_22671# a_7862_34025# 1.02fF
C11992 a_9529_28335# a_17278_28309# 0.41fF
C11993 a_13067_38517# a_12473_41781# 2.03fF
C11994 a_38557_32143# ctopp 2.62fF
C11995 a_27417_32509# a_28430_32143# 0.35fF
C11996 a_33430_59182# a_33430_58178# 1.00fF
C11997 a_12251_39069# a_12381_35836# 0.47fF
C11998 a_10515_63143# a_11067_46823# 0.52fF
C11999 a_17366_22544# a_17366_21540# 1.00fF
C12000 a_36797_27497# a_12899_10927# 0.41fF
C12001 vcm_commonmode a_18278_13874# 0.31fF
C12002 a_1775_67503# VDD 0.73fF
C12003 a_24394_13508# a_25398_13508# 0.97fF
C12004 a_4495_35925# VDD 4.16fF
C12005 a_10975_66407# a_9179_22351# 0.45fF
C12006 vcm_commonmode a_39454_63198# 0.92fF
C12007 a_29414_68218# a_30418_68218# 0.97fF
C12008 a_40491_27247# a_43470_7484# 0.34fF
C12009 a_46482_72234# a_46482_71230# 1.00fF
C12010 a_1923_73087# a_9319_69141# 0.32fF
C12011 config_2_in[11] config_2_in[9] 0.41fF
C12012 a_1823_53885# a_2327_54135# 0.36fF
C12013 a_34482_29941# a_38239_32375# 0.34fF
C12014 a_41462_56170# a_41462_55166# 1.00fF
C12015 a_46390_63198# a_46482_63198# 0.32fF
C12016 a_6607_42167# a_4314_40821# 0.91fF
C12017 a_37446_57174# a_37446_56170# 1.00fF
C12018 vcm_commonmode a_33430_59182# 0.87fF
C12019 a_2606_41079# a_2004_42453# 0.80fF
C12020 a_41427_52263# a_33694_30761# 0.54fF
C12021 vcm_commonmode a_41967_31375# 10.41fF
C12022 a_1591_51183# VDD 0.41fF
C12023 a_11067_13095# a_3987_19623# 0.52fF
C12024 a_33338_21906# a_33430_21540# 0.32fF
C12025 a_42709_29199# a_12877_14441# 0.40fF
C12026 a_12447_29199# a_12263_4391# 0.39fF
C12027 a_1761_39215# a_12381_35836# 3.19fF
C12028 a_32426_60186# ctopp 3.59fF
C12029 a_26748_7638# a_26402_22544# 0.38fF
C12030 a_35438_68218# VDD 0.51fF
C12031 a_2840_66103# a_12755_53030# 1.49fF
C12032 a_35346_7850# VDD 0.61fF
C12033 a_21382_16520# a_21382_15516# 1.00fF
C12034 ctopn a_31422_22544# 3.58fF
C12035 vcm_commonmode a_42374_68218# 0.31fF
C12036 a_40366_59182# a_40458_59182# 0.32fF
C12037 a_6835_46823# a_4191_33449# 1.10fF
C12038 a_2689_65103# VDD 3.37fF
C12039 a_13123_38231# VDD 5.81fF
C12040 a_11067_67279# a_9135_27239# 0.42fF
C12041 vcm_commonmode a_45478_21540# 0.87fF
C12042 a_38358_17890# a_38450_17524# 0.32fF
C12043 a_30764_7638# a_30418_8488# 0.38fF
C12044 a_9503_26151# a_12877_14441# 0.41fF
C12045 a_28547_51175# a_7841_12167# 6.08fF
C12046 a_25306_60186# a_25398_60186# 0.32fF
C12047 a_9223_22895# VDD 0.41fF
C12048 vcm_commonmode a_22386_10496# 0.87fF
C12049 a_11067_13095# a_12899_10927# 1.46fF
C12050 a_24740_7638# a_24394_21540# 0.38fF
C12051 a_7803_55509# VDD 3.52fF
C12052 a_44474_64202# a_44474_63198# 1.23fF
C12053 ctopn a_27406_14512# 3.59fF
C12054 a_2235_41941# a_2401_41941# 0.66fF
C12055 vcm_commonmode a_37446_60186# 0.87fF
C12056 a_41261_28335# a_12981_59343# 0.40fF
C12057 a_49494_13508# VDD 1.10fF
C12058 a_17507_52047# a_12983_63151# 0.40fF
C12059 a_20286_18894# a_20378_18528# 0.32fF
C12060 a_36442_22544# a_36442_21540# 1.00fF
C12061 a_31768_7638# a_31422_16520# 0.38fF
C12062 a_3339_43023# a_1761_50639# 2.56fF
C12063 a_17691_27791# VDD 0.32fF
C12064 a_35438_56170# VDD 0.52fF
C12065 a_39223_32463# a_12985_19087# 0.41fF
C12066 a_43470_13508# a_44474_13508# 0.97fF
C12067 a_26523_29199# a_28841_29575# 1.10fF
C12068 a_18370_8488# VDD 0.58fF
C12069 a_18611_52047# a_12981_62313# 0.40fF
C12070 a_48490_68218# a_49494_68218# 0.97fF
C12071 a_16955_52047# a_20378_63198# 0.42fF
C12072 vcm_commonmode a_33864_28111# 10.30fF
C12073 vcm_commonmode a_42374_56170# 0.31fF
C12074 ctopn a_32426_23548# 3.46fF
C12075 a_3019_13621# VDD 1.02fF
C12076 vcm_commonmode a_25306_8854# 0.31fF
C12077 a_23736_7638# a_12985_16367# 0.41fF
C12078 a_4674_40277# a_6243_30662# 0.40fF
C12079 vcm_commonmode a_17366_15516# 1.82fF
C12080 a_28410_57174# ctopp 3.58fF
C12081 a_29414_56170# a_30418_56170# 0.97fF
C12082 a_16362_14512# a_16746_14510# 2.28fF
C12083 ctopn a_41462_19532# 3.59fF
C12084 vcm_commonmode a_12907_56399# 5.77fF
C12085 a_34434_61190# VDD 0.51fF
C12086 vcm_commonmode a_27406_11500# 0.87fF
C12087 a_33430_58178# a_33430_57174# 1.00fF
C12088 a_49494_56170# m3_49396_56082# 2.78fF
C12089 a_2939_33535# VDD 0.41fF
C12090 a_11067_67279# a_12546_22351# 0.83fF
C12091 a_18611_52047# a_20535_51727# 0.34fF
C12092 vcm_commonmode a_41370_61190# 0.31fF
C12093 a_40458_16520# a_40458_15516# 1.00fF
C12094 vcm_commonmode a_31422_24552# 0.84fF
C12095 a_20635_29415# a_18979_30287# 0.57fF
C12096 a_21371_50959# a_12727_67753# 0.40fF
C12097 a_1591_18543# a_1757_18543# 0.43fF
C12098 a_25398_19532# a_25398_18528# 1.00fF
C12099 a_39223_32463# a_39454_14512# 0.38fF
C12100 a_6831_63303# VDD 13.11fF
C12101 a_29322_10862# a_29414_10496# 0.32fF
C12102 a_42466_62194# ctopp 3.59fF
C12103 a_38450_70226# VDD 0.51fF
C12104 a_7580_61751# a_7210_55081# 0.64fF
C12105 a_15253_37692# VDD 0.96fF
C12106 vcm_commonmode a_41462_55166# 0.84fF
C12107 a_36579_40183# VDD 0.66fF
C12108 vcm_commonmode a_16746_63200# 5.36fF
C12109 vcm_commonmode a_42709_29199# 10.28fF
C12110 vcm_commonmode a_33430_57174# 0.87fF
C12111 a_19374_16520# VDD 0.51fF
C12112 vcm_commonmode a_45386_70226# 0.31fF
C12113 a_5363_30503# a_5441_27791# 0.44fF
C12114 a_44382_60186# a_44474_60186# 0.32fF
C12115 VDD config_1_in[8] 1.12fF
C12116 a_12935_31287# VDD 2.30fF
C12117 vcm_commonmode a_26310_16886# 0.31fF
C12118 a_19720_55394# VDD 6.34fF
C12119 a_20378_15516# a_20378_14512# 1.00fF
C12120 a_48490_71230# ctopp 3.24fF
C12121 ctopn a_44474_20536# 3.59fF
C12122 a_43470_7484# m3_43372_7346# 2.80fF
C12123 a_39362_18894# a_39454_18528# 0.32fF
C12124 a_25517_37455# a_1761_30511# 0.96fF
C12125 vcm_commonmode a_18151_52263# 10.02fF
C12126 a_6327_72917# a_7925_72399# 0.35fF
C12127 a_6831_63303# a_26514_47375# 0.82fF
C12128 a_28410_61190# a_29414_61190# 0.97fF
C12129 a_40458_55166# m3_40360_55078# 2.81fF
C12130 a_4516_55107# VDD 0.64fF
C12131 a_19282_24918# a_19374_24552# 0.32fF
C12132 a_11999_67477# VDD 0.84fF
C12133 a_1803_20719# a_13835_43177# 1.57fF
C12134 a_34434_68218# a_34434_67214# 1.00fF
C12135 vcm_commonmode a_47486_62194# 0.87fF
C12136 vcm_commonmode a_9503_26151# 10.36fF
C12137 a_20635_29415# a_37427_47893# 1.09fF
C12138 vcm_commonmode a_18370_68218# 0.88fF
C12139 a_23395_52047# a_12901_66959# 0.40fF
C12140 a_27406_58178# VDD 0.51fF
C12141 a_10665_20969# VDD 0.78fF
C12142 a_3247_20495# a_2235_30503# 0.36fF
C12143 a_29927_29199# a_32970_31145# 0.42fF
C12144 ctopn a_44474_12504# 3.59fF
C12145 a_36613_48169# a_12907_27023# 0.55fF
C12146 a_16510_8760# a_12895_13967# 1.08fF
C12147 a_48490_56170# a_49494_56170# 0.97fF
C12148 vcm_commonmode a_34342_58178# 0.31fF
C12149 a_75794_38962# VDD 0.73fF
C12150 a_16746_69224# ctopp 1.68fF
C12151 a_18811_41317# VDD 0.92fF
C12152 a_19374_69222# a_19374_68218# 1.00fF
C12153 VDD dummypin[8] 0.87fF
C12154 a_9135_27239# a_21382_8488# 0.38fF
C12155 a_37446_72234# a_38450_72234# 0.97fF
C12156 a_17712_7638# a_12727_15529# 0.40fF
C12157 a_4674_40277# a_5085_23047# 0.55fF
C12158 a_31422_8488# a_32426_8488# 0.97fF
C12159 a_30326_55166# a_30418_55166# 0.32fF
C12160 a_44474_67214# VDD 0.51fF
C12161 a_15439_49525# a_8123_56399# 1.11fF
C12162 a_21290_57174# a_21382_57174# 0.32fF
C12163 a_9011_74879# VDD 0.61fF
C12164 a_24302_15882# a_24394_15516# 0.32fF
C12165 ctopn a_39454_21540# 3.59fF
C12166 a_28757_27247# a_30788_28487# 0.36fF
C12167 a_17863_44211# VDD 1.46fF
C12168 a_32426_70226# a_33430_70226# 0.97fF
C12169 a_44474_19532# a_44474_18528# 1.00fF
C12170 a_37919_28111# a_38450_11500# 0.38fF
C12171 a_2021_22325# a_4798_23759# 0.48fF
C12172 VDD dummypin[7] 0.81fF
C12173 a_8575_74853# a_10055_74031# 0.36fF
C12174 a_32951_27247# a_33430_18528# 0.38fF
C12175 a_30023_41959# a_12381_35836# 0.70fF
C12176 a_48398_10862# a_48490_10496# 0.32fF
C12177 a_41159_28585# VDD 0.42fF
C12178 vcm_commonmode a_32426_13508# 0.87fF
C12179 ctopn a_16362_10496# 1.35fF
C12180 a_10747_68565# VDD 0.80fF
C12181 a_27600_36165# VDD 1.78fF
C12182 ctopn a_44474_17524# 3.59fF
C12183 a_41462_9492# VDD 0.51fF
C12184 a_2021_22325# a_2021_17973# 0.47fF
C12185 a_5024_67885# a_5254_67503# 0.70fF
C12186 a_1591_57711# a_2099_64757# 0.86fF
C12187 vcm_commonmode a_18370_56170# 0.88fF
C12188 a_17039_51157# a_18539_47617# 0.31fF
C12189 a_9989_46831# a_7000_43541# 1.10fF
C12190 a_22294_71230# a_22386_71230# 0.32fF
C12191 vcm_commonmode a_21290_69222# 0.31fF
C12192 a_10515_22671# a_5039_42167# 0.99fF
C12193 a_30418_60186# a_30418_59182# 1.00fF
C12194 a_2163_59585# a_2124_59459# 0.72fF
C12195 a_21382_22544# VDD 0.51fF
C12196 vcm_commonmode a_48398_9858# 0.31fF
C12197 a_9735_63669# VDD 0.98fF
C12198 a_19374_63198# a_19374_62194# 1.00fF
C12199 a_34342_11866# a_34434_11500# 0.32fF
C12200 a_12999_29423# VDD 0.60fF
C12201 a_47486_72234# VDD 1.23fF
C12202 a_39454_15516# a_39454_14512# 1.00fF
C12203 vcm_commonmode a_28318_22910# 0.31fF
C12204 a_16746_70228# ctopp 1.65fF
C12205 a_11067_23759# a_12263_4391# 6.05fF
C12206 a_2411_26133# VDD 10.49fF
C12207 vcm_commonmode a_19282_65206# 0.31fF
C12208 a_31768_55394# a_12355_65103# 0.40fF
C12209 a_2411_18517# a_5363_16367# 0.55fF
C12210 a_1761_30511# a_12713_36483# 0.82fF
C12211 a_12993_50345# VDD 1.33fF
C12212 a_11141_60975# VDD 0.61fF
C12213 a_47486_61190# a_48490_61190# 0.97fF
C12214 a_24394_9492# a_24394_8488# 1.00fF
C12215 a_12082_25077# VDD 0.31fF
C12216 a_38358_24918# a_38450_24552# 0.32fF
C12217 a_1768_13103# a_1591_59343# 0.58fF
C12218 a_12249_43457# a_12641_43124# 0.41fF
C12219 a_49494_7484# VDD 2.17fF
C12220 a_19374_67214# a_20378_67214# 0.97fF
C12221 vcm_commonmode a_17366_61190# 1.83fF
C12222 a_17366_14512# VDD 0.57fF
C12223 a_6467_55527# a_35568_49525# 0.31fF
C12224 a_43470_64202# VDD 0.51fF
C12225 a_35346_62194# a_35438_62194# 0.32fF
C12226 vcm_commonmode a_24302_14878# 0.31fF
C12227 ctopn a_21382_11500# 3.59fF
C12228 a_19743_38007# VDD 0.61fF
C12229 a_11067_67279# a_32951_27247# 0.41fF
C12230 ctopn a_45478_18528# 3.59fF
C12231 a_2539_42106# a_1761_22895# 0.35fF
C12232 a_75628_40594# VDD 0.32fF
C12233 a_38450_69222# a_38450_68218# 1.00fF
C12234 a_5915_30287# a_2787_30503# 0.91fF
C12235 vcm_commonmode a_21382_70226# 0.87fF
C12236 a_21371_52263# a_26402_71230# 0.38fF
C12237 a_38450_58178# vcm_commonmode 0.87fF
C12238 a_28410_8488# a_28410_7484# 1.00fF
C12239 a_49402_55166# a_49494_55166# 0.32fF
C12240 a_22386_23548# VDD 0.52fF
C12241 a_19374_66210# VDD 0.51fF
C12242 a_2223_28617# a_3325_18543# 0.36fF
C12243 a_13716_43047# a_32121_40741# 0.42fF
C12244 a_40366_57174# a_40458_57174# 0.32fF
C12245 a_2843_71829# VDD 3.87fF
C12246 a_36613_48169# a_37446_61190# 0.38fF
C12247 a_12727_15529# a_16362_14512# 1.27fF
C12248 a_43378_15882# a_43470_15516# 0.32fF
C12249 vcm_commonmode a_29322_23914# 0.31fF
C12250 a_21371_50959# a_25398_67214# 0.38fF
C12251 vcm_commonmode a_26310_66210# 0.31fF
C12252 a_40491_27247# a_43470_11500# 0.38fF
C12253 ctopn a_31768_7638# 2.63fF
C12254 a_21382_58178# a_22386_58178# 0.97fF
C12255 a_31422_19532# VDD 0.51fF
C12256 a_4792_52539# VDD 0.62fF
C12257 a_23390_55166# m3_23292_55078# 2.81fF
C12258 a_17366_13508# a_17366_12504# 1.00fF
C12259 vcm_commonmode a_38358_19898# 0.31fF
C12260 a_22386_67214# ctopp 3.59fF
C12261 a_32426_16520# a_33430_16520# 0.97fF
C12262 a_41370_71230# a_41462_71230# 0.32fF
C12263 a_13183_52047# a_17366_69222# 0.38fF
C12264 a_39673_28111# a_40458_13508# 0.38fF
C12265 a_16746_59184# a_16362_59182# 2.28fF
C12266 a_49494_60186# a_49494_59182# 1.00fF
C12267 vcm_commonmode a_39454_8488# 0.86fF
C12268 m3_30320_7346# VDD 0.33fF
C12269 a_38450_63198# a_38450_62194# 1.00fF
C12270 a_6752_29941# VDD 1.07fF
C12271 a_19780_39429# VDD 1.80fF
C12272 a_11067_67279# a_43175_28335# 0.41fF
C12273 ctopn a_30764_7638# 2.62fF
C12274 a_14681_50247# VDD 0.39fF
C12275 a_1586_40455# config_2_in[12] 0.33fF
C12276 a_43470_9492# a_43470_8488# 1.00fF
C12277 a_39362_24918# VDD 0.36fF
C12278 a_19807_28111# a_7862_34025# 0.31fF
C12279 a_38450_67214# a_39454_67214# 0.97fF
C12280 a_31768_55394# ctopp 2.63fF
C12281 a_3417_33231# a_3417_31599# 0.32fF
C12282 vcm_commonmode a_27406_67214# 0.87fF
C12283 a_34434_20536# VDD 0.51fF
C12284 a_23390_63198# VDD 0.57fF
C12285 a_17278_28309# VDD 0.58fF
C12286 a_34780_56398# a_34434_58178# 0.38fF
C12287 a_20286_13874# a_20378_13508# 0.32fF
C12288 vcm_commonmode a_41370_20902# 0.31fF
C12289 a_1761_22895# a_2021_22325# 7.85fF
C12290 a_25306_68218# a_25398_68218# 0.32fF
C12291 vcm_commonmode a_30326_63198# 0.31fF
C12292 a_42466_72234# a_42466_71230# 1.00fF
C12293 a_17366_59182# VDD 0.58fF
C12294 a_47486_8488# a_47486_7484# 1.00fF
C12295 a_24394_7484# a_25398_7484# 0.97fF
C12296 vcm_commonmode a_24394_9492# 0.87fF
C12297 a_41967_31375# a_12899_11471# 0.41fF
C12298 a_2840_53511# a_5653_60039# 0.42fF
C12299 vcm_commonmode a_40458_16520# 0.87fF
C12300 a_21382_64202# ctopp 3.59fF
C12301 ctopn a_26402_13508# 3.59fF
C12302 vcm_commonmode a_24302_59182# 0.31fF
C12303 a_34434_12504# VDD 0.51fF
C12304 a_1761_37039# a_12549_35836# 2.29fF
C12305 a_2872_44111# a_11067_46823# 0.64fF
C12306 a_39673_28111# a_12985_16367# 0.41fF
C12307 a_35438_9492# a_36442_9492# 0.97fF
C12308 a_1591_26159# VDD 0.42fF
C12309 vcm_commonmode a_41370_12870# 0.31fF
C12310 a_18370_64202# a_19374_64202# 0.97fF
C12311 a_36442_13508# a_36442_12504# 1.00fF
C12312 a_31131_35281# VDD 0.43fF
C12313 a_12727_13353# a_12877_14441# 23.46fF
C12314 a_7387_48469# a_7553_48469# 0.58fF
C12315 a_29414_21540# VDD 0.51fF
C12316 vcm_commonmode a_32426_7484# 0.68fF
C12317 a_42718_27497# a_12985_19087# 0.41fF
C12318 a_25744_7638# a_12895_13967# 0.41fF
C12319 a_26748_7638# a_12899_10927# 0.41fF
C12320 a_47486_58178# VDD 0.51fF
C12321 a_7155_55509# a_4758_45369# 0.44fF
C12322 a_5024_67885# a_6417_62215# 0.72fF
C12323 a_22319_38825# VDD 0.64fF
C12324 a_11067_67279# a_43270_27791# 0.41fF
C12325 vcm_commonmode a_36350_21906# 0.31fF
C12326 a_30418_69222# ctopp 3.59fF
C12327 a_1591_40303# VDD 0.46fF
C12328 vcm_commonmode a_26402_64202# 0.87fF
C12329 a_6883_37019# a_6243_30662# 0.36fF
C12330 a_5915_35943# a_2787_30503# 0.35fF
C12331 a_34434_17524# VDD 0.51fF
C12332 a_43378_72234# a_43470_72234# 0.32fF
C12333 a_21382_60186# VDD 0.51fF
C12334 a_39223_32463# VDD 7.02fF
C12335 vcm_commonmode a_41370_17890# 0.31fF
C12336 a_28410_65206# ctopp 3.59fF
C12337 a_26402_67214# a_26402_66210# 1.00fF
C12338 vcm_commonmode a_28318_60186# 0.31fF
C12339 a_34251_52263# a_12981_59343# 0.40fF
C12340 vcm_commonmode a_12947_23413# 1.46fF
C12341 a_37706_44135# VDD 0.55fF
C12342 a_12516_7093# a_12901_66959# 24.02fF
C12343 a_11303_53511# VDD 0.45fF
C12344 a_10055_74031# a_10221_74031# 0.69fF
C12345 a_33864_28111# a_12899_11471# 0.41fF
C12346 a_36629_27791# a_12877_16911# 0.41fF
C12347 a_5671_21495# a_7377_18012# 0.34fF
C12348 a_1823_62589# VDD 1.51fF
C12349 a_22386_65206# a_22386_64202# 1.00fF
C12350 a_39362_13874# a_39454_13508# 0.32fF
C12351 a_24800_43041# a_12549_44212# 0.44fF
C12352 a_44382_68218# a_44474_68218# 0.32fF
C12353 a_2606_41079# a_17488_48731# 0.60fF
C12354 a_30125_47919# VDD 0.48fF
C12355 vcm_commonmode a_35438_69222# 0.87fF
C12356 a_2099_59861# a_2467_47893# 0.40fF
C12357 a_43470_7484# a_44474_7484# 0.97fF
C12358 a_6162_28487# a_8373_26409# 0.51fF
C12359 a_25306_56170# a_25398_56170# 0.32fF
C12360 vcm_commonmode a_42466_22544# 0.87fF
C12361 a_10506_29967# a_14625_30761# 0.36fF
C12362 a_2606_41079# a_1761_41935# 0.82fF
C12363 a_10661_10383# VDD 0.35fF
C12364 vcm_commonmode a_33430_65206# 0.87fF
C12365 a_27406_69222# a_28410_69222# 0.97fF
C12366 a_1591_57711# a_1915_67477# 0.70fF
C12367 a_17039_51157# a_2606_41079# 0.37fF
C12368 a_35438_18528# VDD 0.51fF
C12369 a_16955_52047# a_20378_72234# 0.34fF
C12370 a_18979_30287# a_12899_2767# 0.70fF
C12371 a_22386_61190# a_22386_60186# 1.00fF
C12372 a_11865_24527# VDD 0.74fF
C12373 vcm_commonmode a_18278_11866# 0.31fF
C12374 a_11251_59879# a_3339_43023# 1.24fF
C12375 ctopn a_33430_8488# 3.40fF
C12376 a_42718_27497# a_44474_23548# 0.38fF
C12377 a_1954_61677# VDD 3.08fF
C12378 a_37446_64202# a_38450_64202# 0.97fF
C12379 vcm_commonmode a_42374_18894# 0.31fF
C12380 a_35438_66210# ctopp 3.59fF
C12381 a_21371_52263# a_25419_50959# 0.97fF
C12382 a_1689_10396# a_2339_38129# 1.15fF
C12383 vcm_commonmode a_22294_24918# 0.31fF
C12384 a_6655_46261# VDD 0.54fF
C12385 a_12516_7093# a_16362_70226# 19.89fF
C12386 a_14287_51175# a_12727_67753# 0.40fF
C12387 a_7749_37903# a_5915_35943# 0.40fF
C12388 a_3325_49551# a_1761_50639# 0.59fF
C12389 a_26402_55166# VDD 0.60fF
C12390 a_42709_29199# a_12899_11471# 0.40fF
C12391 a_34434_22544# a_35438_22544# 0.97fF
C12392 a_12889_39889# a_13669_38517# 0.58fF
C12393 a_4339_64521# a_8199_58229# 0.40fF
C12394 a_17366_57174# VDD 0.58fF
C12395 vcm_commonmode a_38450_14512# 0.87fF
C12396 a_7841_12167# a_7987_15431# 0.45fF
C12397 a_25398_65206# a_26402_65206# 0.97fF
C12398 vcm_commonmode a_17366_20536# 1.82fF
C12399 a_7155_55509# a_9695_54965# 0.35fF
C12400 a_44474_10496# VDD 0.51fF
C12401 a_21479_40229# VDD 0.91fF
C12402 a_21382_17524# a_21382_16520# 1.00fF
C12403 a_39673_28111# a_40458_7484# 0.35fF
C12404 vcm_commonmode a_24302_57174# 0.31fF
C12405 a_20359_29199# a_22015_28111# 1.09fF
C12406 a_7571_26151# a_9955_20969# 0.66fF
C12407 a_3247_20495# a_5073_27247# 0.42fF
C12408 a_35601_27497# a_12985_7663# 0.41fF
C12409 a_25398_56170# a_25398_55166# 1.00fF
C12410 a_32970_31145# VDD 2.18fF
C12411 vcm_commonmode a_12727_13353# 6.31fF
C12412 a_2004_42453# a_2339_38129# 1.08fF
C12413 a_4119_70741# VDD 6.58fF
C12414 a_45478_67214# a_45478_66210# 1.00fF
C12415 vcm_commonmode a_43470_23548# 0.87fF
C12416 a_36442_7484# m3_36344_7346# 2.80fF
C12417 vcm_commonmode a_40458_66210# 0.87fF
C12418 a_11067_63143# a_17488_48731# 5.87fF
C12419 a_9503_26151# a_12899_11471# 0.41fF
C12420 a_31422_62194# VDD 0.51fF
C12421 a_24302_61190# a_24394_61190# 0.32fF
C12422 vcm_commonmode a_17366_12504# 1.82fF
C12423 a_8491_57487# a_8123_56399# 0.56fF
C12424 ctopn a_18370_9492# 3.57fF
C12425 a_8531_70543# a_4482_57863# 4.05fF
C12426 a_41462_65206# a_41462_64202# 1.00fF
C12427 a_30311_35877# VDD 1.03fF
C12428 ctopn a_34434_16520# 3.59fF
C12429 a_1803_20719# a_1803_19087# 4.78fF
C12430 a_4443_46607# a_4941_35727# 1.24fF
C12431 vcm_commonmode a_38358_62194# 0.31fF
C12432 a_20359_29199# a_37557_32463# 0.72fF
C12433 a_39454_15516# VDD 0.51fF
C12434 a_16955_52047# a_12901_66959# 0.40fF
C12435 a_25744_7638# a_25398_13508# 0.38fF
C12436 a_25398_19532# a_26402_19532# 0.97fF
C12437 a_8491_27023# a_18370_13508# 0.38fF
C12438 a_35438_23548# a_35438_22544# 1.00fF
C12439 a_6375_64489# VDD 0.34fF
C12440 a_2012_33927# config_2_in[4] 0.58fF
C12441 vcm_commonmode a_46390_15882# 0.31fF
C12442 a_39454_63198# ctopp 3.64fF
C12443 a_1761_41935# a_12889_39889# 0.43fF
C12444 a_44382_56170# a_44474_56170# 0.32fF
C12445 a_37446_71230# VDD 0.58fF
C12446 a_29414_66210# a_29414_65206# 1.00fF
C12447 a_30418_14512# a_31422_14512# 0.97fF
C12448 a_34434_72234# m3_34336_72146# 2.80fF
C12449 a_49494_11500# VDD 1.25fF
C12450 a_5831_39189# a_1761_44111# 0.92fF
C12451 a_1761_46287# a_4500_45289# 0.33fF
C12452 a_12907_56399# a_12355_65103# 1.29fF
C12453 a_46482_69222# a_47486_69222# 0.97fF
C12454 a_1761_31055# a_1761_35407# 0.31fF
C12455 a_12549_35836# a_12663_35431# 0.54fF
C12456 a_6921_72943# a_7289_70767# 0.39fF
C12457 a_34780_56398# a_34251_52263# 0.32fF
C12458 vcm_commonmode a_44382_71230# 0.31fF
C12459 a_41462_61190# a_41462_60186# 1.00fF
C12460 a_27314_8854# a_27406_8488# 0.32fF
C12461 a_33430_59182# ctopp 3.59fF
C12462 a_16917_31573# VDD 0.59fF
C12463 vcm_commonmode a_17366_17524# 1.82fF
C12464 a_14471_28585# a_10873_27497# 0.61fF
C12465 a_16746_57176# a_16362_57174# 2.28fF
C12466 a_10975_66407# a_9367_29397# 1.14fF
C12467 vcm_commonmode a_10515_23975# 6.39fF
C12468 a_16362_13508# VDD 2.47fF
C12469 a_28318_70226# a_28410_70226# 0.32fF
C12470 a_1923_54591# a_4891_47388# 0.32fF
C12471 a_2451_72373# a_1923_73087# 0.98fF
C12472 a_7921_74581# a_6224_73095# 0.62fF
C12473 a_6095_44807# a_4674_40277# 0.50fF
C12474 a_27406_62194# a_27406_61190# 1.00fF
C12475 a_18370_10496# a_18370_9492# 1.00fF
C12476 vcm_commonmode a_23298_13874# 0.31fF
C12477 a_44474_65206# a_45478_65206# 0.97fF
C12478 a_11067_67279# a_12341_3311# 2.04fF
C12479 a_1895_30138# a_1757_29973# 0.46fF
C12480 vcm_commonmode a_44474_63198# 0.92fF
C12481 a_40458_17524# a_40458_16520# 1.00fF
C12482 a_13643_28327# a_16863_29415# 1.49fF
C12483 a_4149_48469# VDD 0.64fF
C12484 a_27406_20536# a_27406_19532# 1.00fF
C12485 a_10526_22057# VDD 1.17fF
C12486 a_35438_23548# a_36442_23548# 0.97fF
C12487 a_43269_29967# a_12899_10927# 0.41fF
C12488 a_9280_65327# VDD 0.48fF
C12489 a_18151_52263# a_11067_46823# 1.79fF
C12490 a_40458_72234# VDD 1.25fF
C12491 a_41872_29423# a_12727_58255# 0.40fF
C12492 a_32426_66210# a_33430_66210# 0.97fF
C12493 vcm_commonmode a_38450_59182# 0.87fF
C12494 a_1923_59583# a_7387_64239# 0.38fF
C12495 a_14926_31849# a_14361_29967# 0.39fF
C12496 vcm_commonmode m3_16264_57086# 3.20fF
C12497 a_32795_42943# VDD 0.92fF
C12498 a_18151_52263# a_12355_65103# 2.75fF
C12499 a_3339_43023# a_19919_38695# 0.40fF
C12500 a_7841_12167# a_13357_32143# 1.28fF
C12501 a_6795_51157# VDD 0.90fF
C12502 vcm_commonmode a_45478_72234# 0.69fF
C12503 a_10515_63143# a_7571_26151# 1.52fF
C12504 a_1586_51335# VDD 8.43fF
C12505 a_8273_42479# a_8117_30287# 0.35fF
C12506 a_43378_61190# a_43470_61190# 0.32fF
C12507 a_3578_25625# VDD 0.40fF
C12508 a_37446_60186# ctopp 3.59fF
C12509 a_40458_68218# VDD 0.51fF
C12510 vcm_commonmode a_18370_18528# 0.88fF
C12511 a_40366_7850# VDD 0.62fF
C12512 ctopn a_36442_22544# 3.58fF
C12513 vcm_commonmode a_47394_68218# 0.31fF
C12514 a_32426_71230# a_32426_70226# 1.00fF
C12515 a_5682_69367# a_3143_66972# 0.86fF
C12516 a_44474_19532# a_45478_19532# 0.97fF
C12517 a_6467_55527# a_27627_51733# 0.72fF
C12518 a_1761_39215# a_13484_39325# 1.79fF
C12519 a_48490_66210# a_48490_65206# 1.00fF
C12520 a_43267_31055# a_46482_59182# 0.38fF
C12521 a_10515_63143# a_9135_29423# 1.05fF
C12522 a_1591_49557# a_1757_49557# 0.72fF
C12523 a_17599_52263# a_22386_71230# 0.38fF
C12524 a_28410_20536# a_29414_20536# 0.97fF
C12525 a_46390_8854# a_46482_8488# 0.32fF
C12526 vcm_commonmode a_27406_10496# 0.87fF
C12527 a_17366_63198# a_18370_63198# 0.97fF
C12528 ctopn a_32426_14512# 3.59fF
C12529 a_25787_28327# a_33430_61190# 0.38fF
C12530 vcm_commonmode a_42466_60186# 0.87fF
C12531 a_33694_30761# a_36507_31573# 0.67fF
C12532 a_30788_28487# a_28446_31375# 0.80fF
C12533 a_16891_44265# VDD 0.64fF
C12534 vcm_commonmode a_16362_66210# 4.47fF
C12535 a_47394_70226# a_47486_70226# 0.32fF
C12536 a_17507_52047# a_21382_67214# 0.38fF
C12537 a_3339_43023# a_15009_40193# 0.40fF
C12538 a_17274_58178# a_17366_58178# 0.32fF
C12539 a_35568_49525# a_35676_49525# 0.84fF
C12540 a_9271_52789# VDD 0.54fF
C12541 a_6098_73095# a_6327_72917# 0.43fF
C12542 a_46482_62194# a_46482_61190# 1.00fF
C12543 a_37446_10496# a_37446_9492# 1.00fF
C12544 a_40458_56170# VDD 0.52fF
C12545 a_5254_67503# a_7210_55081# 0.64fF
C12546 a_35196_35425# VDD 1.54fF
C12547 a_23195_29967# a_23685_29111# 0.45fF
C12548 a_23390_8488# VDD 0.58fF
C12549 a_43362_28879# a_47486_64202# 0.38fF
C12550 a_28318_16886# a_28410_16520# 0.32fF
C12551 vcm_commonmode a_47394_56170# 0.31fF
C12552 a_1689_10396# a_1895_18756# 0.39fF
C12553 ctopn a_37446_23548# 3.40fF
C12554 a_20359_29199# a_22291_29415# 0.92fF
C12555 a_1761_52815# a_1803_20719# 0.30fF
C12556 a_20635_29415# a_18703_29199# 1.05fF
C12557 a_46482_20536# a_46482_19532# 1.00fF
C12558 a_42466_58178# a_41261_28335# 0.38fF
C12559 a_10055_58791# a_4482_57863# 0.54fF
C12560 vcm_commonmode a_30326_8854# 0.31fF
C12561 a_34482_29941# a_32970_31145# 1.29fF
C12562 vcm_commonmode a_22386_15516# 0.87fF
C12563 a_16746_63200# ctopp 1.68fF
C12564 a_33430_57174# ctopp 3.59fF
C12565 a_3983_70767# VDD 0.39fF
C12566 ctopn a_46482_19532# 3.59fF
C12567 vcm_commonmode a_20378_71230# 0.86fF
C12568 a_35601_27497# a_35438_16520# 0.38fF
C12569 a_26402_21540# a_26402_20536# 1.00fF
C12570 a_39454_61190# VDD 0.51fF
C12571 vcm_commonmode a_32426_11500# 0.87fF
C12572 a_41967_31375# a_42466_19532# 0.38fF
C12573 a_4983_66959# VDD 0.93fF
C12574 a_28410_12504# a_29414_12504# 0.97fF
C12575 vcm_commonmode a_46390_61190# 0.31fF
C12576 a_34342_67214# a_34434_67214# 0.32fF
C12577 vcm_commonmode a_36442_24552# 0.84fF
C12578 a_18151_52263# ctopp 2.62fF
C12579 a_19807_28111# a_20267_30503# 0.36fF
C12580 a_1591_45205# VDD 0.38fF
C12581 vcm_commonmode a_18278_67214# 0.31fF
C12582 a_2959_47113# a_29361_51727# 1.36fF
C12583 a_13669_39605# a_13909_38659# 0.57fF
C12584 a_21187_29415# a_28305_28879# 0.94fF
C12585 a_47486_62194# ctopp 3.58fF
C12586 a_77086_40693# a_76971_38925# 1.46fF
C12587 a_12659_54965# a_12755_53030# 1.03fF
C12588 a_43470_70226# VDD 0.51fF
C12589 a_25971_52263# a_30418_58178# 0.38fF
C12590 a_22521_37692# VDD 1.06fF
C12591 a_18370_68218# ctopp 3.58fF
C12592 vcm_commonmode a_46482_55166# 0.84fF
C12593 a_25744_7638# a_25398_7484# 0.34fF
C12594 a_8491_27023# a_18370_7484# 0.34fF
C12595 vcm_commonmode a_38450_57174# 0.87fF
C12596 a_24394_16520# VDD 0.51fF
C12597 a_38450_72234# a_38450_71230# 1.00fF
C12598 a_47486_20536# a_48490_20536# 0.97fF
C12599 a_20286_7850# a_20378_7484# 0.32fF
C12600 a_3247_20495# a_4495_35925# 1.10fF
C12601 a_32426_56170# a_32426_55166# 1.00fF
C12602 a_36442_63198# a_37446_63198# 0.97fF
C12603 vcm_commonmode a_31330_16886# 0.31fF
C12604 a_35099_43447# VDD 0.57fF
C12605 a_37919_28111# a_38450_10496# 0.38fF
C12606 a_36350_58178# a_36442_58178# 0.32fF
C12607 a_34699_37683# a_32971_35281# 0.32fF
C12608 a_15261_51433# VDD 0.39fF
C12609 a_23390_21540# a_24394_21540# 0.97fF
C12610 a_13643_28327# a_19720_7638# 0.64fF
C12611 a_31330_9858# a_31422_9492# 0.32fF
C12612 a_42718_27497# VDD 6.20fF
C12613 a_9123_55223# VDD 0.53fF
C12614 a_10472_26159# a_7841_22895# 0.39fF
C12615 a_16362_68218# VDD 2.48fF
C12616 a_21187_29415# a_4811_34855# 0.78fF
C12617 a_16362_7484# VDD 1.76fF
C12618 a_8583_33551# a_33694_30761# 0.52fF
C12619 a_7580_61751# a_7213_62215# 0.32fF
C12620 a_47394_16886# a_47486_16520# 0.32fF
C12621 a_43267_31055# a_46482_57174# 0.38fF
C12622 a_11803_55311# a_12257_56623# 1.07fF
C12623 a_7939_30503# a_2787_30503# 0.71fF
C12624 a_4674_40277# VDD 13.38fF
C12625 vcm_commonmode a_23390_68218# 0.87fF
C12626 a_32426_58178# VDD 0.51fF
C12627 a_30418_59182# a_31422_59182# 0.97fF
C12628 a_6831_63303# a_26397_51183# 0.79fF
C12629 a_4758_45369# a_19877_52245# 0.35fF
C12630 a_6467_55527# a_19576_51701# 1.10fF
C12631 a_7773_63927# VDD 3.08fF
C12632 a_4685_37583# a_5631_38127# 0.55fF
C12633 a_52778_39198# a_52778_39936# 0.35fF
C12634 a_18370_56170# ctopp 3.28fF
C12635 a_7803_55509# a_4339_64521# 0.50fF
C12636 a_24561_41583# VDD 0.91fF
C12637 vcm_commonmode a_17274_64202# 0.33fF
C12638 a_28410_17524# a_29414_17524# 0.97fF
C12639 a_12341_3311# a_22386_16520# 0.38fF
C12640 a_45478_21540# a_45478_20536# 1.00fF
C12641 a_11067_47695# a_12869_2741# 0.47fF
C12642 a_32426_24552# a_32426_23548# 1.00fF
C12643 a_49494_67214# VDD 1.12fF
C12644 a_17366_12504# a_17366_11500# 1.00fF
C12645 a_47486_12504# a_48490_12504# 0.97fF
C12646 a_32371_32117# VDD 0.47fF
C12647 a_10239_74575# VDD 0.58fF
C12648 a_28756_55394# a_12981_59343# 0.40fF
C12649 ctopn a_44474_21540# 3.59fF
C12650 a_29269_44545# VDD 1.30fF
C12651 a_39673_28111# a_40458_11500# 0.38fF
C12652 a_8575_74853# a_8003_72917# 0.63fF
C12653 a_3301_27791# VDD 0.55fF
C12654 a_16362_56170# VDD 2.48fF
C12655 vcm_commonmode a_37446_13508# 0.87fF
C12656 a_17366_61190# ctopp 3.43fF
C12657 ctopn a_21382_10496# 3.59fF
C12658 a_19374_69222# VDD 0.51fF
C12659 a_46482_9492# VDD 0.51fF
C12660 a_16362_16520# a_12727_13353# 1.27fF
C12661 vcm_commonmode a_23390_56170# 0.87fF
C12662 a_1895_14906# VDD 0.36fF
C12663 vcm_commonmode a_26310_69222# 0.31fF
C12664 a_41261_28335# a_12516_7093# 0.40fF
C12665 a_39362_7850# a_39454_7484# 0.32fF
C12666 a_26402_22544# VDD 0.51fF
C12667 a_6831_63303# a_25419_50959# 0.41fF
C12668 a_17366_65206# VDD 0.57fF
C12669 a_7295_44647# a_3339_30503# 0.69fF
C12670 a_32795_29967# VDD 0.39fF
C12671 a_11902_27497# a_11711_27247# 0.31fF
C12672 a_19967_41781# a_30855_41809# 1.80fF
C12673 a_8531_70543# a_2775_46025# 0.81fF
C12674 vcm_commonmode a_33338_22910# 0.31fF
C12675 a_21382_70226# ctopp 3.58fF
C12676 a_28446_31375# a_23736_7638# 0.87fF
C12677 a_7203_10383# VDD 1.13fF
C12678 a_38450_58178# ctopp 3.59fF
C12679 a_6607_42167# VDD 1.09fF
C12680 vcm_commonmode a_24302_65206# 0.31fF
C12681 a_23298_69222# a_23390_69222# 0.32fF
C12682 a_40491_27247# a_43470_10496# 0.38fF
C12683 a_29414_18528# a_29414_17524# 1.00fF
C12684 a_12641_36596# a_12713_36483# 0.72fF
C12685 a_42466_21540# a_43470_21540# 0.97fF
C12686 a_26523_28111# a_28305_28879# 0.31fF
C12687 a_20635_29415# a_25744_7638# 0.75fF
C12688 a_36797_27497# a_37446_23548# 0.38fF
C12689 a_1923_59583# a_10975_60975# 0.70fF
C12690 a_33338_64202# a_33430_64202# 0.32fF
C12691 a_7862_34025# VDD 10.64fF
C12692 ctopn a_16746_15514# 1.68fF
C12693 vcm_commonmode a_22386_61190# 0.87fF
C12694 a_22386_14512# VDD 0.51fF
C12695 a_12985_19087# a_12899_10927# 0.95fF
C12696 a_17366_55166# VDD 0.65fF
C12697 a_12341_3311# a_1586_18695# 0.85fF
C12698 a_30326_22910# a_30418_22544# 0.32fF
C12699 a_48490_64202# VDD 0.55fF
C12700 a_6835_46823# a_2606_41079# 1.80fF
C12701 a_6417_62215# a_7210_55081# 0.42fF
C12702 a_19374_10496# a_20378_10496# 0.97fF
C12703 vcm_commonmode a_29322_14878# 0.31fF
C12704 ctopn a_26402_11500# 3.59fF
C12705 a_21290_65206# a_21382_65206# 0.32fF
C12706 a_30418_14512# a_30418_13508# 1.00fF
C12707 a_33264_37601# VDD 1.72fF
C12708 a_3663_39991# VDD 0.39fF
C12709 a_12899_11471# a_12727_13353# 23.45fF
C12710 a_47486_17524# a_48490_17524# 0.97fF
C12711 a_7841_12167# a_10899_28879# 0.63fF
C12712 a_2595_47653# a_3983_48469# 0.72fF
C12713 vcm_commonmode a_26402_70226# 0.87fF
C12714 a_34434_60186# a_35438_60186# 0.97fF
C12715 a_27406_23548# VDD 0.52fF
C12716 a_24394_66210# VDD 0.51fF
C12717 a_36442_12504# a_36442_11500# 1.00fF
C12718 a_13143_29575# a_11430_26159# 0.31fF
C12719 a_16928_42919# a_13349_37973# 0.38fF
C12720 a_12947_56817# a_16746_56172# 0.37fF
C12721 vcm_commonmode a_34342_23914# 0.31fF
C12722 a_29414_7484# m3_29316_7346# 2.80fF
C12723 a_2040_43401# VDD 0.31fF
C12724 vcm_commonmode a_31330_66210# 0.31fF
C12725 a_23390_70226# a_23390_69222# 1.00fF
C12726 a_29414_18528# a_30418_18528# 0.97fF
C12727 a_36442_19532# VDD 0.51fF
C12728 a_15285_52245# VDD 0.52fF
C12729 a_3751_72373# a_4031_73095# 0.37fF
C12730 a_29760_7638# a_12877_16911# 0.41fF
C12731 vcm_commonmode a_43378_19898# 0.31fF
C12732 a_27406_67214# ctopp 3.59fF
C12733 a_8485_29673# a_7841_29673# 0.45fF
C12734 a_4811_34855# a_2787_30503# 0.84fF
C12735 a_22176_47919# VDD 0.31fF
C12736 a_21290_19898# a_21382_19532# 0.32fF
C12737 a_5671_21495# VDD 4.08fF
C12738 vcm_commonmode a_44474_8488# 0.86fF
C12739 m3_45380_7346# VDD 0.42fF
C12740 a_36629_27791# a_12895_13967# 0.41fF
C12741 a_17366_23548# m3_17268_23410# 2.77fF
C12742 a_22386_11500# a_22386_10496# 1.00fF
C12743 a_42985_46831# a_10515_22671# 0.40fF
C12744 a_26310_14878# a_26402_14512# 0.32fF
C12745 a_27337_38565# VDD 1.41fF
C12746 a_18127_35797# VDD 4.59fF
C12747 a_11803_55311# a_10975_66407# 1.08fF
C12748 a_42374_69222# a_42466_69222# 0.32fF
C12749 a_48490_18528# a_48490_17524# 1.00fF
C12750 a_2292_17179# VDD 6.63fF
C12751 a_30418_72234# a_31422_72234# 0.97fF
C12752 a_21371_50959# a_36613_48169# 1.04fF
C12753 a_20378_55166# a_21382_55166# 0.97fF
C12754 a_44382_24918# VDD 0.36fF
C12755 a_2840_53511# a_7764_53877# 0.77fF
C12756 a_14298_32143# VDD 0.76fF
C12757 a_8123_56399# a_7479_54439# 0.35fF
C12758 a_1775_60663# result_out[5] 0.31fF
C12759 a_3983_44655# VDD 0.44fF
C12760 vcm_commonmode a_32426_67214# 0.87fF
C12761 a_39454_20536# VDD 0.51fF
C12762 a_49402_22910# a_49494_22544# 0.32fF
C12763 a_28410_63198# VDD 0.57fF
C12764 a_38450_10496# a_39454_10496# 0.97fF
C12765 a_41967_31375# a_12985_7663# 0.41fF
C12766 a_40366_65206# a_40458_65206# 0.32fF
C12767 a_49494_14512# a_49494_13508# 1.00fF
C12768 a_1757_36501# VDD 0.66fF
C12769 vcm_commonmode a_46390_20902# 0.31fF
C12770 a_1761_25071# a_13716_43047# 4.08fF
C12771 a_25263_39913# VDD 0.62fF
C12772 vcm_commonmode a_35346_63198# 0.31fF
C12773 a_16955_52047# a_6835_46823# 1.01fF
C12774 a_32672_49007# VDD 0.47fF
C12775 a_26748_7638# a_26402_13508# 0.38fF
C12776 a_22386_59182# VDD 0.51fF
C12777 vcm_commonmode a_29414_9492# 0.87fF
C12778 m3_30320_72146# VDD 0.33fF
C12779 a_31330_23914# a_31422_23548# 0.32fF
C12780 a_4287_65540# VDD 0.36fF
C12781 a_5254_67503# a_4482_57863# 0.83fF
C12782 a_24394_11500# a_25398_11500# 0.97fF
C12783 vcm_commonmode a_45478_16520# 0.87fF
C12784 a_26402_64202# ctopp 3.59fF
C12785 ctopn a_31422_13508# 3.59fF
C12786 a_15193_41781# a_15931_39859# 0.34fF
C12787 a_33430_72234# VDD 1.62fF
C12788 a_36717_47375# a_12727_58255# 0.40fF
C12789 vcm_commonmode a_29322_59182# 0.31fF
C12790 a_28318_66210# a_28410_66210# 0.32fF
C12791 a_2787_30503# a_12340_29967# 0.36fF
C12792 a_33694_30761# a_38210_30199# 0.34fF
C12793 a_35815_31751# a_34759_31029# 0.31fF
C12794 vcm_commonmode m3_16264_71142# 3.05fF
C12795 a_39454_12504# VDD 0.51fF
C12796 a_15193_42917# VDD 1.75fF
C12797 a_42466_70226# a_42466_69222# 1.00fF
C12798 a_48490_18528# a_49494_18528# 0.97fF
C12799 a_11049_18543# VDD 0.60fF
C12800 a_35382_51157# VDD 0.41fF
C12801 vcm_commonmode a_38450_72234# 0.69fF
C12802 a_16270_72234# a_16362_72234# 0.33fF
C12803 a_24740_7638# a_24394_16520# 0.38fF
C12804 a_7571_29199# a_7755_26703# 0.50fF
C12805 a_12641_37684# a_13097_36367# 0.51fF
C12806 a_8373_26409# VDD 0.42fF
C12807 vcm_commonmode a_46390_12870# 0.31fF
C12808 a_17712_7638# a_17366_23548# 0.38fF
C12809 a_40675_27791# a_41462_23548# 0.38fF
C12810 a_28410_24552# a_29414_24552# 0.97fF
C12811 a_3187_34293# VDD 0.34fF
C12812 a_11067_66191# a_12659_54965# 1.13fF
C12813 a_3247_20495# a_2411_26133# 0.45fF
C12814 a_4191_33449# a_8491_41383# 1.39fF
C12815 a_40366_19898# a_40458_19532# 0.32fF
C12816 a_34434_21540# VDD 0.51fF
C12817 vcm_commonmode a_37446_7484# 0.69fF
C12818 a_2775_46025# a_3325_49551# 0.56fF
C12819 a_25398_62194# a_26402_62194# 0.97fF
C12820 a_41462_11500# a_41462_10496# 1.00fF
C12821 a_41261_28335# a_42466_59182# 0.38fF
C12822 a_45386_14878# a_45478_14512# 0.32fF
C12823 vcm_commonmode a_41370_21906# 0.31fF
C12824 a_35438_69222# ctopp 3.59fF
C12825 a_5441_27791# a_4248_29967# 0.43fF
C12826 vcm_commonmode a_31422_64202# 0.87fF
C12827 a_39454_17524# VDD 0.51fF
C12828 a_40050_48463# a_45478_72234# 0.34fF
C12829 a_14287_51175# a_18370_71230# 0.38fF
C12830 a_24302_20902# a_24394_20536# 0.32fF
C12831 a_26402_60186# VDD 0.51fF
C12832 a_38450_55166# a_39454_55166# 0.97fF
C12833 vcm_commonmode a_18278_10862# 0.31fF
C12834 a_33864_28111# a_12985_7663# 0.41fF
C12835 a_11067_63143# a_15439_49525# 0.31fF
C12836 vcm_commonmode a_46390_17890# 0.31fF
C12837 a_11067_67279# a_4792_20443# 0.31fF
C12838 a_33430_65206# ctopp 3.59fF
C12839 a_30418_57174# a_31422_57174# 0.97fF
C12840 vcm_commonmode a_33338_60186# 0.31fF
C12841 a_29760_55394# a_29414_61190# 0.38fF
C12842 a_33430_15516# a_34434_15516# 0.97fF
C12843 a_8491_27023# a_18370_11500# 0.38fF
C12844 a_25744_7638# a_25398_11500# 0.38fF
C12845 a_8104_18517# VDD 0.62fF
C12846 a_20635_29415# a_29175_28335# 0.50fF
C12847 a_18703_29199# a_12899_2767# 1.02fF
C12848 a_13837_39860# a_13669_37429# 0.61fF
C12849 a_5085_24759# a_4417_22671# 0.41fF
C12850 a_1929_10651# a_3063_9295# 0.40fF
C12851 a_17803_36649# VDD 0.59fF
C12852 vcm_commonmode a_19374_19532# 0.87fF
C12853 a_23395_52047# a_12869_2741# 2.16fF
C12854 a_41872_29423# a_43470_64202# 0.38fF
C12855 a_34711_47375# VDD 0.43fF
C12856 a_31422_71230# a_32426_71230# 0.97fF
C12857 vcm_commonmode a_40458_69222# 0.87fF
C12858 a_42718_27497# a_44474_14512# 0.38fF
C12859 a_38450_58178# a_38557_32143# 0.38fF
C12860 a_2794_62697# a_7523_62581# 0.48fF
C12861 a_43470_11500# a_44474_11500# 0.97fF
C12862 a_25787_28327# a_13643_28327# 1.35fF
C12863 a_47394_66210# a_47486_66210# 0.32fF
C12864 vcm_commonmode a_47486_22544# 0.87fF
C12865 vcm_commonmode m3_16264_18390# 3.21fF
C12866 a_16362_11500# VDD 2.49fF
C12867 a_8491_41383# a_12447_29199# 2.63fF
C12868 a_33819_42359# VDD 0.61fF
C12869 vcm_commonmode a_38450_65206# 0.87fF
C12870 a_40458_18528# VDD 0.51fF
C12871 a_33261_51433# VDD 0.38fF
C12872 a_20378_24552# VDD 0.60fF
C12873 vcm_commonmode a_23298_11866# 0.31fF
C12874 ctopn a_38450_8488# 3.40fF
C12875 a_42709_29199# a_12985_7663# 0.40fF
C12876 a_40675_27791# a_11067_21583# 0.41fF
C12877 a_24302_12870# a_24394_12504# 0.32fF
C12878 a_29119_34473# VDD 0.56fF
C12879 vcm_commonmode a_47394_18894# 0.31fF
C12880 a_40458_66210# ctopp 3.59fF
C12881 a_12907_56399# a_6775_53877# 1.78fF
C12882 vcm_commonmode a_27314_24918# 0.31fF
C12883 a_19374_59182# a_19374_58178# 1.00fF
C12884 a_31422_55166# VDD 0.60fF
C12885 a_44474_62194# a_45478_62194# 0.97fF
C12886 a_23298_28487# VDD 0.48fF
C12887 a_22386_57174# VDD 0.51fF
C12888 vcm_commonmode a_43470_14512# 0.87fF
C12889 a_21371_52263# a_26402_58178# 0.38fF
C12890 a_6883_37019# VDD 2.03fF
C12891 vcm_commonmode a_22386_20536# 0.87fF
C12892 vcm_commonmode a_37354_55166# 0.30fF
C12893 a_49494_10496# VDD 1.12fF
C12894 a_43267_31055# a_46482_65206# 0.38fF
C12895 vcm_commonmode a_29322_57174# 0.31fF
C12896 a_26397_51183# a_30125_47919# 0.35fF
C12897 a_5039_42167# VDD 4.80fF
C12898 a_34434_72234# a_34434_71230# 1.00fF
C12899 a_42985_46831# a_12901_66665# 0.40fF
C12900 a_43378_20902# a_43470_20536# 0.32fF
C12901 a_2865_58799# VDD 0.59fF
C12902 a_2411_26133# a_1591_29973# 0.34fF
C12903 a_9503_26151# a_12985_7663# 0.41fF
C12904 VDD config_1_in[12] 1.05fF
C12905 a_32334_63198# a_32426_63198# 0.32fF
C12906 a_23390_57174# a_23390_56170# 1.00fF
C12907 a_10883_71855# VDD 0.42fF
C12908 vcm_commonmode a_48490_23548# 0.88fF
C12909 a_2235_30503# a_23195_29967# 0.31fF
C12910 a_24515_43493# VDD 1.02fF
C12911 vcm_commonmode a_45478_66210# 0.87fF
C12912 a_2216_28309# a_4242_35407# 0.44fF
C12913 a_38115_52263# VDD 3.21fF
C12914 a_19282_21906# a_19374_21540# 0.32fF
C12915 a_36442_62194# VDD 0.51fF
C12916 a_22808_27497# VDD 0.43fF
C12917 vcm_commonmode a_22386_12504# 0.87fF
C12918 ctopn a_23390_9492# 3.58fF
C12919 a_4211_67655# VDD 1.05fF
C12920 ctopn a_39454_16520# 3.59fF
C12921 a_18151_52263# a_6775_53877# 1.32fF
C12922 a_1761_43567# a_1803_19087# 0.48fF
C12923 vcm_commonmode a_43378_62194# 0.31fF
C12924 a_41261_28335# a_42466_57174# 0.38fF
C12925 a_44474_15516# VDD 0.51fF
C12926 a_43362_28879# a_47486_70226# 0.38fF
C12927 a_8583_33551# a_2021_22325# 0.53fF
C12928 a_26310_59182# a_26402_59182# 0.32fF
C12929 a_6913_64239# VDD 0.39fF
C12930 a_44474_63198# ctopp 3.64fF
C12931 a_11619_3303# a_12349_25847# 0.47fF
C12932 a_42466_71230# VDD 0.58fF
C12933 a_39299_48783# a_12901_58799# 0.40fF
C12934 vcm_commonmode a_17366_21540# 1.82fF
C12935 a_33641_29967# a_34759_31029# 1.48fF
C12936 a_37446_72234# m3_37348_72146# 2.80fF
C12937 a_7464_39215# VDD 0.77fF
C12938 a_33864_28111# a_34434_8488# 0.38fF
C12939 a_24302_17890# a_24394_17524# 0.32fF
C12940 a_26748_7638# a_26402_7484# 0.34fF
C12941 a_14831_50095# a_19885_50095# 0.69fF
C12942 a_36350_72234# a_36442_72234# 0.32fF
C12943 vcm_commonmode a_49402_71230# 0.30fF
C12944 a_5363_30503# a_16917_31573# 0.35fF
C12945 a_38450_59182# ctopp 3.59fF
C12946 a_30418_64202# a_30418_63198# 1.23fF
C12947 a_1923_59583# a_4187_60673# 0.34fF
C12948 a_43378_12870# a_43470_12504# 0.32fF
C12949 a_25321_29673# VDD 3.04fF
C12950 vcm_commonmode a_22386_17524# 0.87fF
C12951 a_5483_74244# VDD 0.47fF
C12952 a_42985_46831# a_48490_62194# 0.38fF
C12953 a_17507_52047# a_12981_59343# 0.40fF
C12954 a_21382_13508# VDD 0.51fF
C12955 a_3987_19623# VDD 11.42fF
C12956 a_2012_33927# a_1761_30511# 0.97fF
C12957 a_22386_22544# a_22386_21540# 1.00fF
C12958 a_1586_36727# a_1683_33237# 0.43fF
C12959 vcm_commonmode a_28318_13874# 0.31fF
C12960 a_29414_13508# a_30418_13508# 0.97fF
C12961 a_20713_36929# VDD 1.72fF
C12962 a_12725_44527# a_12381_43957# 0.63fF
C12963 a_43362_28879# a_12355_15055# 0.40fF
C12964 a_34434_68218# a_35438_68218# 0.97fF
C12965 vcm_commonmode a_49494_63198# 1.06fF
C12966 a_12877_16911# a_12727_15529# 23.51fF
C12967 a_20359_29199# a_12907_27023# 0.58fF
C12968 a_8643_48767# VDD 0.52fF
C12969 vcm_commonmode a_16362_69222# 4.47fF
C12970 a_34251_52263# a_12516_7093# 0.40fF
C12971 a_46482_56170# a_46482_55166# 1.00fF
C12972 a_42466_57174# a_42466_56170# 1.00fF
C12973 a_44382_72234# VDD 0.62fF
C12974 vcm_commonmode a_43470_59182# 0.87fF
C12975 a_37551_42333# VDD 2.00fF
C12976 a_17039_51157# a_26155_50095# 0.70fF
C12977 a_12899_10927# VDD 8.33fF
C12978 vcm_commonmode a_49494_72234# 0.72fF
C12979 a_28756_7638# a_12727_15529# 0.41fF
C12980 a_38358_21906# a_38450_21540# 0.32fF
C12981 a_19807_28111# a_30764_7638# 0.69fF
C12982 a_7343_25615# VDD 0.67fF
C12983 a_19374_58178# a_19374_57174# 1.00fF
C12984 a_42466_60186# ctopp 3.59fF
C12985 ctopn a_12947_8725# 1.23fF
C12986 a_45478_68218# VDD 0.51fF
C12987 vcm_commonmode a_23390_18528# 0.87fF
C12988 a_16362_66210# ctopp 1.35fF
C12989 a_45386_7850# VDD 0.63fF
C12990 a_26402_16520# a_26402_15516# 1.00fF
C12991 ctopn a_41462_22544# 3.58fF
C12992 a_2235_30503# a_16087_31751# 0.36fF
C12993 a_20635_29415# a_26523_28111# 0.48fF
C12994 a_3327_9308# VDD 5.34fF
C12995 a_20267_30503# VDD 12.39fF
C12996 a_45386_59182# a_45478_59182# 0.32fF
C12997 a_28963_28853# VDD 0.45fF
C12998 a_16746_65208# a_16362_65206# 2.28fF
C12999 a_14425_37981# VDD 0.90fF
C13000 vcm_commonmode a_16270_55166# 0.32fF
C13001 a_3024_67191# a_5024_67885# 1.47fF
C13002 a_1586_66567# a_1757_66415# 0.60fF
C13003 a_43378_17890# a_43470_17524# 0.32fF
C13004 vcm_commonmode a_17274_70226# 0.33fF
C13005 a_30326_60186# a_30418_60186# 0.32fF
C13006 vcm_commonmode a_32426_10496# 0.87fF
C13007 a_49494_64202# a_49494_63198# 1.23fF
C13008 a_12355_15055# a_16746_62196# 0.41fF
C13009 a_35431_31751# VDD 0.44fF
C13010 ctopn a_37446_14512# 3.59fF
C13011 a_1586_21959# a_1757_26159# 0.61fF
C13012 a_1586_36727# config_2_in[5] 0.48fF
C13013 a_6271_72943# VDD 0.46fF
C13014 vcm_commonmode a_47486_60186# 0.87fF
C13015 a_20378_71230# ctopp 3.40fF
C13016 ctopn a_16362_20536# 1.35fF
C13017 a_22386_7484# m3_22288_7346# 2.80fF
C13018 a_25306_18894# a_25398_18528# 0.32fF
C13019 a_1923_73087# a_1823_72381# 1.40fF
C13020 a_41462_22544# a_41462_21540# 1.00fF
C13021 a_45478_56170# VDD 0.52fF
C13022 a_48490_13508# a_49494_13508# 0.97fF
C13023 a_28410_8488# VDD 0.58fF
C13024 a_1761_25071# a_32327_40191# 0.40fF
C13025 a_1689_10396# a_2004_42453# 3.70fF
C13026 vcm_commonmode a_19374_62194# 0.87fF
C13027 a_20378_68218# a_20378_67214# 1.00fF
C13028 a_43267_31055# a_12257_56623# 0.40fF
C13029 ctopn a_42466_23548# 3.40fF
C13030 a_16746_19530# a_12895_13967# 2.28fF
C13031 a_11883_58575# VDD 0.40fF
C13032 vcm_commonmode a_35346_8854# 0.31fF
C13033 m3_17268_7346# VDD 0.42fF
C13034 a_2847_30271# VDD 0.39fF
C13035 vcm_commonmode a_27406_15516# 0.87fF
C13036 ctopn a_16362_12504# 1.35fF
C13037 a_38450_57174# ctopp 3.58fF
C13038 a_34434_56170# a_35438_56170# 0.97fF
C13039 a_41427_52263# a_10515_22671# 0.40fF
C13040 a_2292_17179# a_3247_10389# 0.42fF
C13041 a_19626_31751# a_31084_30485# 1.09fF
C13042 a_23395_52047# a_28756_55394# 0.32fF
C13043 vcm_commonmode a_25398_71230# 0.86fF
C13044 a_44474_61190# VDD 0.51fF
C13045 a_17274_55166# a_17366_55166# 0.32fF
C13046 a_17366_8488# a_18370_8488# 0.97fF
C13047 vcm_commonmode a_37446_11500# 0.87fF
C13048 a_11803_55311# a_1803_20719# 0.89fF
C13049 a_12983_63151# VDD 7.28fF
C13050 a_12516_7093# a_12869_2741# 0.47fF
C13051 a_16510_8760# a_11067_21583# 1.09fF
C13052 a_45478_16520# a_45478_15516# 1.00fF
C13053 vcm_commonmode a_41462_24552# 0.84fF
C13054 a_28756_55394# a_8583_33551# 1.05fF
C13055 a_1761_50639# a_1761_43567# 0.31fF
C13056 a_18370_70226# a_19374_70226# 0.97fF
C13057 vcm_commonmode a_23298_67214# 0.31fF
C13058 a_30418_19532# a_30418_18528# 1.00fF
C13059 a_5795_27497# VDD 0.55fF
C13060 a_34342_10862# a_34434_10496# 0.32fF
C13061 a_19720_7638# a_19374_24552# 0.46fF
C13062 a_48490_70226# VDD 0.54fF
C13063 a_28747_37503# VDD 0.92fF
C13064 a_23390_68218# ctopp 3.59fF
C13065 ctopn a_16746_17522# 1.68fF
C13066 a_13669_39605# VDD 5.03fF
C13067 vcm_commonmode a_43470_57174# 0.87fF
C13068 a_29414_16520# VDD 0.51fF
C13069 a_9063_71553# a_9024_71427# 0.75fF
C13070 a_1768_13103# config_2_in[5] 0.63fF
C13071 a_10607_58799# VDD 0.32fF
C13072 a_12727_58255# a_16746_59184# 2.28fF
C13073 a_49402_60186# a_49494_60186# 0.32fF
C13074 vcm_commonmode a_20286_9858# 0.31fF
C13075 a_31768_7638# a_12985_19087# 0.41fF
C13076 a_17488_48731# a_17672_32259# 0.71fF
C13077 a_20286_11866# a_20378_11500# 0.32fF
C13078 a_10055_58791# a_23736_7638# 0.41fF
C13079 vcm_commonmode a_36350_16886# 0.31fF
C13080 a_26402_72234# VDD 1.38fF
C13081 a_29760_55394# a_12727_58255# 0.40fF
C13082 VDD result_out[6] 0.66fF
C13083 a_25398_15516# a_25398_14512# 1.00fF
C13084 a_8583_33551# m2_48260_24282# 0.39fF
C13085 a_12713_43011# VDD 1.07fF
C13086 a_44382_18894# a_44474_18528# 0.32fF
C13087 a_39673_28111# a_40458_10496# 0.38fF
C13088 vcm_commonmode a_31422_72234# 0.69fF
C13089 a_33430_61190# a_34434_61190# 0.97fF
C13090 a_24302_24918# a_24394_24552# 0.32fF
C13091 a_36629_27791# a_36442_23548# 0.38fF
C13092 a_6649_25615# a_7755_26703# 0.56fF
C13093 a_21382_7484# VDD 1.58fF
C13094 a_39454_68218# a_39454_67214# 1.00fF
C13095 a_7862_34025# a_9307_30663# 0.35fF
C13096 VDD result_out[15] 0.59fF
C13097 a_17787_47349# VDD 0.57fF
C13098 vcm_commonmode a_28410_68218# 0.87fF
C13099 a_29760_7638# a_12895_13967# 0.41fF
C13100 a_30764_7638# a_12985_19087# 0.41fF
C13101 a_5490_41365# a_1761_37039# 0.65fF
C13102 a_21290_62194# a_21382_62194# 0.32fF
C13103 a_1643_29397# VDD 0.33fF
C13104 a_11430_26159# a_12349_25847# 1.19fF
C13105 a_23390_56170# ctopp 3.40fF
C13106 a_7213_62215# a_2840_53511# 1.25fF
C13107 a_38557_32143# a_38450_59182# 0.38fF
C13108 ctopn a_17366_18528# 3.43fF
C13109 a_7281_29423# a_6162_28487# 0.69fF
C13110 a_17358_31069# a_17507_30761# 0.48fF
C13111 vcm_commonmode a_22294_64202# 0.31fF
C13112 a_24394_69222# a_24394_68218# 1.00fF
C13113 a_2292_17179# a_3023_16341# 0.34fF
C13114 a_37919_28111# a_38450_15516# 0.38fF
C13115 a_34342_55166# a_34434_55166# 0.33fF
C13116 a_36442_8488# a_37446_8488# 0.97fF
C13117 a_4339_64521# a_9271_52789# 0.34fF
C13118 a_7676_61493# a_2794_62697# 0.55fF
C13119 a_26310_57174# a_26402_57174# 0.32fF
C13120 a_21371_50959# a_25398_61190# 0.38fF
C13121 a_29322_15882# a_29414_15516# 0.32fF
C13122 a_37446_70226# a_38450_70226# 0.97fF
C13123 a_49494_19532# a_49494_18528# 1.00fF
C13124 ctopn a_27752_7638# 2.62fF
C13125 a_19720_7638# a_12877_16911# 0.41fF
C13126 a_7369_24233# VDD 1.28fF
C13127 vcm_commonmode a_42466_13508# 0.87fF
C13128 a_22386_61190# ctopp 3.59fF
C13129 a_48490_59182# a_48490_58178# 1.00fF
C13130 ctopn a_26402_10496# 3.59fF
C13131 a_24394_69222# VDD 0.51fF
C13132 a_1591_36103# VDD 0.41fF
C13133 a_1770_14441# a_1823_54973# 0.84fF
C13134 a_16955_52047# a_12869_2741# 0.79fF
C13135 a_11619_56615# a_12983_63151# 0.32fF
C13136 a_39389_52271# a_39454_64202# 0.38fF
C13137 a_18370_16520# a_19374_16520# 0.97fF
C13138 vcm_commonmode a_28410_56170# 0.87fF
C13139 vcm_commonmode a_31330_69222# 0.31fF
C13140 a_27314_71230# a_27406_71230# 0.32fF
C13141 a_36797_27497# a_37446_14512# 0.38fF
C13142 a_35438_60186# a_35438_59182# 1.00fF
C13143 a_31422_22544# VDD 0.51fF
C13144 a_22386_65206# VDD 0.51fF
C13145 a_24394_63198# a_24394_62194# 1.00fF
C13146 a_7019_30511# VDD 0.56fF
C13147 a_39362_11866# a_39454_11500# 0.32fF
C13148 a_23736_7638# a_23390_23548# 0.38fF
C13149 a_5254_67503# a_7676_61493# 0.37fF
C13150 a_4119_70741# a_6361_57711# 0.38fF
C13151 a_13183_52047# a_12901_58799# 0.40fF
C13152 a_44474_15516# a_44474_14512# 1.00fF
C13153 vcm_commonmode a_38358_22910# 0.31fF
C13154 a_26402_70226# ctopp 3.58fF
C13155 a_8753_31055# a_10506_29967# 0.36fF
C13156 a_1867_10927# VDD 0.51fF
C13157 a_6863_42692# a_1761_22895# 0.62fF
C13158 vcm_commonmode a_29322_65206# 0.31fF
C13159 a_43267_31055# a_10975_66407# 0.40fF
C13160 a_35601_27497# a_12727_13353# 0.41fF
C13161 a_5363_30503# a_7862_34025# 0.57fF
C13162 a_29414_9492# a_29414_8488# 1.00fF
C13163 a_40675_27791# a_12546_22351# 0.41fF
C13164 a_43378_24918# a_43470_24552# 0.32fF
C13165 a_11943_63125# a_10515_63143# 1.06fF
C13166 ctopn a_21382_15516# 3.59fF
C13167 a_21371_50959# a_4215_51157# 0.55fF
C13168 a_1586_36727# a_6725_42479# 0.36fF
C13169 a_24394_67214# a_25398_67214# 0.97fF
C13170 vcm_commonmode a_27406_61190# 0.87fF
C13171 a_4495_35925# a_4248_29967# 0.60fF
C13172 a_27406_14512# VDD 0.51fF
C13173 a_26748_7638# a_26402_11500# 0.38fF
C13174 a_19576_51701# a_27627_51733# 0.34fF
C13175 a_3799_20407# VDD 0.43fF
C13176 a_22294_55166# VDD 0.35fF
C13177 a_24740_7638# a_12899_10927# 0.41fF
C13178 a_21187_29415# a_12899_2767# 0.31fF
C13179 a_7295_44647# a_16101_31029# 0.33fF
C13180 a_40366_62194# a_40458_62194# 0.32fF
C13181 a_9731_22895# VDD 3.77fF
C13182 vcm_commonmode a_34342_14878# 0.31fF
C13183 ctopn a_31422_11500# 3.59fF
C13184 a_17599_52263# a_22386_58178# 0.38fF
C13185 a_41636_37601# VDD 1.83fF
C13186 a_1586_66567# a_9624_65301# 0.34fF
C13187 a_43470_69222# a_43470_68218# 1.00fF
C13188 a_41261_28335# a_42466_65206# 0.38fF
C13189 a_10405_16367# VDD 0.31fF
C13190 a_22989_48437# a_23847_47919# 0.36fF
C13191 vcm_commonmode a_31422_70226# 0.87fF
C13192 a_41427_52263# a_12901_66665# 0.40fF
C13193 a_30418_72234# a_30418_71230# 1.00fF
C13194 a_40491_27247# a_43470_15516# 0.38fF
C13195 a_32426_23548# VDD 0.52fF
C13196 a_33430_8488# a_33430_7484# 1.00fF
C13197 a_29414_66210# VDD 0.51fF
C13198 a_19004_40413# a_19967_41781# 0.44fF
C13199 a_45386_57174# a_45478_57174# 0.32fF
C13200 a_17274_72234# VDD 0.64fF
C13201 a_2191_68565# a_3295_62083# 0.99fF
C13202 a_48398_15882# a_48490_15516# 0.32fF
C13203 vcm_commonmode a_39362_23914# 0.31fF
C13204 a_11455_12157# VDD 0.48fF
C13205 a_1586_36727# VDD 5.33fF
C13206 vcm_commonmode a_36350_66210# 0.31fF
C13207 a_26402_58178# a_27406_58178# 0.97fF
C13208 a_41462_19532# VDD 0.51fF
C13209 a_12869_2741# a_15607_46805# 1.19fF
C13210 a_40491_27247# a_12877_16911# 0.41fF
C13211 a_21382_9492# a_22386_9492# 0.97fF
C13212 a_2840_66103# a_10687_52553# 2.01fF
C13213 a_35601_27497# a_10515_23975# 0.41fF
C13214 a_25300_39655# a_1799_29556# 0.34fF
C13215 a_3983_68591# VDD 0.40fF
C13216 a_7213_62215# a_6417_62215# 0.89fF
C13217 a_22386_13508# a_22386_12504# 1.00fF
C13218 a_20927_35877# VDD 0.85fF
C13219 vcm_commonmode a_48398_19898# 0.31fF
C13220 a_32426_67214# ctopp 3.59fF
C13221 a_13390_29575# a_13239_29575# 0.33fF
C13222 a_37446_16520# a_38450_16520# 0.97fF
C13223 a_12546_22351# a_16362_9492# 19.89fF
C13224 a_38557_32143# a_38450_57174# 0.38fF
C13225 a_46390_71230# a_46482_71230# 0.32fF
C13226 a_41872_29423# a_43470_70226# 0.38fF
C13227 vcm_commonmode a_49494_8488# 0.89fF
C13228 a_4339_64521# a_9431_60214# 0.30fF
C13229 a_43470_63198# a_43470_62194# 1.00fF
C13230 a_27752_7638# a_27406_24552# 0.47fF
C13231 vcm_commonmode a_20378_58178# 0.87fF
C13232 a_36613_48169# a_12901_58799# 0.40fF
C13233 a_35932_38689# VDD 1.58fF
C13234 a_1761_47919# a_13067_38517# 6.11fF
C13235 a_4674_40277# a_3247_20495# 0.92fF
C13236 a_40050_48463# a_45478_66210# 0.38fF
C13237 ctopn a_8491_27023# 2.61fF
C13238 a_2686_70223# a_7289_70767# 0.37fF
C13239 a_3339_43023# a_12907_27023# 0.42fF
C13240 a_48490_9492# a_48490_8488# 1.00fF
C13241 a_25744_7638# a_11067_21583# 0.41fF
C13242 a_27535_30503# a_30788_28487# 0.48fF
C13243 a_48490_58178# a_48490_57174# 1.00fF
C13244 a_43470_67214# a_44474_67214# 0.97fF
C13245 a_39299_48783# a_44474_62194# 0.38fF
C13246 a_7695_31573# a_12215_31573# 0.47fF
C13247 a_4443_46607# a_4563_32900# 0.90fF
C13248 vcm_commonmode a_37446_67214# 0.87fF
C13249 a_12251_39069# a_12621_36091# 0.52fF
C13250 a_44474_20536# VDD 0.51fF
C13251 a_33430_63198# VDD 0.57fF
C13252 a_25306_13874# a_25398_13508# 0.32fF
C13253 a_28757_27247# a_30975_28023# 0.38fF
C13254 a_26523_29199# a_12263_4391# 0.38fF
C13255 a_39449_39868# VDD 1.15fF
C13256 vcm_commonmode a_40366_63198# 0.31fF
C13257 a_39222_48169# a_12355_15055# 0.40fF
C13258 a_30326_68218# a_30418_68218# 0.32fF
C13259 a_28756_55394# a_12516_7093# 0.40fF
C13260 a_17712_7638# a_17366_14512# 0.38fF
C13261 a_40675_27791# a_41462_14512# 0.38fF
C13262 a_27406_59182# VDD 0.51fF
C13263 a_8583_33551# a_8491_41383# 0.44fF
C13264 a_29414_7484# a_30418_7484# 0.97fF
C13265 vcm_commonmode a_34434_9492# 0.87fF
C13266 m3_45380_72146# VDD 0.42fF
C13267 a_7187_23439# a_6816_19355# 0.38fF
C13268 a_1768_13103# VDD 7.85fF
C13269 a_42466_24552# m3_42368_24414# 2.81fF
C13270 a_31422_64202# ctopp 3.59fF
C13271 ctopn a_36442_13508# 3.59fF
C13272 a_37354_72234# VDD 0.63fF
C13273 a_1923_59583# a_3983_65327# 0.34fF
C13274 vcm_commonmode a_34342_59182# 0.31fF
C13275 a_15548_30761# a_13353_30511# 0.84fF
C13276 a_44474_12504# VDD 0.51fF
C13277 a_8491_27023# a_18370_10496# 0.38fF
C13278 a_25744_7638# a_25398_10496# 0.38fF
C13279 a_1761_39215# a_12621_36091# 3.01fF
C13280 a_40458_9492# a_41462_9492# 0.97fF
C13281 a_23390_64202# a_24394_64202# 0.97fF
C13282 a_41462_13508# a_41462_12504# 1.00fF
C13283 a_11521_66567# a_11619_63151# 0.31fF
C13284 a_4812_13879# VDD 3.00fF
C13285 a_1586_45431# a_5831_39189# 0.53fF
C13286 a_5682_69367# a_5213_70223# 0.31fF
C13287 a_39454_21540# VDD 0.51fF
C13288 vcm_commonmode a_42466_7484# 0.69fF
C13289 a_20378_22544# a_21382_22544# 0.97fF
C13290 a_7295_44647# a_14926_31849# 0.38fF
C13291 a_11140_10107# a_11179_9981# 0.76fF
C13292 a_4758_45369# a_10680_52245# 0.73fF
C13293 vcm_commonmode a_46390_21906# 0.31fF
C13294 a_40458_69222# ctopp 3.59fF
C13295 a_16362_10496# VDD 2.47fF
C13296 vcm_commonmode a_36442_64202# 0.87fF
C13297 a_44474_17524# VDD 0.51fF
C13298 a_18151_52263# a_12907_56399# 2.67fF
C13299 a_31422_60186# VDD 0.51fF
C13300 a_2007_21237# VDD 0.41fF
C13301 vcm_commonmode a_23298_10862# 0.31fF
C13302 a_6651_31599# VDD 0.42fF
C13303 a_10515_63143# a_9179_22351# 0.34fF
C13304 a_38450_65206# ctopp 3.59fF
C13305 a_12899_3311# a_28756_7638# 0.67fF
C13306 a_2235_41941# a_2411_26133# 0.34fF
C13307 vcm_commonmode a_38358_60186# 0.31fF
C13308 a_31422_67214# a_31422_66210# 1.00fF
C13309 a_2292_43291# a_1803_20719# 0.51fF
C13310 a_11395_62037# VDD 0.41fF
C13311 a_12907_27023# a_12631_28585# 0.93fF
C13312 a_12641_37684# a_1761_37039# 3.02fF
C13313 a_10055_58791# a_39673_28111# 0.41fF
C13314 a_49494_64202# m3_49396_64114# 2.78fF
C13315 a_27406_65206# a_27406_64202# 1.00fF
C13316 a_44382_13874# a_44474_13508# 0.32fF
C13317 a_29207_36415# VDD 0.86fF
C13318 vcm_commonmode a_24394_19532# 0.87fF
C13319 a_49402_68218# a_49494_68218# 0.32fF
C13320 a_39389_52271# a_12257_56623# 0.40fF
C13321 vcm_commonmode a_45478_69222# 0.87fF
C13322 a_4831_58497# VDD 0.42fF
C13323 a_7571_26151# a_10515_23975# 0.72fF
C13324 a_48490_7484# a_49494_7484# 0.97fF
C13325 m3_49396_21402# VDD 0.34fF
C13326 a_21382_23548# a_21382_22544# 1.00fF
C13327 vcm_commonmode a_18278_15882# 0.31fF
C13328 a_41427_52263# a_19807_28111# 5.99fF
C13329 a_17278_28309# a_17712_7638# 0.51fF
C13330 a_42709_29199# a_9503_26151# 0.35fF
C13331 a_30326_56170# a_30418_56170# 0.32fF
C13332 a_34780_56398# a_10515_22671# 0.40fF
C13333 a_21382_11500# VDD 0.51fF
C13334 a_32426_69222# a_33430_69222# 0.97fF
C13335 vcm_commonmode a_43470_65206# 0.87fF
C13336 a_2952_66139# a_6515_67477# 0.36fF
C13337 a_12895_13967# a_12727_15529# 0.38fF
C13338 a_12473_36341# a_1761_31055# 4.13fF
C13339 a_45478_18528# VDD 0.51fF
C13340 a_35676_49525# a_34145_49007# 0.38fF
C13341 vcm_commonmode a_11803_55311# 16.84fF
C13342 a_23390_72234# a_24394_72234# 0.97fF
C13343 a_12641_37684# a_1761_32143# 1.18fF
C13344 a_1799_29556# a_13669_35253# 0.38fF
C13345 a_27406_61190# a_27406_60186# 1.00fF
C13346 a_25398_24552# VDD 0.60fF
C13347 vcm_commonmode a_28318_11866# 0.31fF
C13348 ctopn a_43470_8488# 3.40fF
C13349 a_1770_14441# VDD 8.36fF
C13350 a_42466_64202# a_43470_64202# 0.97fF
C13351 a_4035_33205# VDD 0.30fF
C13352 a_4528_26159# config_1_in[15] 0.42fF
C13353 a_45478_66210# ctopp 3.59fF
C13354 a_47486_55166# m2_48260_54946# 0.92fF
C13355 a_16510_8760# a_12546_22351# 1.08fF
C13356 vcm_commonmode a_32334_24918# 0.31fF
C13357 a_5239_45717# VDD 0.57fF
C13358 a_1591_18543# a_2411_18517# 0.34fF
C13359 a_35438_55166# VDD 0.60fF
C13360 a_9955_21807# a_5671_21495# 0.59fF
C13361 a_39454_22544# a_40458_22544# 0.97fF
C13362 a_9643_63125# VDD 0.65fF
C13363 a_31768_7638# VDD 6.39fF
C13364 a_27406_57174# VDD 0.51fF
C13365 vcm_commonmode a_48490_14512# 0.87fF
C13366 a_1768_13103# a_2944_64488# 0.40fF
C13367 a_30418_65206# a_31422_65206# 0.97fF
C13368 a_1923_59583# a_2163_63293# 0.32fF
C13369 a_16152_37601# VDD 1.98fF
C13370 vcm_commonmode a_27406_20536# 0.87fF
C13371 vcm_commonmode a_42374_55166# 0.30fF
C13372 a_51330_39932# VDD 0.44fF
C13373 vcm_commonmode a_12981_62313# 6.23fF
C13374 a_26402_17524# a_26402_16520# 1.00fF
C13375 vcm_commonmode a_34342_57174# 0.31fF
C13376 a_20195_49793# a_20156_49667# 0.72fF
C13377 a_1591_71317# a_1757_71317# 0.42fF
C13378 a_4119_70741# a_5208_70063# 0.33fF
C13379 a_7107_58487# VDD 1.00fF
C13380 a_7059_24135# a_6816_19355# 0.61fF
C13381 a_21382_23548# a_22386_23548# 0.97fF
C13382 VDD config_1_in[7] 0.92fF
C13383 a_19807_28111# a_20881_28111# 1.08fF
C13384 a_30418_56170# a_30418_55166# 1.00fF
C13385 a_10506_29967# VDD 1.51fF
C13386 a_12725_44527# a_36708_39655# 0.32fF
C13387 a_19374_72234# VDD 1.23fF
C13388 a_18370_66210# a_19374_66210# 0.97fF
C13389 a_17599_52263# a_12727_58255# 0.40fF
C13390 a_13183_52047# a_2840_66103# 1.72fF
C13391 a_8531_70543# a_11067_67279# 2.26fF
C13392 a_2099_59861# a_2004_42453# 0.54fF
C13393 a_2339_38129# a_5085_24759# 0.40fF
C13394 a_1867_51727# VDD 0.45fF
C13395 vcm_commonmode a_24394_72234# 0.69fF
C13396 a_41462_62194# VDD 0.51fF
C13397 a_29322_61190# a_29414_61190# 0.32fF
C13398 a_30764_7638# VDD 7.67fF
C13399 vcm_commonmode a_27406_12504# 0.87fF
C13400 ctopn a_28410_9492# 3.58fF
C13401 a_8772_63927# VDD 1.89fF
C13402 a_46482_65206# a_46482_64202# 1.00fF
C13403 ctopn a_44474_16520# 3.59fF
C13404 vcm_commonmode a_48398_62194# 0.31fF
C13405 a_11067_67279# a_10975_66407# 0.69fF
C13406 a_49494_15516# VDD 1.13fF
C13407 vcm_commonmode a_19282_68218# 0.31fF
C13408 a_18370_71230# a_18370_70226# 1.00fF
C13409 a_30418_19532# a_31422_19532# 0.97fF
C13410 a_40458_23548# a_40458_22544# 1.00fF
C13411 a_4127_63669# VDD 0.36fF
C13412 a_16746_62196# a_16362_62194# 2.28fF
C13413 m2_48260_54946# VDD 0.40fF
C13414 a_49402_56170# a_49494_56170# 0.32fF
C13415 a_47486_71230# VDD 0.58fF
C13416 a_34780_56398# a_34434_59182# 0.38fF
C13417 a_34434_66210# a_34434_65206# 1.00fF
C13418 a_35438_14512# a_36442_14512# 0.97fF
C13419 vcm_commonmode a_22386_21540# 0.87fF
C13420 a_16362_69222# ctopp 1.35fF
C13421 a_40458_72234# m3_40360_72146# 2.80fF
C13422 a_1586_69367# a_1591_57711# 0.30fF
C13423 a_38557_32143# a_38450_72234# 0.34fF
C13424 a_11521_58951# VDD 0.95fF
C13425 a_46482_61190# a_46482_60186# 1.00fF
C13426 a_32334_8854# a_32426_8488# 0.32fF
C13427 a_43470_59182# ctopp 3.59fF
C13428 vcm_commonmode a_27406_17524# 0.87fF
C13429 a_10109_73487# VDD 0.45fF
C13430 a_17507_52047# a_21382_61190# 0.38fF
C13431 a_20905_32143# a_20881_28111# 0.55fF
C13432 a_26402_13508# VDD 0.51fF
C13433 a_12621_44099# VDD 1.57fF
C13434 a_33338_70226# a_33430_70226# 0.32fF
C13435 a_2124_57979# a_2163_57853# 0.73fF
C13436 a_32426_62194# a_32426_61190# 1.00fF
C13437 a_2959_47113# a_1586_51335# 0.33fF
C13438 a_23390_10496# a_23390_9492# 1.00fF
C13439 a_7265_56053# VDD 1.00fF
C13440 vcm_commonmode a_33338_13874# 0.31fF
C13441 a_49494_58178# m3_49396_58090# 2.78fF
C13442 a_28115_36919# VDD 0.59fF
C13443 a_2021_22325# a_13716_43047# 2.44fF
C13444 a_34251_52263# a_35438_64202# 0.38fF
C13445 a_1586_66567# a_7039_65469# 0.82fF
C13446 a_45478_17524# a_45478_16520# 1.00fF
C13447 a_16955_52047# a_7479_54439# 0.61fF
C13448 vcm_commonmode a_19282_56170# 0.31fF
C13449 a_27535_30503# a_22291_29415# 1.00fF
C13450 a_10515_63143# a_1803_19087# 0.48fF
C13451 a_32426_20536# a_32426_19532# 1.00fF
C13452 a_40458_23548# a_41462_23548# 0.97fF
C13453 a_37919_28111# a_38450_20536# 0.38fF
C13454 a_5595_63125# VDD 1.56fF
C13455 a_49494_56170# a_49494_55166# 1.00fF
C13456 a_17554_30663# VDD 0.45fF
C13457 a_42985_46831# VDD 7.57fF
C13458 a_37446_66210# a_38450_66210# 0.97fF
C13459 vcm_commonmode a_48490_59182# 0.87fF
C13460 ctopn a_18370_19532# 3.58fF
C13461 a_5449_25071# a_5441_27791# 0.35fF
C13462 a_3491_42239# VDD 0.57fF
C13463 a_39389_52271# a_10975_66407# 0.40fF
C13464 a_21371_52263# a_19626_31751# 0.41fF
C13465 a_35676_49525# a_30928_49007# 0.39fF
C13466 a_12641_37684# a_12663_35431# 0.50fF
C13467 a_48398_61190# a_48490_61190# 0.32fF
C13468 a_47486_60186# ctopp 3.58fF
C13469 a_16863_29415# a_4811_34855# 1.75fF
C13470 a_15775_34239# VDD 0.86fF
C13471 vcm_commonmode a_28410_18528# 0.87fF
C13472 a_14287_51175# a_4215_51157# 1.13fF
C13473 a_20286_67214# a_20378_67214# 0.32fF
C13474 vcm_commonmode a_18278_61190# 0.31fF
C13475 ctopn a_46482_22544# 3.58fF
C13476 a_37446_71230# a_37446_70226# 1.00fF
C13477 a_37919_28111# a_38450_12504# 0.38fF
C13478 a_1799_29556# a_1586_21959# 0.55fF
C13479 a_28881_52271# a_29361_51727# 0.48fF
C13480 a_23736_7638# a_12877_14441# 0.41fF
C13481 a_1761_40847# a_13097_37455# 1.29fF
C13482 a_2840_53511# a_5190_59575# 0.63fF
C13483 a_19374_62194# ctopp 3.59fF
C13484 a_41967_31375# a_42466_22544# 0.38fF
C13485 a_9135_27239# a_25744_7638# 4.33fF
C13486 a_49876_41198# a_49876_37608# 0.46fF
C13487 a_14287_51175# a_18370_58178# 0.38fF
C13488 a_23993_37981# VDD 1.00fF
C13489 vcm_commonmode a_19374_55166# 0.84fF
C13490 a_33641_29967# a_37527_29397# 0.51fF
C13491 a_14625_30761# a_20103_30287# 0.38fF
C13492 a_1689_10396# a_1761_25071# 0.84fF
C13493 a_76180_40594# VDD 0.37fF
C13494 a_38557_32143# a_38450_65206# 0.38fF
C13495 a_34780_56398# a_12901_66665# 0.40fF
C13496 a_26402_72234# a_26402_71230# 1.00fF
C13497 vcm_commonmode a_22294_70226# 0.31fF
C13498 a_33430_20536# a_34434_20536# 0.97fF
C13499 a_39362_58178# vcm_commonmode 0.31fF
C13500 vcm_commonmode a_37446_10496# 0.87fF
C13501 a_22386_63198# a_23390_63198# 0.97fF
C13502 ctopn a_42466_14512# 3.59fF
C13503 a_25398_71230# ctopp 3.40fF
C13504 ctopn a_21382_20536# 3.59fF
C13505 a_24959_30503# a_20267_30503# 0.58fF
C13506 a_22294_58178# a_22386_58178# 0.32fF
C13507 a_37919_28111# a_38450_17524# 0.38fF
C13508 a_8295_47388# a_10526_22057# 0.59fF
C13509 a_42466_10496# a_42466_9492# 1.00fF
C13510 a_17274_9858# a_17366_9492# 0.32fF
C13511 a_11067_67279# a_10055_58791# 0.59fF
C13512 a_5024_67885# a_6737_60431# 0.36fF
C13513 a_1761_25071# a_2004_42453# 3.12fF
C13514 a_33430_8488# VDD 0.58fF
C13515 vcm_commonmode a_24394_62194# 0.87fF
C13516 a_33338_16886# a_33430_16520# 0.32fF
C13517 a_34780_56398# a_34434_57174# 0.38fF
C13518 ctopn a_47486_23548# 3.39fF
C13519 a_39389_52271# a_39454_70226# 0.38fF
C13520 a_2944_57960# VDD 0.62fF
C13521 vcm_commonmode a_40366_8854# 0.31fF
C13522 a_19720_7638# a_12895_13967# 0.41fF
C13523 a_40491_27247# a_43470_20536# 0.38fF
C13524 a_41967_31375# a_12727_13353# 0.41fF
C13525 a_1803_20719# a_1761_35407# 0.97fF
C13526 a_6372_38279# a_5631_38127# 0.93fF
C13527 vcm_commonmode a_32426_15516# 0.87fF
C13528 ctopn a_21382_12504# 3.59fF
C13529 a_43470_57174# ctopp 3.58fF
C13530 a_25971_52263# a_12901_58799# 0.40fF
C13531 a_23901_42044# VDD 0.99fF
C13532 a_41427_52263# a_41462_66210# 0.38fF
C13533 a_30764_7638# a_30418_9492# 0.38fF
C13534 a_16902_50639# VDD 0.49fF
C13535 vcm_commonmode a_30418_71230# 0.86fF
C13536 a_29322_72234# a_29414_72234# 0.32fF
C13537 a_5671_21495# a_2143_15271# 0.73fF
C13538 a_31422_21540# a_31422_20536# 1.00fF
C13539 a_49494_61190# VDD 1.12fF
C13540 a_3295_62083# a_1923_54591# 0.33fF
C13541 vcm_commonmode a_42466_11500# 0.87fF
C13542 a_18370_24552# a_18370_23548# 1.00fF
C13543 a_25744_7638# a_12546_22351# 0.41fF
C13544 a_21382_67214# VDD 0.51fF
C13545 a_33430_12504# a_34434_12504# 0.97fF
C13546 a_7281_29423# VDD 1.08fF
C13547 a_41872_29423# a_38115_52263# 1.50fF
C13548 a_1689_10396# a_4578_40455# 1.48fF
C13549 a_39362_67214# a_39454_67214# 0.32fF
C13550 a_39222_48169# a_40458_62194# 0.38fF
C13551 vcm_commonmode a_46482_24552# 0.84fF
C13552 a_28547_51175# a_3339_43023# 0.49fF
C13553 ctopn a_16746_21538# 1.68fF
C13554 vcm_commonmode a_28318_67214# 0.31fF
C13555 a_40491_27247# a_43470_12504# 0.38fF
C13556 a_2143_15271# a_2292_17179# 1.25fF
C13557 a_6831_63303# a_9135_49557# 0.62fF
C13558 a_32772_7638# a_12877_16911# 0.41fF
C13559 a_17222_27247# VDD 1.06fF
C13560 a_3972_25615# a_4417_22671# 0.32fF
C13561 a_39431_37737# VDD 0.62fF
C13562 a_28410_68218# ctopp 3.59fF
C13563 ctopn a_21382_17524# 3.59fF
C13564 a_11719_28023# a_9731_22895# 0.32fF
C13565 a_18370_9492# VDD 0.52fF
C13566 a_1761_47919# a_12473_41781# 1.18fF
C13567 a_2927_39733# a_1761_43567# 0.34fF
C13568 a_3247_20495# a_3987_19623# 1.65fF
C13569 a_13984_43781# a_2021_22325# 0.45fF
C13570 a_25787_28327# a_12355_15055# 0.40fF
C13571 vcm_commonmode a_48490_57174# 0.87fF
C13572 a_25419_50959# a_20267_30503# 0.38fF
C13573 a_34434_16520# VDD 0.51fF
C13574 a_17507_52047# a_12516_7093# 0.40fF
C13575 a_11251_59879# a_11067_46823# 1.10fF
C13576 a_36629_27791# a_36442_14512# 0.38fF
C13577 a_25306_7850# a_25398_7484# 0.32fF
C13578 vcm_commonmode a_25306_9858# 0.31fF
C13579 m3_17268_72146# VDD 0.42fF
C13580 a_35438_24552# m3_35340_24414# 2.81fF
C13581 a_41462_63198# a_42466_63198# 0.97fF
C13582 a_12355_65103# a_11251_59879# 12.67fF
C13583 vcm_commonmode a_41370_16886# 0.31fF
C13584 a_41967_31375# a_10515_23975# 0.41fF
C13585 a_12473_41781# a_12641_42036# 0.83fF
C13586 a_30326_72234# VDD 0.62fF
C13587 vcm_commonmode a_23736_7638# 10.35fF
C13588 a_33864_28111# a_12727_13353# 0.41fF
C13589 a_40675_27791# a_12985_16367# 0.41fF
C13590 a_28410_21540# a_29414_21540# 0.97fF
C13591 a_40491_27247# a_43470_17524# 0.38fF
C13592 a_36350_9858# a_36442_9492# 0.32fF
C13593 a_19282_64202# a_19374_64202# 0.32fF
C13594 a_13143_29575# a_13239_29575# 1.14fF
C13595 a_12549_44212# a_12473_42869# 2.55fF
C13596 a_26402_7484# VDD 1.38fF
C13597 a_46482_58178# a_47486_58178# 0.97fF
C13598 a_1761_49007# a_6863_42692# 1.66fF
C13599 a_22843_29415# a_20267_30503# 7.67fF
C13600 vcm_commonmode a_33430_68218# 0.87fF
C13601 a_35438_59182# a_36442_59182# 0.97fF
C13602 a_6831_63303# a_2595_47653# 0.40fF
C13603 a_16362_22544# a_16746_22542# 2.28fF
C13604 a_40491_27247# a_12895_13967# 0.41fF
C13605 a_20378_64202# VDD 0.51fF
C13606 a_18979_30287# a_28757_27247# 1.47fF
C13607 a_49876_37608# a_49750_39288# 0.40fF
C13608 a_28410_56170# ctopp 3.40fF
C13609 a_1644_70197# VDD 0.31fF
C13610 a_25300_38567# VDD 1.85fF
C13611 ctopn a_22386_18528# 3.59fF
C13612 a_2787_32679# a_1689_10396# 0.44fF
C13613 vcm_commonmode a_27314_64202# 0.31fF
C13614 a_33430_17524# a_34434_17524# 0.97fF
C13615 a_33826_50075# VDD 0.63fF
C13616 a_39673_28111# a_40458_15516# 0.38fF
C13617 a_20378_60186# a_21382_60186# 0.97fF
C13618 a_4798_23759# VDD 1.42fF
C13619 a_37446_24552# a_37446_23548# 1.00fF
C13620 a_22386_12504# a_22386_11500# 1.00fF
C13621 a_27752_7638# a_26748_7638# 0.31fF
C13622 a_15661_29199# a_15681_27497# 0.65fF
C13623 a_1761_22895# a_33155_40191# 0.34fF
C13624 a_2021_17973# VDD 8.21fF
C13625 a_26748_7638# a_26402_10496# 0.38fF
C13626 a_2177_53359# VDD 0.32fF
C13627 a_42709_29199# a_12727_13353# 0.40fF
C13628 a_37919_28111# a_12877_16911# 0.41fF
C13629 a_23736_7638# a_23390_14512# 0.38fF
C13630 a_2605_60975# VDD 0.48fF
C13631 vcm_commonmode a_47486_13508# 0.87fF
C13632 a_27406_61190# ctopp 3.59fF
C13633 ctopn a_31422_10496# 3.59fF
C13634 a_33864_28111# a_10515_23975# 0.40fF
C13635 a_29760_7638# a_29414_24552# 0.46fF
C13636 a_29414_69222# VDD 0.51fF
C13637 a_3668_56311# a_5336_54965# 0.33fF
C13638 a_28547_51175# a_12257_56623# 0.40fF
C13639 vcm_commonmode a_33430_56170# 0.87fF
C13640 a_1591_14741# VDD 0.40fF
C13641 vcm_commonmode a_36350_69222# 0.31fF
C13642 a_36442_22544# VDD 0.51fF
C13643 a_44382_7850# a_44474_7484# 0.32fF
C13644 vcm_commonmode a_16362_8488# 4.46fF
C13645 a_27406_65206# VDD 0.51fF
C13646 a_15290_30761# VDD 0.33fF
C13647 a_32327_40191# a_24029_39355# 1.89fF
C13648 a_23395_52047# a_10515_22671# 0.40fF
C13649 vcm_commonmode a_43378_22910# 0.31fF
C13650 a_31422_70226# ctopp 3.58fF
C13651 a_25313_31599# a_23736_7638# 0.38fF
C13652 a_1761_50639# a_19629_39631# 0.61fF
C13653 a_22411_42359# VDD 0.60fF
C13654 vcm_commonmode a_34342_65206# 0.31fF
C13655 a_28318_69222# a_28410_69222# 0.32fF
C13656 a_9135_27239# a_21382_9492# 0.38fF
C13657 a_34434_18528# a_34434_17524# 1.00fF
C13658 a_1591_16917# a_1757_16917# 0.62fF
C13659 a_13097_36367# a_12889_35537# 0.66fF
C13660 a_8295_47388# a_4674_40277# 0.50fF
C13661 a_19720_55394# a_17599_52263# 0.37fF
C13662 a_16955_52047# a_17507_52047# 0.68fF
C13663 a_47486_21540# a_48490_21540# 0.97fF
C13664 a_9503_26151# a_12727_13353# 0.41fF
C13665 a_16270_24918# VDD 0.46fF
C13666 a_10515_22671# a_8491_27023# 1.01fF
C13667 a_36629_27791# a_11067_21583# 0.41fF
C13668 a_38358_64202# a_38450_64202# 0.32fF
C13669 ctopn a_26402_15516# 3.59fF
C13670 a_1761_4399# VDD 0.62fF
C13671 vcm_commonmode a_32426_61190# 0.87fF
C13672 a_32426_14512# VDD 0.51fF
C13673 a_7407_46529# VDD 0.47fF
C13674 a_40050_48463# a_45478_69222# 0.38fF
C13675 a_27314_55166# VDD 0.35fF
C13676 a_35346_22910# a_35438_22544# 0.32fF
C13677 a_24394_10496# a_25398_10496# 0.97fF
C13678 vcm_commonmode a_39362_14878# 0.31fF
C13679 ctopn a_36442_11500# 3.59fF
C13680 a_42709_29199# a_10515_23975# 0.40fF
C13681 a_7841_12167# a_9275_15253# 0.34fF
C13682 a_26310_65206# a_26402_65206# 0.32fF
C13683 a_35438_14512# a_35438_13508# 1.00fF
C13684 vcm_commonmode a_18278_20902# 0.31fF
C13685 vcm_commonmode a_33338_55166# 0.30fF
C13686 a_24423_40229# VDD 1.08fF
C13687 vcm_commonmode a_36442_70226# 0.87fF
C13688 a_39454_60186# a_40458_60186# 0.97fF
C13689 a_37446_23548# VDD 0.52fF
C13690 a_20378_58178# ctopp 3.59fF
C13691 a_17274_23914# a_17366_23548# 0.32fF
C13692 a_34434_66210# VDD 0.51fF
C13693 a_27535_30503# a_27797_29423# 0.39fF
C13694 a_41462_12504# a_41462_11500# 1.00fF
C13695 vcm_commonmode a_17366_16520# 1.82fF
C13696 vcm_commonmode a_44382_23914# 0.31fF
C13697 a_28410_70226# a_28410_69222# 1.00fF
C13698 a_41872_29423# a_12983_63151# 0.40fF
C13699 vcm_commonmode a_41370_66210# 0.31fF
C13700 a_34434_18528# a_35438_18528# 0.97fF
C13701 a_37307_51339# a_37423_51335# 0.37fF
C13702 a_46482_19532# VDD 0.51fF
C13703 a_27167_52271# VDD 0.35fF
C13704 vcm_commonmode a_17366_72234# 0.69fF
C13705 a_2686_70223# a_6921_72943# 0.42fF
C13706 vcm_commonmode a_18278_12870# 0.31fF
C13707 a_8491_57487# a_8132_53511# 0.87fF
C13708 a_9503_26151# a_10515_23975# 0.41fF
C13709 a_3040_68425# VDD 0.32fF
C13710 a_11067_13095# a_11067_63143# 1.48fF
C13711 a_11803_64239# a_11759_63927# 0.36fF
C13712 a_37446_67214# ctopp 3.59fF
C13713 a_12621_44099# a_12663_40871# 0.60fF
C13714 a_40050_48463# a_12981_62313# 0.40fF
C13715 a_26310_19898# a_26402_19532# 0.32fF
C13716 a_7050_53333# a_4215_51157# 0.31fF
C13717 a_7567_64391# VDD 0.36fF
C13718 a_27406_11500# a_27406_10496# 1.00fF
C13719 a_25971_29967# VDD 0.44fF
C13720 a_25971_52263# a_18703_29199# 0.82fF
C13721 a_19629_39631# a_23789_39100# 0.39fF
C13722 a_25971_52263# a_30418_59182# 0.38fF
C13723 vcm_commonmode a_25398_58178# 0.87fF
C13724 a_31330_14878# a_31422_14512# 0.32fF
C13725 a_11803_55311# a_12355_65103# 1.74fF
C13726 a_47394_69222# a_47486_69222# 0.32fF
C13727 a_39673_28111# a_12877_14441# 0.41fF
C13728 a_12447_29199# a_28817_29111# 0.49fF
C13729 a_2411_19605# VDD 4.10fF
C13730 a_25398_55166# a_26402_55166# 0.97fF
C13731 vcm_commonmode a_18278_17890# 0.31fF
C13732 a_19374_15516# a_20378_15516# 0.97fF
C13733 a_9367_29397# a_9405_31599# 0.42fF
C13734 a_1761_22895# VDD 9.24fF
C13735 a_43362_28879# a_12727_67753# 0.40fF
C13736 vcm_commonmode a_42466_67214# 0.87fF
C13737 a_49494_20536# VDD 1.12fF
C13738 a_12683_51329# a_13445_50639# 0.50fF
C13739 a_10055_58791# a_1586_18695# 0.32fF
C13740 a_8575_74853# a_6224_73095# 0.48fF
C13741 a_38450_63198# VDD 0.57fF
C13742 a_43470_10496# a_44474_10496# 0.97fF
C13743 a_45386_65206# a_45478_65206# 0.32fF
C13744 a_31768_55394# a_31422_64202# 0.38fF
C13745 vcm_commonmode a_45386_63198# 0.31fF
C13746 a_2235_30503# a_7939_30503# 0.95fF
C13747 a_16863_29415# a_20635_29415# 1.04fF
C13748 a_17366_71230# a_18370_71230# 0.97fF
C13749 a_28547_51175# a_8531_70543# 1.99fF
C13750 a_32426_59182# VDD 0.51fF
C13751 vcm_commonmode a_39454_9492# 0.87fF
C13752 a_36350_23914# a_36442_23548# 0.32fF
C13753 a_10975_65327# VDD 0.48fF
C13754 a_13643_28327# a_32970_31145# 0.53fF
C13755 a_21187_29415# a_32823_29397# 0.41fF
C13756 a_29414_11500# a_30418_11500# 0.97fF
C13757 a_36442_64202# ctopp 3.59fF
C13758 ctopn a_41462_13508# 3.59fF
C13759 a_41427_52263# VDD 10.59fF
C13760 a_33338_66210# a_33430_66210# 0.32fF
C13761 vcm_commonmode a_39362_59182# 0.31fF
C13762 a_4429_14191# a_4812_13879# 1.56fF
C13763 vcm_commonmode a_19374_22544# 0.87fF
C13764 a_11719_28023# a_10506_29967# 0.38fF
C13765 vcm_commonmode m3_16264_56082# 3.05fF
C13766 a_49494_12504# VDD 1.12fF
C13767 a_28547_51175# a_10975_66407# 0.40fF
C13768 a_16746_69224# a_16362_69222# 2.28fF
C13769 a_47486_70226# a_47486_69222# 1.00fF
C13770 a_1761_37039# a_15968_36061# 2.06fF
C13771 a_30757_37455# a_32327_35839# 0.42fF
C13772 a_11711_50645# a_11877_50645# 0.42fF
C13773 a_7073_51433# VDD 0.41fF
C13774 vcm_commonmode a_43267_31055# 10.10fF
C13775 a_5309_25853# VDD 0.51fF
C13776 a_9955_20969# a_7187_23439# 0.30fF
C13777 a_33430_24552# a_34434_24552# 0.97fF
C13778 a_16510_8760# a_12985_16367# 1.08fF
C13779 a_17366_56170# m3_17268_56082# 2.77fF
C13780 a_25447_34743# VDD 0.63fF
C13781 vcm_commonmode a_19282_18894# 0.31fF
C13782 a_20359_29199# a_18979_30287# 1.20fF
C13783 a_45386_19898# a_45478_19532# 0.32fF
C13784 a_44474_21540# VDD 0.51fF
C13785 vcm_commonmode a_47486_7484# 0.69fF
C13786 a_30418_62194# a_31422_62194# 0.97fF
C13787 a_23928_28585# VDD 0.82fF
C13788 a_46482_11500# a_46482_10496# 1.00fF
C13789 a_13349_37973# a_1761_39215# 0.60fF
C13790 a_45478_69222# ctopp 3.59fF
C13791 a_3339_43023# a_12621_36091# 0.36fF
C13792 a_21382_10496# VDD 0.51fF
C13793 a_24331_40767# VDD 1.06fF
C13794 a_34780_56398# a_34434_65206# 0.38fF
C13795 vcm_commonmode a_41462_64202# 0.87fF
C13796 a_2143_15271# a_3327_9308# 0.35fF
C13797 a_1591_49557# a_2292_43291# 0.33fF
C13798 a_49494_17524# VDD 1.10fF
C13799 a_10391_49855# VDD 0.62fF
C13800 a_23395_52047# a_12901_66665# 0.40fF
C13801 a_22386_72234# a_22386_71230# 1.00fF
C13802 a_8491_27023# a_18370_15516# 0.38fF
C13803 a_25744_7638# a_25398_15516# 0.38fF
C13804 a_29322_20902# a_29414_20536# 0.32fF
C13805 a_36442_60186# VDD 0.51fF
C13806 a_12447_29199# a_37699_27221# 0.33fF
C13807 a_43470_55166# a_44474_55166# 0.97fF
C13808 vcm_commonmode a_28318_10862# 0.31fF
C13809 a_18278_63198# a_18370_63198# 0.32fF
C13810 a_20881_28111# VDD 2.03fF
C13811 a_43470_65206# ctopp 3.59fF
C13812 a_35438_57174# a_36442_57174# 0.97fF
C13813 vcm_commonmode a_43378_60186# 0.31fF
C13814 a_38450_15516# a_39454_15516# 0.97fF
C13815 VDD start_conversion_in 1.23fF
C13816 vcm_commonmode a_20378_23548# 0.87fF
C13817 a_2292_43291# a_1761_43567# 0.40fF
C13818 a_17803_44265# VDD 0.59fF
C13819 vcm_commonmode a_17366_66210# 1.83fF
C13820 a_10503_52828# VDD 4.77fF
C13821 a_4758_45369# VDD 9.04fF
C13822 a_31263_27221# VDD 0.46fF
C13823 a_41999_36367# VDD 0.47fF
C13824 vcm_commonmode a_29414_19532# 0.87fF
C13825 a_38450_58178# a_38450_59182# 1.00fF
C13826 vcm_commonmode a_39673_28111# 10.35fF
C13827 a_25971_52263# a_30418_57174# 0.38fF
C13828 a_16746_15514# VDD 33.20fF
C13829 VDD config_2_in[8] 0.79fF
C13830 a_34251_52263# a_35438_70226# 0.38fF
C13831 a_36442_71230# a_37446_71230# 0.97fF
C13832 a_7571_29199# a_2787_30503# 0.36fF
C13833 a_48490_11500# a_49494_11500# 0.97fF
C13834 vcm_commonmode a_23298_15882# 0.31fF
C13835 a_12981_62313# ctopp 3.23fF
C13836 a_1586_21959# a_1591_23445# 0.80fF
C13837 a_42985_46831# a_48490_60186# 0.38fF
C13838 a_18611_52047# a_12901_58799# 0.40fF
C13839 a_12985_19087# a_12947_8725# 23.40fF
C13840 a_12585_39069# VDD 1.06fF
C13841 a_26402_11500# VDD 0.51fF
C13842 vcm_commonmode a_48490_65206# 0.87fF
C13843 a_36613_48169# a_37446_66210# 0.38fF
C13844 vcm_commonmode a_21290_71230# 0.31fF
C13845 a_12947_8725# a_16746_8486# 2.25fF
C13846 a_30418_24552# VDD 0.60fF
C13847 vcm_commonmode a_33338_11866# 0.31fF
C13848 ctopn a_48490_8488# 3.24fF
C13849 a_4425_32687# VDD 0.59fF
C13850 a_29322_12870# a_29414_12504# 0.32fF
C13851 a_36717_47375# a_36442_62194# 0.38fF
C13852 vcm_commonmode a_37354_24918# 0.31fF
C13853 a_24394_59182# a_24394_58178# 1.00fF
C13854 a_40458_55166# VDD 0.60fF
C13855 a_7295_44647# a_23736_7638# 2.54fF
C13856 a_32426_57174# VDD 0.51fF
C13857 a_11067_23759# a_12985_19087# 0.36fF
C13858 a_12516_7093# a_10515_22671# 0.43fF
C13859 vcm_commonmode a_32426_20536# 0.87fF
C13860 vcm_commonmode a_47394_55166# 0.30fF
C13861 a_1761_47919# a_27245_41829# 0.31fF
C13862 a_20378_68218# a_21382_68218# 0.97fF
C13863 a_21371_52263# a_12355_15055# 0.44fF
C13864 vcm_commonmode a_21382_63198# 0.92fF
C13865 vcm_commonmode a_39362_57174# 0.31fF
C13866 a_4811_34855# a_2235_30503# 0.99fF
C13867 a_27535_30503# a_12907_27023# 0.31fF
C13868 a_11067_46823# a_22015_28111# 1.00fF
C13869 a_48398_20902# a_48490_20536# 0.32fF
C13870 a_23736_7638# a_12899_11471# 0.41fF
C13871 a_28410_24552# m3_28312_24414# 2.81fF
C13872 a_37354_63198# a_37446_63198# 0.32fF
C13873 a_6467_55527# a_7479_54439# 0.52fF
C13874 a_28410_57174# a_28410_56170# 1.00fF
C13875 a_23298_72234# VDD 0.61fF
C13876 a_1761_52815# a_4123_37013# 1.16fF
C13877 a_37939_43455# VDD 0.60fF
C13878 a_13925_51727# VDD 0.91fF
C13879 a_6559_59879# a_18501_50645# 0.60fF
C13880 a_24302_21906# a_24394_21540# 0.32fF
C13881 a_46482_62194# VDD 0.51fF
C13882 a_12641_37684# a_27600_36165# 0.30fF
C13883 a_2235_30503# config_2_in[0] 0.44fF
C13884 a_9695_54965# VDD 0.46fF
C13885 vcm_commonmode a_32426_12504# 0.87fF
C13886 ctopn a_33430_9492# 3.58fF
C13887 a_2840_66103# a_4215_51157# 0.76fF
C13888 a_17366_68218# VDD 0.57fF
C13889 a_18627_35327# VDD 0.89fF
C13890 a_2021_17973# a_12663_40871# 1.67fF
C13891 a_17274_7850# VDD 0.64fF
C13892 a_3143_66972# a_2840_53511# 1.80fF
C13893 a_3024_67191# a_7213_62215# 0.39fF
C13894 vcm_commonmode a_24302_68218# 0.31fF
C13895 a_31330_59182# a_31422_59182# 0.32fF
C13896 a_1761_52815# a_2872_44111# 1.28fF
C13897 a_8636_63669# VDD 0.32fF
C13898 a_51330_39932# a_51422_39932# 0.44fF
C13899 a_1923_59583# a_1823_63677# 0.31fF
C13900 vcm_commonmode a_27406_21540# 0.87fF
C13901 a_43470_72234# m3_43372_72146# 2.80fF
C13902 a_25987_41317# VDD 0.97fF
C13903 a_29322_17890# a_29414_17524# 0.32fF
C13904 vcm_commonmode a_45478_58178# 0.87fF
C13905 a_4191_33449# VDD 9.17fF
C13906 a_13183_52047# a_17366_71230# 0.38fF
C13907 a_16746_60188# a_12727_58255# 0.41fF
C13908 a_48490_59182# ctopp 3.43fF
C13909 a_10515_23975# a_12947_23413# 23.33fF
C13910 a_35438_64202# a_35438_63198# 1.23fF
C13911 a_31964_30485# VDD 0.74fF
C13912 a_48398_12870# a_48490_12504# 0.32fF
C13913 vcm_commonmode a_32426_17524# 0.87fF
C13914 a_12473_42869# a_13576_42589# 0.40fF
C13915 a_13067_38517# a_33764_41831# 0.52fF
C13916 vcm_commonmode a_19374_60186# 0.87fF
C13917 a_31422_13508# VDD 0.51fF
C13918 a_1761_52815# a_1761_40847# 0.53fF
C13919 a_38450_58178# a_38450_57174# 1.00fF
C13920 a_31004_44869# VDD 1.78fF
C13921 a_6738_19783# VDD 1.44fF
C13922 a_4240_53083# VDD 0.57fF
C13923 a_27406_22544# a_27406_21540# 1.00fF
C13924 a_11067_63143# a_10515_22671# 0.96fF
C13925 a_10515_63143# a_11251_59879# 0.91fF
C13926 a_17366_56170# VDD 0.58fF
C13927 vcm_commonmode a_38358_13874# 0.31fF
C13928 a_34434_13508# a_35438_13508# 0.97fF
C13929 a_40895_36919# VDD 0.64fF
C13930 a_3339_30503# a_25462_27497# 0.32fF
C13931 a_39454_68218# a_40458_68218# 0.97fF
C13932 vcm_commonmode a_24302_56170# 0.31fF
C13933 a_21371_50959# a_12257_56623# 0.40fF
C13934 a_5639_15279# VDD 0.39fF
C13935 a_32772_7638# a_12895_13967# 0.41fF
C13936 a_39673_28111# a_40458_20536# 0.38fF
C13937 a_23395_52047# a_19807_28111# 1.04fF
C13938 a_12985_25615# a_10964_25615# 0.32fF
C13939 a_20378_56170# a_21382_56170# 0.97fF
C13940 a_47486_57174# a_47486_56170# 1.00fF
C13941 a_16955_52047# a_10515_22671# 0.40fF
C13942 ctopn a_23390_19532# 3.59fF
C13943 a_43362_28879# a_41842_27221# 0.68fF
C13944 a_25744_7638# a_12985_16367# 0.41fF
C13945 a_43378_21906# a_43470_21540# 0.32fF
C13946 a_12981_59343# VDD 7.05fF
C13947 a_20635_29415# a_40491_27247# 0.78fF
C13948 a_8583_33551# a_19807_28111# 0.65fF
C13949 a_24394_58178# a_24394_57174# 1.00fF
C13950 a_36629_27791# a_12546_22351# 0.41fF
C13951 a_18627_34239# VDD 0.72fF
C13952 vcm_commonmode a_33430_18528# 0.87fF
C13953 vcm_commonmode a_23298_61190# 0.31fF
C13954 a_31422_16520# a_31422_15516# 1.00fF
C13955 a_13183_52047# a_12659_54965# 0.38fF
C13956 a_12447_29199# VDD 9.90fF
C13957 a_41427_52263# a_41462_69222# 0.38fF
C13958 a_39673_28111# a_40458_12504# 0.38fF
C13959 a_12895_13967# a_16362_18528# 19.89fF
C13960 a_18611_52047# a_16510_8760# 2.01fF
C13961 a_18602_55312# VDD 0.45fF
C13962 a_49402_64202# VDD 0.32fF
C13963 a_20286_10862# a_20378_10496# 0.32fF
C13964 a_8123_56399# VDD 7.46fF
C13965 a_24394_62194# ctopp 3.59fF
C13966 a_20378_70226# VDD 0.51fF
C13967 a_37446_58178# VDD 0.51fF
C13968 vcm_commonmode a_24394_55166# 0.84fF
C13969 a_2952_46805# a_1761_43567# 0.31fF
C13970 a_3305_38671# VDD 4.51fF
C13971 a_1586_66567# a_2840_66103# 0.34fF
C13972 a_48398_17890# a_48490_17524# 0.32fF
C13973 a_5529_16367# VDD 0.65fF
C13974 a_30525_49551# VDD 0.83fF
C13975 vcm_commonmode a_27314_70226# 0.31fF
C13976 a_35346_60186# a_35438_60186# 0.32fF
C13977 vcm_commonmode a_42466_10496# 0.87fF
C13978 a_37919_28111# a_38450_21540# 0.38fF
C13979 a_27752_7638# a_12985_19087# 0.41fF
C13980 a_8491_27023# a_7377_18012# 0.90fF
C13981 ctopn a_47486_14512# 3.58fF
C13982 a_7707_70741# VDD 2.80fF
C13983 a_30418_71230# ctopp 3.40fF
C13984 ctopn a_26402_20536# 3.59fF
C13985 a_2592_43023# VDD 0.44fF
C13986 a_36717_47375# a_12983_63151# 0.40fF
C13987 a_30326_18894# a_30418_18528# 0.32fF
C13988 a_3751_72373# a_6327_72917# 0.41fF
C13989 a_2124_73211# a_2163_73085# 0.76fF
C13990 a_46482_22544# a_46482_21540# 1.00fF
C13991 a_39673_28111# a_40458_17524# 0.38fF
C13992 a_19374_61190# a_20378_61190# 0.97fF
C13993 a_1853_27247# VDD 0.43fF
C13994 a_14258_34191# VDD 0.69fF
C13995 a_38450_8488# VDD 0.58fF
C13996 a_38557_32143# a_12981_62313# 0.40fF
C13997 a_25398_68218# a_25398_67214# 1.00fF
C13998 vcm_commonmode a_29414_62194# 0.87fF
C13999 a_2606_41079# a_6863_42692# 0.48fF
C14000 a_11067_46823# a_22291_29415# 6.57fF
C14001 a_26917_47919# VDD 0.50fF
C14002 vcm_commonmode a_11067_67279# 6.37fF
C14003 a_12901_66665# a_12516_7093# 24.86fF
C14004 a_49494_17524# m3_49396_17386# 2.78fF
C14005 a_7050_53333# a_15557_52245# 0.30fF
C14006 vcm_commonmode a_45386_8854# 0.31fF
C14007 a_37919_28111# a_12895_13967# 0.41fF
C14008 a_12024_30199# VDD 0.43fF
C14009 vcm_commonmode a_37446_15516# 0.87fF
C14010 ctopn a_26402_12504# 3.59fF
C14011 a_48490_57174# ctopp 3.43fF
C14012 a_39454_56170# a_40458_56170# 0.97fF
C14013 a_21371_52263# a_26402_59182# 0.38fF
C14014 a_10975_66407# a_1586_21959# 1.22fF
C14015 a_26433_39631# VDD 2.88fF
C14016 a_7649_17455# VDD 0.44fF
C14017 vcm_commonmode a_35438_71230# 0.86fF
C14018 a_31768_55394# a_31422_72234# 0.34fF
C14019 a_10515_63143# a_8566_39215# 2.06fF
C14020 a_21290_55166# a_21382_55166# 0.32fF
C14021 a_22386_8488# a_23390_8488# 0.97fF
C14022 vcm_commonmode a_47486_11500# 0.87fF
C14023 a_29760_7638# a_11067_21583# 0.41fF
C14024 a_26402_67214# VDD 0.51fF
C14025 a_8132_53511# a_7479_54439# 1.73fF
C14026 a_4351_67279# a_6831_63303# 0.38fF
C14027 ctopn a_21382_21540# 3.59fF
C14028 a_1586_45431# a_1757_45205# 0.60fF
C14029 vcm_commonmode a_33338_67214# 0.31fF
C14030 a_39222_48169# a_12727_67753# 0.40fF
C14031 a_23390_70226# a_24394_70226# 0.97fF
C14032 a_35438_19532# a_35438_18528# 1.00fF
C14033 a_21371_52263# a_7939_30503# 1.78fF
C14034 a_40458_58178# a_41462_58178# 0.97fF
C14035 a_5441_72399# a_5475_74895# 0.35fF
C14036 a_17712_7638# a_12899_10927# 0.40fF
C14037 a_2411_19605# a_1591_19631# 0.33fF
C14038 a_20635_29415# a_12899_3311# 1.76fF
C14039 a_16863_29415# a_12899_2767# 1.16fF
C14040 a_39362_10862# a_39454_10496# 0.32fF
C14041 a_5823_28585# VDD 0.30fF
C14042 a_33430_68218# ctopp 3.59fF
C14043 ctopn a_26402_17524# 3.59fF
C14044 a_23390_9492# VDD 0.51fF
C14045 a_28931_39679# VDD 0.97fF
C14046 a_23395_52047# a_27406_64202# 0.38fF
C14047 a_5915_35943# a_12935_31287# 0.32fF
C14048 a_39454_16520# VDD 0.51fF
C14049 a_32227_48169# VDD 0.70fF
C14050 a_4298_58951# a_2606_41079# 0.54fF
C14051 a_21382_60186# a_21382_59182# 1.00fF
C14052 vcm_commonmode a_30326_9858# 0.31fF
C14053 a_40491_27247# a_43470_21540# 0.38fF
C14054 a_25306_11866# a_25398_11500# 0.32fF
C14055 vcm_commonmode a_46390_16886# 0.31fF
C14056 a_34780_56398# VDD 6.52fF
C14057 a_30418_15516# a_30418_14512# 1.00fF
C14058 a_35815_31751# a_32823_29397# 0.79fF
C14059 a_4495_35925# a_7461_27247# 0.39fF
C14060 a_7862_34025# a_23195_29967# 0.37fF
C14061 vcm_commonmode m3_16264_70138# 3.20fF
C14062 a_8958_65961# a_9914_68279# 0.37fF
C14063 a_21371_50959# a_10975_66407# 0.40fF
C14064 a_49402_18894# a_49494_18528# 0.32fF
C14065 a_11067_47695# a_17449_46831# 0.42fF
C14066 a_37534_51701# VDD 0.87fF
C14067 vcm_commonmode a_39389_52271# 10.02fF
C14068 a_15607_46805# a_26748_7638# 1.49fF
C14069 a_38450_61190# a_39454_61190# 0.97fF
C14070 a_29322_24918# a_29414_24552# 0.32fF
C14071 a_3063_34319# VDD 0.42fF
C14072 a_31422_7484# VDD 1.23fF
C14073 a_44474_68218# a_44474_67214# 1.00fF
C14074 vcm_commonmode a_38450_68218# 0.87fF
C14075 a_41261_28335# a_12901_66959# 0.40fF
C14076 a_8491_27023# a_12985_19087# 0.41fF
C14077 a_25398_64202# VDD 0.51fF
C14078 a_20267_30503# a_14646_29423# 0.77fF
C14079 a_26310_62194# a_26402_62194# 0.32fF
C14080 a_33430_56170# ctopp 3.51fF
C14081 a_32795_38591# VDD 0.83fF
C14082 ctopn a_27406_18528# 3.59fF
C14083 a_29414_69222# a_29414_68218# 1.00fF
C14084 a_25971_52263# a_30418_65206# 0.38fF
C14085 vcm_commonmode a_32334_64202# 0.31fF
C14086 a_2473_34293# a_1761_34319# 0.36fF
C14087 a_1586_40455# VDD 5.06fF
C14088 a_16955_52047# a_12901_66665# 0.40fF
C14089 a_18370_72234# a_18370_71230# 1.00fF
C14090 a_40050_48463# a_43267_31055# 2.39fF
C14091 a_39362_55166# a_39454_55166# 0.32fF
C14092 a_9971_23439# VDD 0.39fF
C14093 a_41462_8488# a_42466_8488# 0.97fF
C14094 a_19374_8488# a_19374_7484# 1.00fF
C14095 a_1849_31599# VDD 0.51fF
C14096 a_31330_57174# a_31422_57174# 0.32fF
C14097 a_34342_15882# a_34434_15516# 0.32fF
C14098 a_11619_56615# a_12024_30199# 0.44fF
C14099 a_2663_43541# VDD 0.43fF
C14100 a_43267_31055# a_46482_68218# 0.38fF
C14101 a_42466_70226# a_43470_70226# 0.97fF
C14102 a_39673_28111# a_12899_11471# 0.41fF
C14103 a_3016_60949# VDD 4.24fF
C14104 a_20359_27791# VDD 0.49fF
C14105 a_32426_61190# ctopp 3.59fF
C14106 ctopn a_36442_10496# 3.59fF
C14107 a_42709_29199# a_48490_23548# 0.42fF
C14108 a_32951_27247# a_33430_24552# 0.42fF
C14109 a_34434_69222# VDD 0.51fF
C14110 vcm_commonmode a_20286_19898# 0.31fF
C14111 a_12947_8725# VDD 4.18fF
C14112 a_23390_16520# a_24394_16520# 0.97fF
C14113 vcm_commonmode a_38450_56170# 0.87fF
C14114 a_21371_52263# a_26402_57174# 0.38fF
C14115 a_9379_15039# VDD 0.38fF
C14116 vcm_commonmode a_41370_69222# 0.31fF
C14117 a_32334_71230# a_32426_71230# 0.32fF
C14118 a_31768_55394# a_31422_70226# 0.38fF
C14119 a_40458_60186# a_40458_59182# 1.00fF
C14120 a_41462_22544# VDD 0.51fF
C14121 vcm_commonmode a_21382_8488# 0.86fF
C14122 a_8491_27023# a_18370_20536# 0.38fF
C14123 a_25744_7638# a_25398_20536# 0.38fF
C14124 a_32426_65206# VDD 0.51fF
C14125 a_6835_46823# a_17039_51157# 1.94fF
C14126 a_29414_63198# a_29414_62194# 1.00fF
C14127 a_44382_11866# a_44474_11500# 0.32fF
C14128 a_10055_58791# a_1586_21959# 0.38fF
C14129 a_39299_48783# a_44474_60186# 0.38fF
C14130 a_49494_15516# a_49494_14512# 1.00fF
C14131 vcm_commonmode a_48398_22910# 0.31fF
C14132 a_36442_70226# ctopp 3.58fF
C14133 vcm_commonmode m3_16264_17386# 3.21fF
C14134 a_37885_42333# VDD 0.88fF
C14135 a_25787_28327# a_33430_66210# 0.38fF
C14136 vcm_commonmode a_39362_65206# 0.31fF
C14137 a_43267_31055# a_12355_65103# 0.40fF
C14138 a_32772_7638# a_32426_8488# 0.38fF
C14139 a_1761_30511# a_1761_31055# 1.76fF
C14140 a_22294_72234# a_22386_72234# 0.32fF
C14141 a_26748_7638# a_26402_15516# 0.38fF
C14142 a_34434_9492# a_34434_8488# 1.00fF
C14143 a_21290_24918# VDD 0.36fF
C14144 a_39223_32463# a_39454_18528# 0.38fF
C14145 a_12355_15055# a_6831_63303# 1.96fF
C14146 a_11067_23759# VDD 26.03fF
C14147 ctopn a_31422_15516# 3.59fF
C14148 a_9529_28335# a_14471_28585# 0.55fF
C14149 a_2787_32679# a_4578_40455# 0.55fF
C14150 a_12663_40871# a_37939_43455# 0.43fF
C14151 m2_15446_73620# VDD 0.60fF
C14152 vcm_commonmode a_37446_61190# 0.87fF
C14153 a_29414_67214# a_30418_67214# 0.97fF
C14154 a_28547_51175# a_32426_62194# 0.38fF
C14155 a_43267_31055# a_46482_56170# 0.38fF
C14156 a_37446_14512# VDD 0.51fF
C14157 a_8491_27023# a_18370_12504# 0.38fF
C14158 a_25744_7638# a_25398_12504# 0.38fF
C14159 a_21371_52263# a_4811_34855# 0.53fF
C14160 a_16362_20536# VDD 2.47fF
C14161 a_11067_47695# VDD 11.35fF
C14162 a_2944_63400# VDD 0.48fF
C14163 a_45386_62194# a_45478_62194# 0.32fF
C14164 a_6467_55527# a_6559_59879# 0.53fF
C14165 vcm_commonmode a_44382_14878# 0.31fF
C14166 ctopn a_41462_11500# 3.59fF
C14167 a_43269_29967# a_47486_23548# 0.38fF
C14168 vcm_commonmode a_23298_20902# 0.31fF
C14169 a_31243_40183# VDD 0.65fF
C14170 a_48490_69222# a_48490_68218# 1.00fF
C14171 a_19720_55394# a_12355_15055# 0.40fF
C14172 a_16746_68220# a_12727_67753# 0.41fF
C14173 a_1761_49007# VDD 7.56fF
C14174 vcm_commonmode a_41462_70226# 0.87fF
C14175 a_7571_29199# a_10472_26159# 0.61fF
C14176 a_42466_23548# VDD 0.52fF
C14177 a_38450_8488# a_38450_7484# 1.00fF
C14178 a_25398_58178# ctopp 3.59fF
C14179 a_39454_66210# VDD 0.51fF
C14180 VDD config_1_in[10] 1.38fF
C14181 a_21382_24552# m3_21284_24414# 2.81fF
C14182 vcm_commonmode a_22386_16520# 0.87fF
C14183 a_12899_2767# a_19720_7638# 2.44fF
C14184 vcm_commonmode a_49402_23914# 0.30fF
C14185 a_16362_12504# VDD 2.47fF
C14186 vcm_commonmode a_46390_66210# 0.31fF
C14187 a_31422_58178# a_32426_58178# 0.97fF
C14188 a_4242_35407# a_4495_35925# 0.45fF
C14189 a_25744_7638# a_25398_17524# 0.38fF
C14190 a_8491_27023# a_18370_17524# 0.38fF
C14191 a_11067_46823# a_39673_28111# 0.60fF
C14192 a_26402_9492# a_27406_9492# 0.97fF
C14193 vcm_commonmode a_23298_12870# 0.31fF
C14194 a_20359_29199# a_16510_8760# 0.50fF
C14195 a_8531_70543# a_2419_48783# 3.18fF
C14196 a_27406_13508# a_27406_12504# 1.00fF
C14197 a_42466_67214# ctopp 3.59fF
C14198 a_32121_44545# a_32695_43455# 0.58fF
C14199 a_42466_16520# a_43470_16520# 0.97fF
C14200 a_11803_64239# VDD 0.39fF
C14201 a_48490_63198# a_48490_62194# 1.00fF
C14202 a_17696_29967# VDD 0.37fF
C14203 vcm_commonmode a_30418_58178# 0.87fF
C14204 a_77664_39480# VDD 0.46fF
C14205 vcm_commonmode a_18278_21906# 0.31fF
C14206 a_8384_40303# VDD 0.74fF
C14207 a_27869_50095# a_20359_29199# 1.27fF
C14208 a_16746_17522# VDD 33.20fF
C14209 a_9577_60437# VDD 0.40fF
C14210 a_39223_32463# a_12877_16911# 0.41fF
C14211 a_25953_32143# VDD 0.57fF
C14212 vcm_commonmode a_23298_17890# 0.31fF
C14213 a_12357_37999# a_13349_37973# 0.73fF
C14214 a_48490_67214# a_49494_67214# 0.97fF
C14215 a_17366_67214# a_17366_66210# 1.00fF
C14216 a_43267_31055# ctopp 2.63fF
C14217 a_4443_46607# a_5831_39189# 1.19fF
C14218 a_4839_43780# VDD 0.52fF
C14219 vcm_commonmode a_47486_67214# 0.87fF
C14220 a_43470_63198# VDD 0.57fF
C14221 a_30326_13874# a_30418_13508# 0.32fF
C14222 a_22448_37253# VDD 1.81fF
C14223 a_1761_44111# a_1803_20719# 4.71fF
C14224 a_35346_68218# a_35438_68218# 0.32fF
C14225 a_40050_48463# a_45478_58178# 0.38fF
C14226 a_14287_51175# a_12257_56623# 0.40fF
C14227 a_20359_29199# a_18703_29199# 1.25fF
C14228 vcm_commonmode a_17366_69222# 1.83fF
C14229 a_37446_59182# VDD 0.51fF
C14230 a_34434_7484# a_35438_7484# 0.97fF
C14231 vcm_commonmode a_44474_9492# 0.87fF
C14232 m3_49396_59094# VDD 0.34fF
C14233 a_5915_30511# VDD 0.34fF
C14234 a_11067_67279# a_16746_20534# 2.28fF
C14235 a_41462_64202# ctopp 3.59fF
C14236 ctopn a_46482_13508# 3.59fF
C14237 a_16955_52047# a_19807_28111# 0.31fF
C14238 a_2315_24540# a_3143_22364# 1.22fF
C14239 vcm_commonmode a_44382_59182# 0.31fF
C14240 a_1768_16367# a_1768_13103# 0.85fF
C14241 vcm_commonmode a_24394_22544# 0.87fF
C14242 a_3339_30503# a_20505_29967# 0.48fF
C14243 a_42099_43177# VDD 0.69fF
C14244 a_18370_69222# a_19374_69222# 0.97fF
C14245 a_17366_18528# VDD 0.57fF
C14246 a_41967_31375# a_42466_13508# 0.38fF
C14247 a_22015_28111# a_35601_27497# 0.31fF
C14248 a_45478_9492# a_46482_9492# 0.97fF
C14249 a_28410_64202# a_29414_64202# 0.97fF
C14250 a_46482_13508# a_46482_12504# 1.00fF
C14251 vcm_commonmode a_24302_18894# 0.31fF
C14252 a_17366_66210# ctopp 3.43fF
C14253 a_2830_15431# a_2926_15253# 0.44fF
C14254 a_35079_46831# VDD 0.38fF
C14255 a_36613_48169# a_37446_69222# 0.38fF
C14256 a_49494_21540# VDD 1.21fF
C14257 a_25398_22544# a_26402_22544# 0.97fF
C14258 a_27752_7638# VDD 7.35fF
C14259 vcm_commonmode a_20378_14512# 0.87fF
C14260 a_8958_65961# VDD 1.06fF
C14261 a_26402_10496# VDD 0.51fF
C14262 a_32887_40767# VDD 0.97fF
C14263 a_1586_66567# a_1923_59583# 0.49fF
C14264 vcm_commonmode a_46482_64202# 0.87fF
C14265 a_11067_13095# a_6473_40277# 0.31fF
C14266 a_41462_60186# VDD 0.51fF
C14267 a_5363_30503# a_20881_28111# 0.41fF
C14268 vcm_commonmode a_33338_10862# 0.31fF
C14269 a_36507_31573# VDD 0.74fF
C14270 a_1768_16367# a_2007_21237# 0.61fF
C14271 a_48490_65206# ctopp 3.43fF
C14272 a_4351_67279# a_11303_53511# 0.63fF
C14273 a_2317_28892# a_2315_24540# 0.33fF
C14274 a_32121_42369# a_32887_42405# 0.34fF
C14275 a_1586_36727# config_2_in[2] 0.36fF
C14276 a_1586_66567# a_9485_62613# 0.50fF
C14277 a_36442_67214# a_36442_66210# 1.00fF
C14278 vcm_commonmode a_48398_60186# 0.31fF
C14279 vcm_commonmode a_25398_23548# 0.87fF
C14280 a_27359_43985# VDD 0.96fF
C14281 a_29760_55394# a_12983_63151# 0.40fF
C14282 vcm_commonmode a_22386_66210# 0.87fF
C14283 a_24029_39355# a_1761_27791# 1.09fF
C14284 a_32426_65206# a_32426_64202# 1.00fF
C14285 a_49402_13874# a_49494_13508# 0.32fF
C14286 vcm_commonmode a_34434_19532# 0.87fF
C14287 ctopn a_16746_16518# 1.68fF
C14288 a_31768_55394# a_12981_62313# 0.40fF
C14289 vcm_commonmode a_20286_62194# 0.31fF
C14290 a_19807_28111# a_15607_46805# 0.78fF
C14291 a_21382_15516# VDD 0.51fF
C14292 a_11035_47893# VDD 0.40fF
C14293 a_10055_58791# a_2419_48783# 0.63fF
C14294 a_26402_23548# a_26402_22544# 1.00fF
C14295 vcm_commonmode a_28318_15882# 0.31fF
C14296 a_21382_63198# ctopp 3.64fF
C14297 a_39299_48783# a_16863_29415# 0.54fF
C14298 a_35346_56170# a_35438_56170# 0.32fF
C14299 a_19374_71230# VDD 0.58fF
C14300 a_20378_66210# a_20378_65206# 1.00fF
C14301 a_17599_52263# a_22386_59182# 0.38fF
C14302 a_21382_14512# a_22386_14512# 0.97fF
C14303 a_7910_38671# VDD 0.52fF
C14304 a_31422_11500# VDD 0.51fF
C14305 a_18045_41281# VDD 1.38fF
C14306 a_37446_69222# a_38450_69222# 0.97fF
C14307 a_12889_35537# a_12663_35431# 0.39fF
C14308 a_12792_51017# VDD 0.33fF
C14309 vcm_commonmode a_26310_71230# 0.31fF
C14310 a_32426_61190# a_32426_60186# 1.00fF
C14311 a_18278_8854# a_18370_8488# 0.32fF
C14312 a_35438_24552# VDD 0.60fF
C14313 vcm_commonmode a_38358_11866# 0.31fF
C14314 a_2840_66103# a_34411_50613# 0.35fF
C14315 a_2191_68565# a_4500_45289# 0.32fF
C14316 a_29760_7638# a_12546_22351# 0.41fF
C14317 a_4563_32900# a_4495_35925# 0.71fF
C14318 a_47486_64202# a_48490_64202# 0.97fF
C14319 a_7695_31573# VDD 3.53fF
C14320 a_41427_52263# a_25419_50959# 7.84fF
C14321 a_12899_3311# a_12899_2767# 18.97fF
C14322 a_1770_14441# a_1768_16367# 2.16fF
C14323 a_12877_16911# a_16362_13508# 1.27fF
C14324 vcm_commonmode a_42374_24918# 0.31fF
C14325 a_7862_34025# a_19626_31751# 1.21fF
C14326 a_7939_30503# a_12935_31287# 0.93fF
C14327 a_4443_46607# a_7571_29199# 0.74fF
C14328 a_19282_70226# a_19374_70226# 0.32fF
C14329 a_25787_28327# a_12727_67753# 0.40fF
C14330 a_45478_55166# VDD 0.60fF
C14331 a_44474_22544# a_45478_22544# 0.97fF
C14332 a_18370_62194# a_18370_61190# 1.00fF
C14333 a_9361_28335# VDD 0.58fF
C14334 a_37446_57174# VDD 0.51fF
C14335 a_23736_7638# a_12985_7663# 0.41fF
C14336 a_49402_70226# VDD 0.31fF
C14337 a_35438_65206# a_36442_65206# 0.97fF
C14338 a_27981_37477# VDD 1.43fF
C14339 vcm_commonmode a_37446_20536# 0.87fF
C14340 a_13837_39860# VDD 2.24fF
C14341 a_18611_52047# a_23390_64202# 0.38fF
C14342 vcm_commonmode a_26402_63198# 0.92fF
C14343 a_31422_17524# a_31422_16520# 1.00fF
C14344 vcm_commonmode a_44382_57174# 0.31fF
C14345 a_23019_48463# VDD 0.38fF
C14346 a_14287_51175# a_8531_70543# 0.31fF
C14347 a_18370_20536# a_18370_19532# 1.00fF
C14348 a_1768_13103# config_2_in[2] 1.89fF
C14349 a_11067_63143# a_12985_19087# 0.44fF
C14350 a_26402_23548# a_27406_23548# 0.97fF
C14351 a_45478_58178# ctopp 3.59fF
C14352 a_23395_52047# VDD 12.87fF
C14353 vcm_commonmode a_20378_59182# 0.87fF
C14354 a_23390_66210# a_24394_66210# 0.97fF
C14355 VDD dummypin[3] 0.86fF
C14356 a_6559_22671# a_2787_32679# 0.47fF
C14357 a_14287_51175# a_10975_66407# 0.42fF
C14358 a_41427_52263# a_23395_32463# 0.54fF
C14359 a_12473_37429# a_12663_35431# 0.47fF
C14360 vcm_commonmode a_28547_51175# 10.08fF
C14361 a_36629_27791# a_12985_16367# 0.41fF
C14362 a_34342_61190# a_34434_61190# 0.32fF
C14363 a_8491_27023# VDD 13.37fF
C14364 a_8583_33551# VDD 15.84fF
C14365 vcm_commonmode a_37446_12504# 0.87fF
C14366 a_19374_60186# ctopp 3.59fF
C14367 ctopn a_38450_9492# 3.58fF
C14368 a_22386_68218# VDD 0.51fF
C14369 a_28195_35327# VDD 1.03fF
C14370 a_22294_7850# VDD 0.62fF
C14371 ctopn a_18370_22544# 3.57fF
C14372 VDD dummypin[1] 1.00fF
C14373 a_7387_46831# a_6559_22671# 0.35fF
C14374 a_18539_47617# VDD 0.36fF
C14375 a_23390_71230# a_23390_70226# 1.00fF
C14376 vcm_commonmode a_29322_68218# 0.31fF
C14377 a_34251_52263# a_12901_66959# 0.40fF
C14378 a_35438_19532# a_36442_19532# 0.97fF
C14379 a_3247_20495# a_5309_25853# 0.43fF
C14380 a_45478_23548# a_45478_22544# 1.00fF
C14381 a_2467_29397# VDD 0.37fF
C14382 a_12349_25847# a_10964_25615# 1.32fF
C14383 a_3143_22364# a_3355_25071# 0.31fF
C14384 a_39454_66210# a_39454_65206# 1.00fF
C14385 a_40458_14512# a_41462_14512# 0.97fF
C14386 vcm_commonmode a_32426_21540# 0.87fF
C14387 a_46482_72234# m3_46384_72146# 2.80fF
C14388 a_33543_41271# VDD 0.67fF
C14389 a_21371_52263# a_26402_65206# 0.38fF
C14390 a_41462_72234# a_42466_72234# 0.97fF
C14391 a_19374_20536# a_20378_20536# 0.97fF
C14392 a_1757_23445# VDD 0.58fF
C14393 a_37354_8854# a_37446_8488# 0.32fF
C14394 a_4339_64521# a_4758_45369# 0.39fF
C14395 vcm_commonmode a_37446_17524# 0.87fF
C14396 a_7499_74031# VDD 0.40fF
C14397 vcm_commonmode a_24394_60186# 0.87fF
C14398 a_2787_30503# a_15548_30761# 0.71fF
C14399 a_36442_13508# VDD 0.51fF
C14400 a_34222_43439# VDD 0.53fF
C14401 a_38358_70226# a_38450_70226# 0.32fF
C14402 a_41261_28335# a_42466_68218# 0.38fF
C14403 a_41967_31375# a_42466_7484# 0.34fF
C14404 a_19807_28111# a_15681_27497# 0.68fF
C14405 a_1761_40847# a_12381_35836# 0.31fF
C14406 a_1586_51335# a_8500_58799# 0.89fF
C14407 a_37446_62194# a_37446_61190# 1.00fF
C14408 a_10515_63143# a_5190_59575# 0.94fF
C14409 a_12707_26159# VDD 1.07fF
C14410 a_28410_10496# a_28410_9492# 1.00fF
C14411 a_22386_56170# VDD 0.52fF
C14412 vcm_commonmode a_43378_13874# 0.31fF
C14413 a_19282_16886# a_19374_16520# 0.32fF
C14414 vcm_commonmode a_29322_56170# 0.31fF
C14415 a_17599_52263# a_22386_57174# 0.38fF
C14416 ctopn a_19374_23548# 3.39fF
C14417 a_11067_46823# a_12907_27023# 0.43fF
C14418 a_23395_52047# a_27406_70226# 0.38fF
C14419 a_37446_20536# a_37446_19532# 1.00fF
C14420 a_6559_22671# a_5531_22895# 0.31fF
C14421 a_45478_23548# a_46482_23548# 0.97fF
C14422 a_39222_48169# a_40458_60186# 0.38fF
C14423 a_42466_66210# a_43470_66210# 0.97fF
C14424 a_18151_52263# a_11251_59879# 6.21fF
C14425 ctopn a_28410_19532# 3.59fF
C14426 a_1761_49007# a_12663_40871# 0.55fF
C14427 a_5179_10927# VDD 0.41fF
C14428 a_16707_42359# VDD 0.62fF
C14429 a_29760_55394# a_29414_66210# 0.38fF
C14430 a_39389_52271# a_12355_65103# 0.40fF
C14431 a_33864_28111# a_34434_9492# 0.38fF
C14432 a_28968_50871# VDD 0.43fF
C14433 a_17366_21540# a_17366_20536# 1.00fF
C14434 a_21382_61190# VDD 0.51fF
C14435 a_4417_22671# VDD 2.57fF
C14436 a_19720_7638# a_11067_21583# 0.41fF
C14437 a_4674_40277# a_5915_30287# 0.31fF
C14438 a_29513_34428# VDD 0.74fF
C14439 a_19374_12504# a_20378_12504# 0.97fF
C14440 vcm_commonmode a_38450_18528# 0.87fF
C14441 a_3987_19623# a_5490_41365# 0.68fF
C14442 a_12447_29199# a_5363_30503# 0.46fF
C14443 vcm_commonmode a_28318_61190# 0.31fF
C14444 a_28756_55394# a_28410_62194# 0.38fF
C14445 a_25306_67214# a_25398_67214# 0.32fF
C14446 vcm_commonmode a_18370_24552# 0.84fF
C14447 a_41261_28335# a_42466_56170# 0.38fF
C14448 a_14354_32117# a_12412_32143# 0.64fF
C14449 a_15607_46805# a_29927_29199# 0.33fF
C14450 a_42466_71230# a_42466_70226# 1.00fF
C14451 a_14471_28585# VDD 0.77fF
C14452 a_29414_62194# ctopp 3.59fF
C14453 a_4555_55233# a_4516_55107# 0.72fF
C14454 a_25398_70226# VDD 0.51fF
C14455 a_42466_58178# VDD 0.51fF
C14456 vcm_commonmode a_29414_55166# 0.84fF
C14457 a_41842_27221# a_12899_3311# 0.65fF
C14458 vcm_commonmode a_20378_57174# 0.87fF
C14459 a_24556_49551# VDD 0.47fF
C14460 vcm_commonmode a_32334_70226# 0.31fF
C14461 a_38450_20536# a_39454_20536# 0.97fF
C14462 vcm_commonmode a_47486_10496# 0.87fF
C14463 a_26748_7638# a_26402_20536# 0.38fF
C14464 a_39673_28111# a_40458_21540# 0.38fF
C14465 a_27406_63198# a_28410_63198# 0.97fF
C14466 a_1591_63151# VDD 2.31fF
C14467 a_35438_71230# ctopp 3.40fF
C14468 ctopn a_31422_20536# 3.59fF
C14469 a_27314_58178# a_27406_58178# 0.32fF
C14470 a_18835_52465# VDD 0.34fF
C14471 a_42718_27497# a_12877_16911# 0.41fF
C14472 a_15607_46805# a_28817_29111# 0.33fF
C14473 a_22294_9858# a_22386_9492# 0.32fF
C14474 a_47486_10496# a_47486_9492# 1.00fF
C14475 a_31422_55166# m3_31324_55078# 2.81fF
C14476 a_8782_65015# VDD 1.43fF
C14477 a_3143_22364# config_1_in[15] 0.33fF
C14478 a_43470_8488# VDD 0.58fF
C14479 vcm_commonmode a_34434_62194# 0.87fF
C14480 a_38358_16886# a_38450_16520# 0.32fF
C14481 a_26748_7638# a_26402_12504# 0.38fF
C14482 a_21382_59182# a_22386_59182# 0.97fF
C14483 a_1643_64213# VDD 0.38fF
C14484 a_8491_41383# a_8461_32937# 0.34fF
C14485 a_20103_30287# VDD 0.42fF
C14486 vcm_commonmode a_42466_15516# 0.87fF
C14487 ctopn a_31422_12504# 3.59fF
C14488 vcm_commonmode a_21290_58178# 0.31fF
C14489 a_38345_42044# VDD 1.00fF
C14490 a_4351_67279# a_4983_66959# 0.39fF
C14491 a_19374_17524# a_20378_17524# 0.97fF
C14492 vcm_commonmode a_40458_71230# 0.86fF
C14493 a_36442_21540# a_36442_20536# 1.00fF
C14494 a_9135_27239# a_12727_15529# 0.41fF
C14495 a_6607_42167# a_5449_25071# 0.37fF
C14496 a_3339_43023# a_18703_29199# 1.91fF
C14497 a_23390_24552# a_23390_23548# 1.00fF
C14498 a_40491_27247# a_11067_21583# 0.41fF
C14499 a_31422_67214# VDD 0.51fF
C14500 a_38450_12504# a_39454_12504# 0.97fF
C14501 a_12257_56623# a_12947_56817# 23.39fF
C14502 a_44382_67214# a_44474_67214# 0.32fF
C14503 a_9513_65301# a_9624_65301# 0.42fF
C14504 a_39389_52271# ctopp 2.62fF
C14505 ctopn a_26402_21540# 3.59fF
C14506 a_3339_30503# a_14926_31849# 0.85fF
C14507 a_1823_72381# a_1823_66941# 0.47fF
C14508 vcm_commonmode a_38358_67214# 0.31fF
C14509 a_3325_49551# a_4127_50069# 0.66fF
C14510 a_1643_54421# VDD 0.37fF
C14511 a_2411_19605# a_2143_15271# 0.34fF
C14512 a_26748_7638# a_26402_17524# 0.38fF
C14513 a_22015_28111# a_12899_3855# 1.05fF
C14514 vcm_commonmode a_19374_13508# 0.87fF
C14515 a_2847_69439# VDD 0.42fF
C14516 a_38450_68218# ctopp 3.59fF
C14517 ctopn a_31422_17524# 3.59fF
C14518 a_28410_9492# VDD 0.51fF
C14519 a_39836_38567# VDD 1.81fF
C14520 a_3247_20495# a_6738_19783# 0.54fF
C14521 a_44474_16520# VDD 0.51fF
C14522 a_12907_56399# a_11803_55311# 7.29fF
C14523 a_30326_7850# a_30418_7484# 0.32fF
C14524 vcm_commonmode a_35346_9858# 0.31fF
C14525 a_46482_63198# a_47486_63198# 0.97fF
C14526 a_38210_30199# VDD 1.48fF
C14527 a_1761_52815# a_30757_37455# 0.60fF
C14528 a_20378_18528# a_20378_17524# 1.00fF
C14529 a_11067_47695# a_21095_47919# 0.62fF
C14530 a_2847_51157# VDD 0.36fF
C14531 a_33430_21540# a_34434_21540# 0.97fF
C14532 a_41370_9858# a_41462_9492# 0.32fF
C14533 a_43270_27791# a_45478_23548# 0.38fF
C14534 a_24302_64202# a_24394_64202# 0.32fF
C14535 a_14951_34743# VDD 0.60fF
C14536 a_36442_7484# VDD 1.25fF
C14537 a_43362_28879# a_47486_63198# 0.42fF
C14538 a_12907_56399# a_12981_62313# 0.34fF
C14539 a_4995_13103# VDD 0.41fF
C14540 ctopn m3_18272_24702# 0.35fF
C14541 a_25787_28327# a_33430_69222# 0.38fF
C14542 vcm_commonmode a_43470_68218# 0.87fF
C14543 a_40458_59182# a_41462_59182# 0.97fF
C14544 a_21290_22910# a_21382_22544# 0.32fF
C14545 a_30764_7638# a_30418_19532# 0.38fF
C14546 a_30418_64202# VDD 0.51fF
C14547 a_12447_29199# a_23395_32463# 0.31fF
C14548 a_38450_56170# ctopp 3.40fF
C14549 a_12516_7093# VDD 20.34fF
C14550 a_13183_52047# a_17366_58178# 0.38fF
C14551 a_21382_14512# a_21382_13508# 1.00fF
C14552 ctopn a_32426_18528# 3.59fF
C14553 a_2539_42106# a_1761_25071# 0.99fF
C14554 vcm_commonmode a_37354_64202# 0.31fF
C14555 a_38450_17524# a_39454_17524# 0.97fF
C14556 a_21187_29415# a_20359_29199# 0.97fF
C14557 a_2606_41079# VDD 16.25fF
C14558 a_47394_72234# a_47486_72234# 0.32fF
C14559 a_42709_29199# a_48490_14512# 0.38fF
C14560 a_25398_60186# a_26402_60186# 0.97fF
C14561 a_42466_24552# a_42466_23548# 1.00fF
C14562 a_39673_28111# a_12985_7663# 0.41fF
C14563 a_8491_41383# a_7598_36103# 0.38fF
C14564 a_16746_63200# a_12981_62313# 0.41fF
C14565 a_8117_30287# VDD 1.03fF
C14566 a_27406_12504# a_27406_11500# 1.00fF
C14567 a_41872_29423# a_12981_59343# 0.40fF
C14568 a_28757_27247# a_30440_31573# 0.32fF
C14569 a_17599_52263# a_12983_63151# 0.40fF
C14570 a_20378_18528# a_21382_18528# 0.97fF
C14571 a_18370_19532# VDD 0.52fF
C14572 a_13445_50639# a_12993_50345# 0.62fF
C14573 a_10975_60975# a_11141_60975# 0.66fF
C14574 a_10055_58791# a_40675_27791# 0.41fF
C14575 a_37446_61190# ctopp 3.59fF
C14576 ctopn a_41462_10496# 3.59fF
C14577 a_39223_32463# a_12895_13967# 0.41fF
C14578 a_39454_69222# VDD 0.51fF
C14579 vcm_commonmode a_25306_19898# 0.31fF
C14580 a_18151_52263# a_12981_62313# 0.40fF
C14581 vcm_commonmode a_43470_56170# 0.87fF
C14582 a_1761_34319# a_36890_34191# 0.44fF
C14583 a_2467_47893# VDD 0.50fF
C14584 vcm_commonmode a_46390_69222# 0.31fF
C14585 a_49402_7850# a_49494_7484# 0.32fF
C14586 a_46482_22544# VDD 0.51fF
C14587 vcm_commonmode a_26402_8488# 0.86fF
C14588 a_37446_65206# VDD 0.51fF
C14589 a_30891_28309# VDD 0.49fF
C14590 a_17222_27247# a_17712_7638# 0.31fF
C14591 a_14287_51175# a_18370_59182# 0.38fF
C14592 a_17274_14878# a_17366_14512# 0.32fF
C14593 a_41462_70226# ctopp 3.58fF
C14594 a_32970_31145# a_34759_31029# 3.39fF
C14595 a_33338_69222# a_33430_69222# 0.32fF
C14596 vcm_commonmode a_44382_65206# 0.31fF
C14597 a_39454_18528# a_39454_17524# 1.00fF
C14598 a_12641_36596# a_1761_31055# 2.59fF
C14599 a_18151_52263# a_24394_72234# 0.35fF
C14600 vcm_commonmode a_16362_71230# 4.46fF
C14601 a_10515_63143# a_3339_32463# 2.01fF
C14602 a_43269_29967# a_47486_14512# 0.38fF
C14603 a_26310_24918# VDD 0.36fF
C14604 a_43378_64202# a_43470_64202# 0.32fF
C14605 a_5595_33205# VDD 0.90fF
C14606 ctopn a_36442_15516# 3.59fF
C14607 a_1586_21959# a_3325_18543# 1.41fF
C14608 vcm_commonmode a_42466_61190# 0.87fF
C14609 a_8123_14741# a_8289_14741# 0.57fF
C14610 a_42466_14512# VDD 0.51fF
C14611 a_8263_45908# VDD 0.31fF
C14612 a_21371_52263# a_12727_67753# 0.40fF
C14613 a_13123_38231# a_12473_37429# 1.25fF
C14614 a_21382_20536# VDD 0.51fF
C14615 a_36350_55166# VDD 0.35fF
C14616 a_40366_22910# a_40458_22544# 0.32fF
C14617 a_11067_63143# VDD 5.57fF
C14618 a_29414_10496# a_30418_10496# 0.97fF
C14619 vcm_commonmode a_49402_14878# 0.30fF
C14620 ctopn a_46482_11500# 3.59fF
C14621 a_15397_39631# a_13576_40413# 0.32fF
C14622 a_31330_65206# a_31422_65206# 0.32fF
C14623 a_40458_14512# a_40458_13508# 1.00fF
C14624 vcm_commonmode a_28318_20902# 0.31fF
C14625 a_12889_39889# VDD 2.12fF
C14626 a_19720_55394# a_19374_64202# 0.38fF
C14627 vcm_commonmode a_17274_63198# 0.33fF
C14628 vcm_commonmode a_46482_70226# 0.87fF
C14629 a_41967_31375# a_42466_11500# 0.38fF
C14630 a_44474_60186# a_45478_60186# 0.97fF
C14631 a_53260_40156# a_7841_12167# 1.08fF
C14632 a_47486_23548# VDD 0.52fF
C14633 a_30418_58178# ctopp 3.59fF
C14634 a_25744_7638# a_25398_21540# 0.38fF
C14635 a_22294_23914# a_22386_23548# 0.32fF
C14636 a_8491_27023# a_18370_21540# 0.38fF
C14637 a_44474_66210# VDD 0.51fF
C14638 VDD dummypin[15] 0.65fF
C14639 a_46482_12504# a_46482_11500# 1.00fF
C14640 vcm_commonmode a_27406_16520# 0.87fF
C14641 a_16955_52047# VDD 15.48fF
C14642 a_19282_66210# a_19374_66210# 0.32fF
C14643 a_44474_7484# m3_44376_7346# 2.80fF
C14644 a_3607_34639# a_7841_29673# 0.34fF
C14645 a_21382_12504# VDD 0.51fF
C14646 a_33430_70226# a_33430_69222# 1.00fF
C14647 a_12516_7093# a_11619_56615# 2.16fF
C14648 a_3143_66972# a_3024_67191# 0.65fF
C14649 a_39454_18528# a_40458_18528# 0.97fF
C14650 a_2872_44111# a_2292_43291# 0.80fF
C14651 a_8051_52047# VDD 0.43fF
C14652 vcm_commonmode a_21371_50959# 10.02fF
C14653 a_41462_55166# m3_41364_55078# 2.81fF
C14654 vcm_commonmode a_28318_12870# 0.31fF
C14655 a_19374_24552# a_20378_24552# 0.97fF
C14656 a_5211_24759# a_7059_24135# 0.58fF
C14657 a_47486_67214# ctopp 3.58fF
C14658 a_12549_44212# a_22671_43439# 0.30fF
C14659 a_3024_67191# a_1823_65853# 0.72fF
C14660 a_27535_30503# a_18979_30287# 0.87fF
C14661 a_20359_29199# a_26523_28111# 1.16fF
C14662 a_28756_55394# a_12901_66959# 0.40fF
C14663 a_31330_19898# a_31422_19532# 0.32fF
C14664 a_16746_21538# VDD 33.21fF
C14665 vcm_commonmode a_19374_7484# 0.69fF
C14666 a_9135_27239# a_21382_19532# 0.38fF
C14667 a_4647_63937# VDD 0.49fF
C14668 a_19807_28111# a_30565_30199# 0.64fF
C14669 a_32038_29575# VDD 0.63fF
C14670 a_32426_11500# a_32426_10496# 1.00fF
C14671 a_38557_32143# a_12907_27023# 0.72fF
C14672 a_1761_41935# a_14293_39631# 1.94fF
C14673 vcm_commonmode a_35438_58178# 0.87fF
C14674 a_36350_14878# a_36442_14512# 0.32fF
C14675 vcm_commonmode a_23298_21906# 0.31fF
C14676 a_17366_69222# ctopp 3.43fF
C14677 a_33694_30761# a_41597_29967# 0.31fF
C14678 a_1761_47919# a_1803_19087# 1.30fF
C14679 a_17599_52263# a_22386_65206# 0.38fF
C14680 a_21382_17524# VDD 0.51fF
C14681 a_23631_50069# VDD 0.72fF
C14682 a_38557_32143# a_39389_52271# 0.31fF
C14683 a_32951_27247# a_12727_15529# 0.41fF
C14684 a_30418_55166# a_31422_55166# 0.97fF
C14685 a_12869_2741# a_10873_27497# 0.52fF
C14686 a_2124_63419# a_2163_63293# 0.73fF
C14687 a_30052_32117# VDD 2.66fF
C14688 vcm_commonmode a_28318_17890# 0.31fF
C14689 a_21382_57174# a_22386_57174# 0.97fF
C14690 a_24394_15516# a_25398_15516# 0.97fF
C14691 a_1586_40455# a_3247_20495# 0.36fF
C14692 a_38557_32143# a_38450_68218# 0.38fF
C14693 a_48490_63198# VDD 0.60fF
C14694 a_12447_29199# a_18162_31055# 0.55fF
C14695 a_48490_10496# a_49494_10496# 0.97fF
C14696 a_11067_13095# a_16362_64202# 19.83fF
C14697 a_31847_36893# VDD 2.01fF
C14698 a_15851_27791# a_15661_29199# 0.73fF
C14699 a_1761_44111# a_1761_43567# 1.15fF
C14700 a_5682_69367# a_6515_62037# 1.30fF
C14701 a_14287_51175# a_18370_57174# 0.38fF
C14702 a_15607_46805# VDD 15.02fF
C14703 vcm_commonmode a_22386_69222# 0.87fF
C14704 a_18611_52047# a_23390_70226# 0.38fF
C14705 a_22386_71230# a_23390_71230# 0.97fF
C14706 a_42466_59182# VDD 0.51fF
C14707 vcm_commonmode a_49494_9492# 0.89fF
C14708 a_41370_23914# a_41462_23548# 0.32fF
C14709 a_12869_2741# a_19889_27497# 0.59fF
C14710 a_20946_30669# VDD 1.21fF
C14711 a_34434_11500# a_35438_11500# 0.97fF
C14712 a_9642_10357# a_10259_10703# 0.40fF
C14713 a_46482_64202# ctopp 3.59fF
C14714 a_48490_72234# VDD 1.28fF
C14715 a_11619_56615# a_11067_63143# 6.13fF
C14716 vcm_commonmode a_49402_59182# 0.30fF
C14717 a_36717_47375# a_36442_60186# 0.38fF
C14718 a_38358_66210# a_38450_66210# 0.32fF
C14719 a_11067_67279# a_10515_63143# 0.45fF
C14720 vcm_commonmode a_29414_22544# 0.87fF
C14721 a_28547_51175# a_12355_65103# 0.40fF
C14722 vcm_commonmode a_20378_65206# 0.87fF
C14723 a_21371_50959# a_25398_66210# 0.38fF
C14724 a_22386_18528# VDD 0.51fF
C14725 a_37919_28111# a_38450_16520# 0.38fF
C14726 a_29760_7638# a_12985_16367# 0.41fF
C14727 a_43175_28335# a_12727_15529# 0.41fF
C14728 ctopn a_20378_8488# 3.40fF
C14729 a_19720_7638# a_12546_22351# 0.41fF
C14730 a_38450_24552# a_39454_24552# 0.97fF
C14731 a_12869_2741# a_12263_4391# 2.17fF
C14732 vcm_commonmode a_29322_18894# 0.31fF
C14733 a_22386_66210# ctopp 3.59fF
C14734 a_18151_52263# a_24394_62194# 0.38fF
C14735 a_38557_32143# a_38450_56170# 0.38fF
C14736 a_2840_53511# a_6559_59663# 0.71fF
C14737 a_35438_62194# a_36442_62194# 0.97fF
C14738 a_5291_56765# VDD 0.41fF
C14739 vcm_commonmode a_25398_14512# 0.87fF
C14740 a_24768_27247# a_24683_27497# 0.36fF
C14741 a_1586_21959# a_6816_19355# 0.98fF
C14742 a_12135_69109# VDD 0.51fF
C14743 a_22411_38007# VDD 0.59fF
C14744 a_11067_67279# a_35601_27497# 0.41fF
C14745 vcm_commonmode a_20286_55166# 0.30fF
C14746 a_2787_32679# a_2021_22325# 0.43fF
C14747 a_31422_10496# VDD 0.51fF
C14748 a_77086_40693# VDD 119.67fF
C14749 a_8531_70543# a_2840_66103# 1.04fF
C14750 a_34342_20902# a_34434_20536# 0.32fF
C14751 a_46482_60186# VDD 0.51fF
C14752 vcm_commonmode a_38358_10862# 0.31fF
C14753 a_23298_63198# a_23390_63198# 0.32fF
C14754 a_11067_67279# a_12985_7663# 25.91fF
C14755 a_11902_27497# a_17278_28309# 0.40fF
C14756 a_1803_19087# a_23789_39100# 0.49fF
C14757 a_40458_57174# a_41462_57174# 0.97fF
C14758 a_43470_15516# a_44474_15516# 0.97fF
C14759 vcm_commonmode a_30418_23548# 0.87fF
C14760 vcm_commonmode a_27406_66210# 0.87fF
C14761 a_18370_62194# VDD 0.52fF
C14762 a_3987_19623# a_5449_25071# 1.79fF
C14763 a_15607_46805# a_18053_28879# 0.68fF
C14764 a_24394_55166# m3_24296_55078# 2.81fF
C14765 a_7841_12167# a_1929_12131# 0.51fF
C14766 a_10055_58791# a_16510_8760# 1.07fF
C14767 vcm_commonmode a_39454_19532# 0.87fF
C14768 ctopn a_21382_16520# 3.59fF
C14769 a_12381_43957# a_12357_37999# 0.36fF
C14770 vcm_commonmode a_25306_62194# 0.31fF
C14771 a_26402_15516# VDD 0.51fF
C14772 a_41462_71230# a_42466_71230# 0.97fF
C14773 a_17274_59182# a_17366_59182# 0.32fF
C14774 a_1681_5175# a_1761_6031# 0.45fF
C14775 m3_34336_7346# VDD 0.33fF
C14776 a_3339_32463# a_9135_29423# 0.31fF
C14777 a_19807_28111# a_26523_29199# 0.36fF
C14778 a_7479_54439# a_17039_51157# 0.35fF
C14779 a_9963_29967# VDD 0.39fF
C14780 vcm_commonmode a_33338_15882# 0.31fF
C14781 a_26402_63198# ctopp 3.64fF
C14782 a_24394_71230# VDD 0.58fF
C14783 a_21479_39141# VDD 0.84fF
C14784 a_36442_11500# VDD 0.51fF
C14785 a_43175_28335# a_46482_8488# 0.38fF
C14786 a_3987_19623# a_5239_20693# 0.31fF
C14787 a_5691_36727# a_3339_30503# 0.48fF
C14788 vcm_commonmode a_31330_71230# 0.31fF
C14789 a_43270_27791# a_12727_15529# 0.41fF
C14790 a_40491_27247# a_43470_16520# 0.38fF
C14791 a_3016_60949# a_4674_57685# 0.53fF
C14792 a_40458_24552# VDD 0.60fF
C14793 vcm_commonmode a_43378_11866# 0.31fF
C14794 a_20378_59182# ctopp 3.59fF
C14795 a_40491_27247# a_12546_22351# 0.41fF
C14796 a_6835_46823# a_12869_2741# 0.44fF
C14797 a_21382_64202# a_21382_63198# 1.23fF
C14798 a_34342_12870# a_34434_12504# 0.32fF
C14799 a_7565_31751# VDD 0.46fF
C14800 vcm_commonmode a_47394_24918# 0.30fF
C14801 a_28547_51175# ctopp 2.66fF
C14802 a_29414_59182# a_29414_58178# 1.00fF
C14803 a_1761_52815# a_1761_50639# 2.34fF
C14804 a_6831_63303# a_9301_49557# 0.62fF
C14805 a_15681_27497# VDD 2.32fF
C14806 a_42466_57174# VDD 0.51fF
C14807 a_6095_44807# a_7891_64213# 0.38fF
C14808 a_40343_37737# VDD 0.60fF
C14809 a_20378_13508# a_21382_13508# 0.97fF
C14810 vcm_commonmode a_42466_20536# 0.87fF
C14811 a_38210_30199# a_38436_29941# 0.83fF
C14812 a_12725_44527# a_17863_44211# 0.97fF
C14813 a_21387_39679# VDD 0.87fF
C14814 vcm_commonmode a_31422_63198# 0.92fF
C14815 a_25398_68218# a_26402_68218# 0.97fF
C14816 vcm_commonmode a_49402_57174# 0.30fF
C14817 a_37446_56170# a_37446_55166# 1.00fF
C14818 a_42374_63198# a_42466_63198# 0.32fF
C14819 a_42466_58178# a_43470_58178# 0.97fF
C14820 a_23928_28585# a_17712_7638# 2.50fF
C14821 a_33430_57174# a_33430_56170# 1.00fF
C14822 vcm_commonmode a_25398_59182# 0.87fF
C14823 a_1761_50639# a_12641_42036# 0.34fF
C14824 a_30663_51727# VDD 0.60fF
C14825 a_29322_21906# a_29414_21540# 0.32fF
C14826 a_7571_29199# a_12899_3311# 2.36fF
C14827 a_2847_26133# VDD 0.46fF
C14828 vcm_commonmode a_42466_12504# 0.87fF
C14829 a_24394_60186# ctopp 3.59fF
C14830 ctopn a_43470_9492# 3.58fF
C14831 a_32772_7638# a_11067_21583# 0.41fF
C14832 a_27406_68218# VDD 0.51fF
C14833 a_11711_12559# a_11416_12283# 0.57fF
C14834 a_27314_7850# VDD 0.61fF
C14835 a_47394_58178# a_47486_58178# 0.32fF
C14836 a_41872_29423# a_43470_63198# 0.42fF
C14837 a_5024_67885# a_7213_62215# 1.14fF
C14838 a_17366_16520# a_17366_15516# 1.00fF
C14839 ctopn a_23390_22544# 3.58fF
C14840 a_34482_29941# a_15607_46805# 1.64fF
C14841 vcm_commonmode a_34342_68218# 0.31fF
C14842 a_29760_55394# a_29414_69222# 0.38fF
C14843 a_36350_59182# a_36442_59182# 0.32fF
C14844 a_10687_52553# a_29361_51727# 0.73fF
C14845 a_16746_22542# a_11067_21583# 2.28fF
C14846 a_28756_7638# a_12899_10927# 0.41fF
C14847 a_42718_27497# a_12895_13967# 0.41fF
C14848 a_26523_28111# a_28446_31375# 0.44fF
C14849 a_8531_70543# a_14831_50095# 1.06fF
C14850 a_12349_25847# a_9135_27239# 0.31fF
C14851 a_2656_70197# VDD 0.31fF
C14852 vcm_commonmode a_37446_21540# 0.87fF
C14853 a_1761_50639# a_14963_39783# 0.75fF
C14854 a_1591_9839# VDD 0.43fF
C14855 a_2847_40277# VDD 0.51fF
C14856 a_34342_17890# a_34434_17524# 0.32fF
C14857 a_35224_49871# VDD 0.55fF
C14858 a_21290_60186# a_21382_60186# 0.32fF
C14859 a_11067_67279# a_7571_26151# 2.64fF
C14860 a_40458_64202# a_40458_63198# 1.23fF
C14861 config_2_in[2] start_conversion_in 0.41fF
C14862 vcm_commonmode a_42466_17524# 0.87fF
C14863 ctopn a_19374_14512# 3.59fF
C14864 vcm_commonmode a_29414_60186# 0.87fF
C14865 a_36717_47375# a_12981_59343# 0.40fF
C14866 a_13357_32143# a_25313_31599# 0.42fF
C14867 a_14646_29423# a_20881_28111# 0.35fF
C14868 a_3339_30503# a_17358_31069# 0.44fF
C14869 a_41462_13508# VDD 0.51fF
C14870 a_13716_43047# VDD 6.41fF
C14871 a_16362_18528# a_16746_18526# 2.28fF
C14872 a_1586_9991# VDD 5.55fF
C14873 a_2952_53333# VDD 1.50fF
C14874 a_42718_27497# a_44474_18528# 0.38fF
C14875 a_32426_22544# a_32426_21540# 1.00fF
C14876 a_5535_18012# a_7377_18012# 1.68fF
C14877 a_1761_40847# a_1761_35407# 1.52fF
C14878 a_8583_33551# a_26397_51183# 0.85fF
C14879 a_27406_56170# VDD 0.52fF
C14880 vcm_commonmode a_48398_13874# 0.31fF
C14881 a_39454_13508# a_40458_13508# 0.97fF
C14882 a_28756_55394# a_28410_55166# 0.46fF
C14883 a_44474_68218# a_45478_68218# 0.97fF
C14884 vcm_commonmode a_34342_56170# 0.31fF
C14885 ctopn a_24394_23548# 3.40fF
C14886 a_7939_30503# a_7862_34025# 1.18fF
C14887 a_26417_47919# VDD 1.71fF
C14888 vcm_commonmode a_17274_8854# 0.33fF
C14889 a_20378_57174# ctopp 3.58fF
C14890 a_25398_56170# a_26402_56170# 0.97fF
C14891 ctopn a_33430_19532# 3.59fF
C14892 vcm_commonmode m3_16264_23410# 3.05fF
C14893 a_26815_42405# VDD 1.00fF
C14894 a_28756_7638# a_28410_8488# 0.38fF
C14895 a_12641_36596# a_19096_36513# 2.46fF
C14896 a_48398_21906# a_48490_21540# 0.32fF
C14897 a_26402_61190# VDD 0.51fF
C14898 vcm_commonmode a_19374_11500# 0.87fF
C14899 a_29414_58178# a_29414_57174# 1.00fF
C14900 a_37919_28111# a_11067_21583# 0.41fF
C14901 vcm_commonmode a_43470_18528# 0.87fF
C14902 a_2127_4943# VDD 0.45fF
C14903 vcm_commonmode a_33338_61190# 0.31fF
C14904 a_36442_16520# a_36442_15516# 1.00fF
C14905 vcm_commonmode a_23390_24552# 0.84fF
C14906 a_26514_47375# a_26417_47919# 1.53fF
C14907 a_19720_55394# a_12727_67753# 0.40fF
C14908 a_21382_19532# a_21382_18528# 1.00fF
C14909 a_8295_47388# a_4191_33449# 1.29fF
C14910 a_6831_63303# a_19885_50095# 0.59fF
C14911 a_8583_33551# a_25419_50959# 1.37fF
C14912 a_25306_10862# a_25398_10496# 0.32fF
C14913 a_34434_62194# ctopp 3.59fF
C14914 a_30418_70226# VDD 0.51fF
C14915 a_32367_28309# a_28817_29111# 0.86fF
C14916 a_2235_30503# a_9135_27239# 0.44fF
C14917 vcm_commonmode a_25398_57174# 0.87fF
C14918 a_2467_48981# VDD 0.43fF
C14919 a_1823_72381# a_1586_66567# 0.52fF
C14920 vcm_commonmode a_37354_70226# 0.31fF
C14921 a_12341_3311# a_12727_15529# 0.41fF
C14922 a_11067_47695# a_2143_15271# 0.69fF
C14923 a_7210_55081# a_4482_57863# 0.42fF
C14924 a_40366_60186# a_40458_60186# 0.32fF
C14925 a_10515_63143# a_1586_18695# 0.98fF
C14926 a_10515_63143# a_9240_53877# 1.03fF
C14927 a_7571_29199# a_2235_30503# 0.67fF
C14928 vcm_commonmode a_18278_16886# 0.31fF
C14929 a_2004_42453# a_4314_40821# 0.39fF
C14930 a_10147_71855# VDD 0.33fF
C14931 a_40458_71230# ctopp 3.40fF
C14932 ctopn a_36442_20536# 3.59fF
C14933 a_37446_7484# m3_37348_7346# 2.80fF
C14934 a_4563_32900# a_4674_40277# 1.58fF
C14935 a_35346_18894# a_35438_18528# 0.32fF
C14936 vcm_commonmode a_14287_51175# 10.02fF
C14937 a_6453_71855# a_6921_72943# 0.30fF
C14938 a_24394_61190# a_25398_61190# 0.97fF
C14939 a_18007_27441# VDD 0.59fF
C14940 a_34434_55166# m3_34336_55078# 2.45fF
C14941 a_10055_58791# a_25744_7638# 0.41fF
C14942 a_3693_68047# VDD 0.86fF
C14943 a_1768_16367# a_1853_27247# 0.37fF
C14944 a_4443_46607# a_1761_39215# 4.21fF
C14945 a_48490_8488# VDD 0.61fF
C14946 a_30418_68218# a_30418_67214# 1.00fF
C14947 vcm_commonmode a_39454_62194# 0.87fF
C14948 a_17507_52047# a_12901_66959# 0.40fF
C14949 a_19374_58178# VDD 0.51fF
C14950 a_32029_38565# a_32795_38591# 0.32fF
C14951 a_13669_38517# a_13837_38772# 2.20fF
C14952 a_7891_64213# VDD 0.32fF
C14953 vcm_commonmode a_47486_15516# 0.87fF
C14954 ctopn a_36442_12504# 3.59fF
C14955 a_44474_56170# a_45478_56170# 0.97fF
C14956 vcm_commonmode a_26310_58178# 0.31fF
C14957 a_2339_38129# VDD 7.07fF
C14958 a_14287_51175# a_18370_65206# 0.38fF
C14959 a_12663_35431# a_13743_35836# 0.30fF
C14960 a_34579_50613# VDD 0.89fF
C14961 a_28547_51175# a_38557_32143# 1.72fF
C14962 vcm_commonmode a_45478_71230# 0.86fF
C14963 a_34434_72234# a_35438_72234# 0.97fF
C14964 a_23395_52047# a_41872_29423# 7.46fF
C14965 a_40675_27791# a_12877_14441# 0.41fF
C14966 a_3295_54421# VDD 6.63fF
C14967 a_27406_8488# a_28410_8488# 0.97fF
C14968 a_26310_55166# a_26402_55166# 0.32fF
C14969 a_26748_7638# a_26402_21540# 0.38fF
C14970 a_36442_67214# VDD 0.51fF
C14971 a_17274_57174# a_17366_57174# 0.32fF
C14972 a_20286_15882# a_20378_15516# 0.32fF
C14973 a_41872_29423# a_8583_33551# 0.80fF
C14974 ctopn a_31422_21540# 3.59fF
C14975 a_9779_47919# a_9945_47919# 0.62fF
C14976 a_13984_43781# VDD 1.28fF
C14977 vcm_commonmode a_43378_67214# 0.31fF
C14978 a_1950_59887# a_10379_66389# 0.33fF
C14979 a_28410_70226# a_29414_70226# 0.97fF
C14980 a_34780_56398# a_34434_68218# 0.38fF
C14981 a_40458_19532# a_40458_18528# 1.00fF
C14982 a_1586_69367# a_1591_64239# 1.03fF
C14983 a_15607_46805# a_38436_29941# 0.48fF
C14984 a_44382_10862# a_44474_10496# 0.32fF
C14985 vcm_commonmode a_24394_13508# 0.87fF
C14986 a_10286_26311# a_10472_26159# 0.73fF
C14987 a_7369_24233# a_7841_22895# 0.32fF
C14988 a_12039_69367# VDD 0.76fF
C14989 a_43470_68218# ctopp 3.59fF
C14990 ctopn a_36442_17524# 3.59fF
C14991 a_8491_41383# a_8273_42479# 0.60fF
C14992 a_33430_9492# VDD 0.51fF
C14993 a_4811_34855# a_7862_34025# 0.48fF
C14994 a_49494_16520# VDD 1.24fF
C14995 a_18278_71230# a_18370_71230# 0.32fF
C14996 a_19720_55394# a_19374_70226# 0.38fF
C14997 a_43270_27791# a_45478_14512# 0.38fF
C14998 a_26402_60186# a_26402_59182# 1.00fF
C14999 vcm_commonmode a_40366_9858# 0.31fF
C15000 a_11141_65327# VDD 0.63fF
C15001 a_2411_26133# a_2012_33927# 0.57fF
C15002 a_30326_11866# a_30418_11500# 0.32fF
C15003 a_41462_72234# VDD 1.64fF
C15004 a_39299_48783# a_12727_58255# 0.40fF
C15005 a_28547_51175# a_32426_60186# 0.38fF
C15006 a_5959_13621# a_4812_13879# 0.56fF
C15007 a_35438_15516# a_35438_14512# 1.00fF
C15008 a_12727_15529# a_16746_13506# 0.41fF
C15009 vcm_commonmode a_20286_22910# 0.31fF
C15010 a_1823_77821# VDD 1.16fF
C15011 a_35463_42943# VDD 0.83fF
C15012 a_42985_46831# a_48490_67214# 0.38fF
C15013 a_21371_50959# a_12355_65103# 0.40fF
C15014 a_17507_52047# a_21382_66210# 0.38fF
C15015 a_7479_17607# VDD 0.73fF
C15016 vcm_commonmode a_46482_72234# 0.69fF
C15017 a_43470_61190# a_44474_61190# 0.97fF
C15018 a_10570_25625# VDD 0.36fF
C15019 a_20378_9492# a_20378_8488# 1.00fF
C15020 a_9503_26151# a_20378_23548# 0.38fF
C15021 a_34342_24918# a_34434_24552# 0.33fF
C15022 a_29943_34789# VDD 0.88fF
C15023 a_21371_52263# a_10687_52553# 3.13fF
C15024 a_18829_29423# a_19459_29423# 0.34fF
C15025 a_41462_7484# VDD 1.64fF
C15026 a_49494_68218# a_49494_67214# 1.00fF
C15027 a_16955_52047# a_20378_62194# 0.38fF
C15028 a_34780_56398# a_34434_56170# 0.36fF
C15029 a_21187_29415# a_38805_47081# 0.30fF
C15030 ctopn m3_33332_24990# 0.31fF
C15031 vcm_commonmode a_48490_68218# 0.87fF
C15032 a_3247_20495# a_4417_22671# 0.37fF
C15033 a_49494_59182# m3_49396_59094# 2.78fF
C15034 a_35438_64202# VDD 0.51fF
C15035 a_3016_60949# a_2959_47113# 0.51fF
C15036 a_31330_62194# a_31422_62194# 0.32fF
C15037 a_28841_29575# VDD 1.32fF
C15038 a_43470_56170# ctopp 3.40fF
C15039 a_3325_69135# VDD 1.30fF
C15040 ctopn a_37446_18528# 3.59fF
C15041 vcm_commonmode a_42374_64202# 0.31fF
C15042 a_34434_69222# a_34434_68218# 1.00fF
C15043 a_19594_35823# a_1761_32143# 1.26fF
C15044 a_46482_8488# a_47486_8488# 0.97fF
C15045 a_24394_8488# a_24394_7484# 1.00fF
C15046 a_44382_55166# a_44474_55166# 0.32fF
C15047 a_1768_16367# a_1586_40455# 1.05fF
C15048 a_4811_65871# VDD 0.63fF
C15049 a_7479_54439# a_6236_54421# 0.31fF
C15050 a_23626_31573# VDD 0.77fF
C15051 a_2840_53511# a_6646_54135# 0.74fF
C15052 a_36350_57174# a_36442_57174# 0.32fF
C15053 a_39362_15882# a_39454_15516# 0.32fF
C15054 vcm_commonmode a_21290_23914# 0.31fF
C15055 a_16362_71230# ctopp 1.17fF
C15056 vcm_commonmode a_18278_66210# 0.31fF
C15057 a_47486_70226# a_48490_70226# 0.97fF
C15058 a_17366_58178# a_18370_58178# 0.97fF
C15059 a_23390_19532# VDD 0.51fF
C15060 a_6467_55527# VDD 13.27fF
C15061 a_42466_61190# ctopp 3.59fF
C15062 ctopn a_46482_10496# 3.59fF
C15063 a_44474_69222# VDD 0.51fF
C15064 a_36395_36649# VDD 0.66fF
C15065 vcm_commonmode a_30326_19898# 0.31fF
C15066 a_6095_44807# a_8132_53511# 1.24fF
C15067 a_34780_56398# a_8295_47388# 0.39fF
C15068 a_28410_16520# a_29414_16520# 0.97fF
C15069 vcm_commonmode a_40675_27791# 10.35fF
C15070 vcm_commonmode a_48490_56170# 0.88fF
C15071 a_3607_34639# a_4903_31849# 0.45fF
C15072 VDD config_2_in[6] 0.85fF
C15073 a_37354_71230# a_37446_71230# 0.32fF
C15074 a_41967_31375# a_42466_10496# 0.38fF
C15075 a_45478_60186# a_45478_59182# 1.00fF
C15076 vcm_commonmode a_31422_8488# 0.86fF
C15077 a_1952_60431# a_2177_53359# 0.36fF
C15078 a_23736_7638# a_12727_13353# 0.41fF
C15079 a_42466_65206# VDD 0.51fF
C15080 a_34434_63198# a_34434_62194# 1.00fF
C15081 a_30565_30199# VDD 3.47fF
C15082 a_49402_11866# a_49494_11500# 0.32fF
C15083 a_41427_52263# a_13643_28327# 0.32fF
C15084 a_7289_70767# VDD 0.74fF
C15085 a_1768_13103# config_1_in[14] 0.51fF
C15086 a_1591_38677# VDD 0.44fF
C15087 a_46482_70226# ctopp 3.58fF
C15088 vcm_commonmode a_49402_65206# 0.30fF
C15089 a_1950_59887# a_6095_44807# 0.88fF
C15090 VDD config_2_in[15] 1.52fF
C15091 a_4187_60673# a_4148_60547# 0.72fF
C15092 a_39454_9492# a_39454_8488# 1.00fF
C15093 a_31330_24918# VDD 0.36fF
C15094 a_11521_66567# VDD 2.93fF
C15095 a_38115_52263# a_34759_31029# 0.62fF
C15096 ctopn a_41462_15516# 3.59fF
C15097 a_12473_42869# a_12713_43011# 2.08fF
C15098 a_6835_46823# a_7479_54439# 0.49fF
C15099 a_34434_67214# a_35438_67214# 0.97fF
C15100 vcm_commonmode a_47486_61190# 0.87fF
C15101 a_11067_67279# a_41967_31375# 0.41fF
C15102 a_21371_50959# ctopp 2.62fF
C15103 a_47486_14512# VDD 0.51fF
C15104 a_2847_45503# VDD 0.64fF
C15105 vcm_commonmode a_19374_67214# 0.87fF
C15106 a_26402_20536# VDD 0.51fF
C15107 a_41370_55166# VDD 0.35fF
C15108 a_2775_46025# a_19478_51959# 0.32fF
C15109 a_11067_21583# a_12166_21501# 0.32fF
C15110 a_5254_67503# a_3295_62083# 0.53fF
C15111 a_22127_37737# VDD 0.60fF
C15112 vcm_commonmode a_33338_20902# 0.31fF
C15113 vcm_commonmode a_22294_63198# 0.31fF
C15114 a_21290_68218# a_21382_68218# 0.32fF
C15115 a_2289_35113# a_2503_34319# 0.56fF
C15116 a_4758_45369# a_1761_46287# 0.76fF
C15117 a_1823_58773# VDD 1.75fF
C15118 a_43470_8488# a_43470_7484# 1.00fF
C15119 a_20378_7484# a_21382_7484# 0.97fF
C15120 vcm_commonmode a_16362_9492# 4.47fF
C15121 a_35438_58178# ctopp 3.59fF
C15122 a_11067_66191# a_5039_42167# 0.37fF
C15123 a_49494_66210# VDD 1.10fF
C15124 vcm_commonmode a_32426_16520# 0.87fF
C15125 ctopn a_18370_13508# 3.58fF
C15126 a_17507_52047# a_34145_49007# 0.60fF
C15127 a_23736_7638# a_10515_23975# 0.41fF
C15128 vcm_commonmode a_12901_58799# 6.22fF
C15129 a_4443_46607# a_5715_44343# 0.87fF
C15130 a_7295_44647# a_18979_30287# 3.54fF
C15131 a_26402_12504# VDD 0.51fF
C15132 a_32327_40191# VDD 1.71fF
C15133 a_1895_18756# VDD 0.58fF
C15134 a_19720_7638# a_12985_16367# 0.41fF
C15135 a_1761_39215# a_13097_36367# 0.39fF
C15136 a_31422_9492# a_32426_9492# 0.97fF
C15137 vcm_commonmode a_33338_12870# 0.31fF
C15138 a_32772_7638# a_12546_22351# 0.41fF
C15139 a_32426_13508# a_32426_12504# 1.00fF
C15140 a_13716_43047# a_12663_40871# 0.63fF
C15141 a_39389_52271# a_39454_63198# 0.42fF
C15142 a_47486_16520# a_48490_16520# 0.97fF
C15143 a_21371_50959# a_25398_69222# 0.38fF
C15144 a_21382_21540# VDD 0.51fF
C15145 vcm_commonmode a_24394_7484# 0.69fF
C15146 a_41261_28335# ctopn 4.67fF
C15147 a_8491_27023# a_2143_15271# 1.30fF
C15148 a_3143_66972# a_6737_60431# 0.49fF
C15149 a_11067_67279# a_33864_28111# 0.41fF
C15150 vcm_commonmode a_28318_21906# 0.31fF
C15151 a_22386_69222# ctopp 3.59fF
C15152 a_7736_10499# VDD 0.70fF
C15153 vcm_commonmode a_18370_64202# 0.88fF
C15154 vcm_commonmode a_46390_58178# 0.31fF
C15155 a_26402_17524# VDD 0.51fF
C15156 a_26155_50095# VDD 0.49fF
C15157 a_40366_72234# a_40458_72234# 0.32fF
C15158 a_12727_58255# a_16362_60186# 19.89fF
C15159 a_11067_47695# a_8295_47388# 4.51fF
C15160 a_32426_55166# a_33430_55166# 0.97fF
C15161 a_16510_8760# a_12877_14441# 1.08fF
C15162 a_2840_53511# a_3295_62083# 0.30fF
C15163 a_32367_28309# VDD 2.92fF
C15164 vcm_commonmode a_33338_17890# 0.31fF
C15165 a_20378_65206# ctopp 3.59fF
C15166 a_1644_74005# VDD 0.32fF
C15167 a_29760_55394# a_12981_59343# 0.40fF
C15168 vcm_commonmode a_20286_60186# 0.31fF
C15169 a_22386_67214# a_22386_66210# 1.00fF
C15170 a_1586_9991# a_3247_10389# 0.79fF
C15171 a_1586_40455# config_2_in[11] 0.67fF
C15172 a_10394_19605# VDD 1.10fF
C15173 a_36797_27497# a_37446_18528# 0.38fF
C15174 a_24959_30503# a_32038_29575# 0.52fF
C15175 a_18370_65206# a_18370_64202# 1.00fF
C15176 a_35346_13874# a_35438_13508# 0.32fF
C15177 a_18151_52263# a_24394_55166# 0.46fF
C15178 a_24800_43041# a_34222_43439# 0.46fF
C15179 a_40366_68218# a_40458_68218# 0.32fF
C15180 a_17039_51157# a_23763_47381# 0.70fF
C15181 a_5805_15279# VDD 0.59fF
C15182 a_41872_29423# a_12516_7093# 0.40fF
C15183 vcm_commonmode a_27406_69222# 0.87fF
C15184 a_47486_59182# VDD 0.51fF
C15185 a_39454_7484# a_40458_7484# 0.97fF
C15186 a_20267_30503# a_7939_30503# 1.63fF
C15187 a_26523_29199# VDD 7.82fF
C15188 a_21290_56170# a_21382_56170# 0.32fF
C15189 a_2840_66103# a_8999_61493# 0.38fF
C15190 a_11067_67279# a_42709_29199# 0.40fF
C15191 vcm_commonmode a_34434_22544# 0.87fF
C15192 a_23395_32463# a_30891_28309# 0.34fF
C15193 a_9219_11471# VDD 1.52fF
C15194 a_6473_40277# VDD 1.48fF
C15195 vcm_commonmode a_25398_65206# 0.87fF
C15196 a_23390_69222# a_24394_69222# 0.97fF
C15197 a_23749_36929# a_24055_36415# 0.30fF
C15198 a_27406_18528# VDD 0.51fF
C15199 a_40491_27247# a_12985_16367# 0.41fF
C15200 a_39673_28111# a_40458_16520# 0.38fF
C15201 a_6372_38279# a_6662_34025# 0.74fF
C15202 a_18370_61190# a_18370_60186# 1.00fF
C15203 ctopn a_25398_8488# 3.40fF
C15204 a_37919_28111# a_12546_22351# 0.41fF
C15205 a_33430_64202# a_34434_64202# 0.97fF
C15206 vcm_commonmode a_34342_18894# 0.31fF
C15207 a_27406_66210# ctopp 3.59fF
C15208 a_11067_46823# a_18979_30287# 1.36fF
C15209 a_12895_13967# a_12899_10927# 23.48fF
C15210 a_19478_51959# a_20535_51727# 0.51fF
C15211 a_18370_55166# VDD 0.61fF
C15212 a_31768_7638# a_12877_16911# 0.41fF
C15213 a_30418_22544# a_31422_22544# 0.97fF
C15214 a_8132_53511# VDD 2.80fF
C15215 vcm_commonmode a_30418_14512# 0.87fF
C15216 a_14287_51175# a_7295_44647# 5.11fF
C15217 a_21382_65206# a_22386_65206# 0.97fF
C15218 a_35647_38053# VDD 0.86fF
C15219 a_11067_67279# a_9503_26151# 0.44fF
C15220 vcm_commonmode a_25306_55166# 0.30fF
C15221 a_36442_10496# VDD 0.51fF
C15222 a_17366_17524# a_17366_16520# 1.00fF
C15223 vcm_commonmode a_12947_56817# 1.43fF
C15224 a_1761_35407# a_1761_34319# 1.20fF
C15225 a_1761_27791# a_6243_30662# 0.46fF
C15226 vcm_commonmode a_43378_10862# 0.31fF
C15227 a_16863_29415# a_28757_27247# 0.72fF
C15228 a_21382_56170# a_21382_55166# 1.00fF
C15229 a_25263_29981# VDD 1.94fF
C15230 a_17507_52047# a_30928_49007# 1.00fF
C15231 a_1950_59887# VDD 8.68fF
C15232 a_13183_52047# a_12727_58255# 0.40fF
C15233 a_41462_67214# a_41462_66210# 1.00fF
C15234 vcm_commonmode a_35438_23548# 0.87fF
C15235 a_30418_7484# m3_30320_7346# 2.80fF
C15236 a_4535_43031# VDD 0.31fF
C15237 vcm_commonmode a_32426_66210# 0.87fF
C15238 a_13123_38231# a_13743_35836# 0.42fF
C15239 a_2775_46025# a_1761_50639# 0.67fF
C15240 a_30764_7638# a_12877_16911# 0.41fF
C15241 a_23390_62194# VDD 0.51fF
C15242 a_20286_61190# a_20378_61190# 0.32fF
C15243 a_37446_65206# a_37446_64202# 1.00fF
C15244 vcm_commonmode a_44474_19532# 0.87fF
C15245 ctopn a_26402_16520# 3.59fF
C15246 vcm_commonmode a_30326_62194# 0.31fF
C15247 a_11067_46823# a_37427_47893# 0.61fF
C15248 a_31422_15516# VDD 0.51fF
C15249 a_31186_48169# VDD 0.50fF
C15250 a_21382_19532# a_22386_19532# 0.97fF
C15251 vcm_commonmode a_16510_8760# 19.82fF
C15252 a_5535_18012# VDD 3.85fF
C15253 m3_49396_7346# VDD 0.50fF
C15254 a_31422_23548# a_31422_22544# 1.00fF
C15255 vcm_commonmode a_38358_15882# 0.31fF
C15256 a_31422_63198# ctopp 3.64fF
C15257 a_12899_3311# a_12341_3311# 0.83fF
C15258 a_40366_56170# a_40458_56170# 0.32fF
C15259 a_29414_71230# VDD 0.58fF
C15260 vcm_commonmode a_16362_58178# 4.47fF
C15261 a_25398_66210# a_25398_65206# 1.00fF
C15262 a_29072_38567# VDD 1.58fF
C15263 a_26402_14512# a_27406_14512# 0.97fF
C15264 a_2656_45895# a_2539_42106# 0.49fF
C15265 a_4563_32900# a_3987_19623# 0.93fF
C15266 a_1761_50639# a_19919_38695# 0.72fF
C15267 a_41462_11500# VDD 0.51fF
C15268 a_30855_41809# VDD 2.31fF
C15269 a_42466_69222# a_43470_69222# 0.97fF
C15270 a_1591_16917# VDD 0.72fF
C15271 vcm_commonmode a_36350_71230# 0.31fF
C15272 a_37446_61190# a_37446_60186# 1.00fF
C15273 a_23298_8854# a_23390_8488# 0.32fF
C15274 a_45478_24552# VDD 0.60fF
C15275 vcm_commonmode a_48398_11866# 0.31fF
C15276 a_25398_59182# ctopp 3.59fF
C15277 a_6095_44807# a_12202_54599# 0.69fF
C15278 a_23395_52047# a_2959_47113# 0.44fF
C15279 a_23395_32463# a_30052_32117# 0.31fF
C15280 a_13643_28327# a_12447_29199# 0.61fF
C15281 a_2292_43291# a_6559_45205# 0.56fF
C15282 a_25971_52263# a_30418_68218# 0.38fF
C15283 a_24302_70226# a_24394_70226# 0.32fF
C15284 a_41370_58178# a_41462_58178# 0.32fF
C15285 a_5599_74549# a_1586_69367# 0.39fF
C15286 a_40675_27791# a_41462_18528# 0.38fF
C15287 a_17712_7638# a_17366_18528# 0.38fF
C15288 a_23390_62194# a_23390_61190# 1.00fF
C15289 a_47486_57174# VDD 0.51fF
C15290 a_40458_65206# a_41462_65206# 0.97fF
C15291 vcm_commonmode a_47486_20536# 0.87fF
C15292 vcm_commonmode a_36442_63198# 0.92fF
C15293 a_36442_17524# a_36442_16520# 1.00fF
C15294 a_22843_29415# a_15607_46805# 1.03fF
C15295 a_1761_52815# a_2927_39733# 1.64fF
C15296 a_40050_48463# a_45478_71230# 0.38fF
C15297 a_23390_20536# a_23390_19532# 1.00fF
C15298 m3_34336_72146# VDD 0.33fF
C15299 a_31422_23548# a_32426_23548# 0.97fF
C15300 a_9263_24501# a_10275_21495# 0.58fF
C15301 a_5239_65301# VDD 0.58fF
C15302 a_34434_72234# VDD 1.37fF
C15303 a_28756_55394# a_28410_60186# 0.38fF
C15304 a_28410_66210# a_29414_66210# 0.97fF
C15305 a_36613_48169# a_12727_58255# 0.40fF
C15306 vcm_commonmode a_30418_59182# 0.87fF
C15307 vcm_commonmode m3_16264_69134# 3.21fF
C15308 a_18627_42943# VDD 0.84fF
C15309 a_14287_51175# a_12355_65103# 0.89fF
C15310 a_4351_67279# a_8772_63927# 0.39fF
C15311 a_39299_48783# a_44474_67214# 0.38fF
C15312 a_13097_37455# a_1761_35407# 0.35fF
C15313 a_35568_49525# VDD 2.10fF
C15314 vcm_commonmode a_39454_72234# 0.69fF
C15315 a_39673_28111# a_12727_13353# 0.41fF
C15316 a_39362_61190# a_39454_61190# 0.32fF
C15317 vcm_commonmode a_47486_12504# 0.87fF
C15318 a_29414_60186# ctopp 3.59fF
C15319 ctopn a_48490_9492# 3.42fF
C15320 a_32426_68218# VDD 0.51fF
C15321 a_32334_7850# VDD 0.62fF
C15322 a_25971_52263# a_30418_56170# 0.38fF
C15323 ctopn a_28410_22544# 3.58fF
C15324 vcm_commonmode a_39362_68218# 0.31fF
C15325 a_28410_71230# a_28410_70226# 1.00fF
C15326 a_40458_19532# a_41462_19532# 0.97fF
C15327 a_4674_40277# a_18328_31573# 0.88fF
C15328 a_34482_29941# a_26523_29199# 0.33fF
C15329 a_8491_41383# a_33694_30761# 1.08fF
C15330 a_41872_29423# a_15607_46805# 0.32fF
C15331 a_15189_39889# a_12889_39889# 0.87fF
C15332 a_2952_66139# VDD 5.18fF
C15333 a_44474_66210# a_44474_65206# 1.00fF
C15334 a_33727_38825# VDD 0.64fF
C15335 a_45478_14512# a_46482_14512# 0.97fF
C15336 vcm_commonmode a_42466_21540# 0.87fF
C15337 a_1586_9991# a_4429_14191# 0.39fF
C15338 a_1895_49722# VDD 0.78fF
C15339 a_8575_74853# a_10699_69679# 0.36fF
C15340 a_24394_20536# a_25398_20536# 0.97fF
C15341 a_25744_7638# a_12877_14441# 0.41fF
C15342 a_42374_8854# a_42466_8488# 0.32fF
C15343 vcm_commonmode a_19374_10496# 0.87fF
C15344 a_11710_58487# a_11883_58575# 0.32fF
C15345 vcm_commonmode a_47486_17524# 0.87fF
C15346 ctopn a_24394_14512# 3.59fF
C15347 a_3137_73493# VDD 0.70fF
C15348 vcm_commonmode a_34434_60186# 0.87fF
C15349 a_46482_13508# VDD 0.51fF
C15350 a_4535_43567# VDD 0.47fF
C15351 a_43378_70226# a_43470_70226# 0.32fF
C15352 a_40675_27791# a_12899_11471# 0.41fF
C15353 a_42466_62194# a_42466_61190# 1.00fF
C15354 a_33430_10496# a_33430_9492# 1.00fF
C15355 a_32426_56170# VDD 0.52fF
C15356 a_10055_58791# a_36629_27791# 0.41fF
C15357 a_39673_28111# a_10515_23975# 0.41fF
C15358 a_20563_36649# VDD 0.56fF
C15359 a_11067_13095# a_6835_46823# 0.83fF
C15360 m2_48260_24282# m3_48392_24414# 0.85fF
C15361 a_24302_16886# a_24394_16520# 0.32fF
C15362 vcm_commonmode a_39362_56170# 0.31fF
C15363 ctopn a_29414_23548# 3.40fF
C15364 a_9865_14441# VDD 0.57fF
C15365 a_42466_20536# a_42466_19532# 1.00fF
C15366 vcm_commonmode a_22294_8854# 0.31fF
C15367 a_10975_66407# a_9275_15253# 0.30fF
C15368 a_3339_32463# a_3339_30503# 0.60fF
C15369 a_25398_57174# ctopp 3.58fF
C15370 a_47486_66210# a_48490_66210# 0.97fF
C15371 ctopn a_38450_19532# 3.59fF
C15372 vcm_commonmode m3_16264_16382# 3.21fF
C15373 a_36579_42359# VDD 0.62fF
C15374 a_35676_49525# VDD 1.56fF
C15375 a_25744_7638# a_25398_16520# 0.38fF
C15376 a_22386_21540# a_22386_20536# 1.00fF
C15377 a_8491_27023# a_18370_16520# 0.38fF
C15378 a_31422_61190# VDD 0.51fF
C15379 vcm_commonmode a_24394_11500# 0.87fF
C15380 a_24394_12504# a_25398_12504# 0.97fF
C15381 vcm_commonmode a_48490_18528# 0.87fF
C15382 a_13390_29575# a_18126_28023# 0.53fF
C15383 a_12663_40871# a_32327_40191# 0.73fF
C15384 vcm_commonmode a_38358_61190# 0.31fF
C15385 a_30326_67214# a_30418_67214# 0.32fF
C15386 vcm_commonmode a_28410_24552# 0.84fF
C15387 a_14287_51175# ctopp 2.61fF
C15388 m2_48260_54946# inp_analog 0.75fF
C15389 a_47486_71230# a_47486_70226# 1.00fF
C15390 a_32426_55166# VDD 0.60fF
C15391 a_12546_22351# a_12166_21501# 0.45fF
C15392 a_6835_46823# a_23830_49525# 0.88fF
C15393 a_39454_62194# ctopp 3.59fF
C15394 a_35438_70226# VDD 0.51fF
C15395 vcm_commonmode a_38450_55166# 0.84fF
C15396 a_30115_38695# VDD 2.18fF
C15397 a_12727_67753# a_16362_68218# 19.89fF
C15398 vcm_commonmode a_30418_57174# 0.87fF
C15399 a_26397_51183# a_26417_47919# 0.55fF
C15400 a_20359_29199# a_16863_29415# 1.05fF
C15401 a_16746_16518# VDD 33.21fF
C15402 vcm_commonmode a_42374_70226# 0.31fF
C15403 a_43470_20536# a_44474_20536# 0.97fF
C15404 a_2775_46025# a_4482_57863# 0.94fF
C15405 a_16270_7850# a_16362_7484# 0.33fF
C15406 VDD config_1_in[5] 0.96fF
C15407 a_32426_63198# a_33430_63198# 0.97fF
C15408 vcm_commonmode a_23298_16886# 0.31fF
C15409 a_45478_71230# ctopp 3.40fF
C15410 ctopn a_41462_20536# 3.59fF
C15411 a_27183_43493# VDD 0.93fF
C15412 a_32334_58178# a_32426_58178# 0.32fF
C15413 a_19374_21540# a_20378_21540# 0.97fF
C15414 a_24683_27497# VDD 0.45fF
C15415 a_27314_9858# a_27406_9492# 0.32fF
C15416 a_12202_54599# VDD 1.22fF
C15417 a_7624_68021# VDD 0.32fF
C15418 a_43267_31055# a_46482_55166# 0.55fF
C15419 a_34251_52263# a_35438_63198# 0.42fF
C15420 vcm_commonmode a_44474_62194# 0.87fF
C15421 a_43378_16886# a_43470_16520# 0.32fF
C15422 vcm_commonmode a_25744_7638# 10.35fF
C15423 a_12901_66665# a_16362_70226# 1.15fF
C15424 a_17507_52047# a_21382_69222# 0.38fF
C15425 a_1586_18695# a_1757_18543# 0.60fF
C15426 a_24394_58178# VDD 0.51fF
C15427 a_26402_59182# a_27406_59182# 0.97fF
C15428 a_13669_38517# a_13909_38659# 0.56fF
C15429 a_33864_28111# a_34434_19532# 0.38fF
C15430 ctopn a_41462_12504# 3.59fF
C15431 a_3949_41935# a_1761_39215# 0.31fF
C15432 a_5490_41365# a_3305_38671# 1.45fF
C15433 vcm_commonmode a_31330_58178# 0.31fF
C15434 a_40050_48463# a_12901_58799# 0.40fF
C15435 a_24394_17524# a_25398_17524# 0.97fF
C15436 a_27535_30503# a_21187_29415# 1.03fF
C15437 a_41462_21540# a_41462_20536# 1.00fF
C15438 a_3339_43023# a_4443_46607# 1.46fF
C15439 a_28410_24552# a_28410_23548# 1.00fF
C15440 a_30764_7638# a_30418_22544# 0.38fF
C15441 a_41462_67214# VDD 0.51fF
C15442 a_13643_28327# a_11067_23759# 0.35fF
C15443 a_43470_12504# a_44474_12504# 0.97fF
C15444 a_5441_72399# VDD 1.04fF
C15445 a_17599_52263# a_12981_59343# 0.40fF
C15446 a_49402_67214# a_49494_67214# 0.32fF
C15447 ctopn a_36442_21540# 3.59fF
C15448 vcm_commonmode a_48398_67214# 0.31fF
C15449 a_1591_51183# a_1757_51183# 0.69fF
C15450 a_2775_46025# a_32582_51701# 0.82fF
C15451 a_2473_34293# config_2_in[3] 0.70fF
C15452 a_1591_54447# VDD 1.07fF
C15453 vcm_commonmode a_29414_13508# 0.87fF
C15454 a_38557_32143# a_18979_30287# 2.43fF
C15455 a_31768_7638# a_31422_23548# 0.38fF
C15456 a_3305_38671# a_4941_35727# 0.52fF
C15457 a_12907_56399# a_4891_47388# 0.48fF
C15458 a_48490_68218# ctopp 3.43fF
C15459 ctopn a_41462_17524# 3.59fF
C15460 a_16955_52047# a_20378_55166# 0.47fF
C15461 a_38450_9492# VDD 0.51fF
C15462 a_42985_46831# a_12355_15055# 0.40fF
C15463 a_11067_67279# a_3339_30503# 0.57fF
C15464 a_36717_47375# a_12516_7093# 0.40fF
C15465 vcm_commonmode a_18278_69222# 0.31fF
C15466 a_9503_26151# a_20378_14512# 0.38fF
C15467 a_35346_7850# a_35438_7484# 0.32fF
C15468 a_18370_22544# VDD 0.52fF
C15469 vcm_commonmode a_45386_9858# 0.31fF
C15470 a_1689_10396# a_2011_34837# 0.31fF
C15471 a_9204_30663# VDD 0.30fF
C15472 a_39223_32463# a_11067_21583# 0.41fF
C15473 a_2315_24540# a_3325_18543# 0.88fF
C15474 a_16746_56172# a_16362_56170# 2.28fF
C15475 a_45386_72234# VDD 0.63fF
C15476 vcm_commonmode a_25306_22910# 0.31fF
C15477 a_7155_55509# a_7479_54439# 0.71fF
C15478 a_14926_31849# a_17358_31069# 1.21fF
C15479 a_12343_42333# VDD 2.07fF
C15480 a_19282_69222# a_19374_69222# 0.32fF
C15481 a_25398_18528# a_25398_17524# 1.00fF
C15482 a_38450_21540# a_39454_21540# 0.97fF
C15483 a_5411_59317# VDD 0.44fF
C15484 a_46390_9858# a_46482_9492# 0.32fF
C15485 a_29322_64202# a_29414_64202# 0.32fF
C15486 a_7580_61751# a_7519_59575# 0.58fF
C15487 a_46482_7484# VDD 1.35fF
C15488 ctopn m3_48392_24414# 0.35fF
C15489 a_45478_59182# a_46482_59182# 0.97fF
C15490 a_26310_22910# a_26402_22544# 0.32fF
C15491 a_40458_64202# VDD 0.51fF
C15492 a_1643_56597# VDD 0.35fF
C15493 vcm_commonmode a_21290_14878# 0.31fF
C15494 ctopn a_18370_11500# 3.58fF
C15495 a_48490_56170# ctopp 3.46fF
C15496 a_17274_65206# a_17366_65206# 0.32fF
C15497 a_14031_38007# VDD 0.59fF
C15498 a_26402_14512# a_26402_13508# 1.00fF
C15499 ctopn a_42466_18528# 3.59fF
C15500 a_6559_45205# a_6725_45205# 0.42fF
C15501 a_32121_40741# VDD 1.87fF
C15502 vcm_commonmode a_47394_64202# 0.31fF
C15503 a_43470_17524# a_44474_17524# 0.97fF
C15504 a_14831_50095# a_32134_49159# 0.31fF
C15505 a_15103_49525# VDD 0.49fF
C15506 vcm_commonmode a_18370_70226# 0.88fF
C15507 a_1923_54591# a_1591_51183# 0.34fF
C15508 a_30418_60186# a_31422_60186# 0.97fF
C15509 a_19374_23548# VDD 0.52fF
C15510 a_47486_24552# a_47486_23548# 1.00fF
C15511 a_16746_66212# VDD 33.19fF
C15512 a_5547_31599# VDD 0.49fF
C15513 a_32426_12504# a_32426_11500# 1.00fF
C15514 a_1761_43567# a_19245_39747# 0.53fF
C15515 a_6921_72943# VDD 1.87fF
C15516 vcm_commonmode a_26310_23914# 0.31fF
C15517 a_23390_7484# m3_23292_7346# 2.80fF
C15518 a_29391_44031# VDD 0.84fF
C15519 vcm_commonmode a_23298_66210# 0.31fF
C15520 a_19374_70226# a_19374_69222# 1.00fF
C15521 a_25398_18528# a_26402_18528# 0.97fF
C15522 a_28410_19532# VDD 0.51fF
C15523 a_32772_7638# a_12985_16367# 0.41fF
C15524 a_1761_40847# a_13669_35253# 1.22fF
C15525 a_47486_61190# ctopp 3.58fF
C15526 a_16510_8760# a_12899_11471# 1.08fF
C15527 a_13909_39747# a_1761_27791# 5.71fF
C15528 a_49494_69222# VDD 1.24fF
C15529 vcm_commonmode a_35346_19898# 0.31fF
C15530 a_19374_67214# ctopp 3.59fF
C15531 a_43362_28879# a_12257_56623# 0.40fF
C15532 a_2292_43291# a_1761_47919# 0.32fF
C15533 a_27535_30503# a_26523_28111# 3.52fF
C15534 a_12489_47919# VDD 0.62fF
C15535 a_17274_19898# a_17366_19532# 0.32fF
C15536 a_6559_22671# a_10073_23439# 0.51fF
C15537 vcm_commonmode a_36442_8488# 0.86fF
C15538 m3_21284_7346# VDD 0.39fF
C15539 a_47486_65206# VDD 0.51fF
C15540 a_18370_11500# a_18370_10496# 1.00fF
C15541 a_41261_28335# a_10515_22671# 0.40fF
C15542 a_22294_14878# a_22386_14512# 0.32fF
C15543 a_19967_41781# VDD 7.31fF
C15544 a_2191_68565# a_1954_61677# 0.90fF
C15545 a_38358_69222# a_38450_69222# 0.32fF
C15546 a_44474_18528# a_44474_17524# 1.00fF
C15547 a_2595_47653# a_1586_40455# 0.44fF
C15548 a_27406_72234# a_28410_72234# 0.97fF
C15549 a_36350_24918# VDD 0.36fF
C15550 a_12901_58799# ctopp 3.23fF
C15551 a_5531_22895# a_6451_22895# 0.40fF
C15552 a_9135_27239# a_21382_22544# 0.38fF
C15553 a_48398_64202# a_48490_64202# 0.32fF
C15554 a_8461_32937# VDD 1.50fF
C15555 ctopn a_46482_15516# 3.59fF
C15556 a_12516_7093# a_8295_47388# 0.74fF
C15557 a_3247_20495# a_2339_38129# 0.66fF
C15558 a_3019_13621# a_2873_13879# 0.90fF
C15559 a_7939_30503# a_10506_29967# 1.50fF
C15560 a_18703_29199# a_7295_44647# 6.01fF
C15561 a_1689_10396# VDD 13.96fF
C15562 vcm_commonmode a_24394_67214# 0.87fF
C15563 a_21371_52263# a_26402_68218# 0.38fF
C15564 a_18611_52047# a_2235_30503# 2.10fF
C15565 a_8295_47388# a_2606_41079# 3.80fF
C15566 a_31422_20536# VDD 0.51fF
C15567 a_46390_55166# VDD 0.35fF
C15568 a_41967_31375# a_42466_15516# 0.38fF
C15569 a_45386_22910# a_45478_22544# 0.32fF
C15570 a_36629_27791# a_36442_18528# 0.38fF
C15571 a_20378_63198# VDD 0.57fF
C15572 a_24959_30503# a_30565_30199# 0.32fF
C15573 a_34434_10496# a_35438_10496# 0.97fF
C15574 a_36350_65206# a_36442_65206# 0.32fF
C15575 a_7155_55509# a_9526_61751# 0.53fF
C15576 a_29679_37737# VDD 0.63fF
C15577 a_45478_14512# a_45478_13508# 1.00fF
C15578 vcm_commonmode a_38358_20902# 0.31fF
C15579 vcm_commonmode a_27314_63198# 0.31fF
C15580 a_24683_48463# VDD 0.32fF
C15581 a_41427_52263# a_41462_71230# 0.38fF
C15582 vcm_commonmode a_21382_9492# 0.87fF
C15583 a_27314_23914# a_27406_23548# 0.32fF
C15584 a_31768_7638# a_12895_13967# 0.41fF
C15585 a_11067_47695# a_11619_3303# 0.73fF
C15586 a_20378_11500# a_21382_11500# 0.97fF
C15587 vcm_commonmode a_37446_16520# 0.87fF
C15588 a_18370_64202# ctopp 3.58fF
C15589 ctopn a_23390_13508# 3.59fF
C15590 a_12671_42134# a_12473_41781# 0.30fF
C15591 a_27406_72234# VDD 1.23fF
C15592 a_18151_52263# a_24394_60186# 0.38fF
C15593 a_24302_66210# a_24394_66210# 0.32fF
C15594 a_25971_52263# a_12727_58255# 0.40fF
C15595 vcm_commonmode a_21290_59182# 0.31fF
C15596 a_7281_29423# a_4427_30511# 0.42fF
C15597 a_31422_12504# VDD 0.51fF
C15598 a_2004_42453# VDD 9.10fF
C15599 a_39222_48169# a_40458_67214# 0.38fF
C15600 a_3143_66972# a_5024_67885# 0.98fF
C15601 a_38450_70226# a_38450_69222# 1.00fF
C15602 a_32772_7638# a_32426_9492# 0.38fF
C15603 a_44474_18528# a_45478_18528# 0.97fF
C15604 a_27627_51733# VDD 0.34fF
C15605 vcm_commonmode a_32426_72234# 0.69fF
C15606 a_37919_28111# a_12985_16367# 0.41fF
C15607 a_49494_55166# m3_49396_55078# 2.81fF
C15608 vcm_commonmode a_38358_12870# 0.31fF
C15609 a_24394_24552# a_25398_24552# 0.97fF
C15610 a_21371_52263# a_26402_56170# 0.38fF
C15611 a_36350_19898# a_36442_19532# 0.32fF
C15612 a_1803_20719# a_1761_25615# 0.39fF
C15613 a_26402_21540# VDD 0.51fF
C15614 vcm_commonmode a_29414_7484# 0.69fF
C15615 a_30764_7638# a_12895_13967# 0.41fF
C15616 a_16362_64202# VDD 2.48fF
C15617 a_2787_32679# a_6243_30662# 1.46fF
C15618 a_22843_29415# a_28841_29575# 0.46fF
C15619 a_4314_40821# a_5993_37039# 0.33fF
C15620 a_18979_30287# a_30155_32375# 0.73fF
C15621 a_21382_62194# a_22386_62194# 0.97fF
C15622 a_37446_11500# a_37446_10496# 1.00fF
C15623 a_4497_29673# VDD 0.34fF
C15624 a_44474_58178# VDD 0.51fF
C15625 a_41370_14878# a_41462_14512# 0.32fF
C15626 a_17799_38591# VDD 0.86fF
C15627 vcm_commonmode a_33338_21906# 0.31fF
C15628 a_27406_69222# ctopp 3.59fF
C15629 a_3339_43023# a_13097_36367# 3.76fF
C15630 a_40921_41245# VDD 1.06fF
C15631 vcm_commonmode a_23390_64202# 0.87fF
C15632 a_1761_31055# a_1761_32143# 1.14fF
C15633 a_32327_35839# a_13669_35253# 0.79fF
C15634 a_31422_17524# VDD 0.51fF
C15635 a_41261_28335# a_42466_72234# 0.34fF
C15636 a_20286_20902# a_20378_20536# 0.32fF
C15637 a_18370_60186# VDD 0.52fF
C15638 a_34434_55166# a_35438_55166# 0.97fF
C15639 a_11067_63143# a_8295_47388# 0.33fF
C15640 a_23736_7638# a_23390_18528# 0.38fF
C15641 a_3339_32463# a_2473_34293# 0.71fF
C15642 a_7676_61493# a_7523_62581# 0.60fF
C15643 a_11067_13095# a_5085_24759# 0.43fF
C15644 vcm_commonmode a_38358_17890# 0.31fF
C15645 a_25398_65206# ctopp 3.59fF
C15646 a_28305_28879# a_31768_7638# 0.38fF
C15647 a_26402_57174# a_27406_57174# 0.97fF
C15648 vcm_commonmode a_25306_60186# 0.31fF
C15649 a_29414_15516# a_30418_15516# 0.97fF
C15650 a_8295_47388# a_16753_49007# 0.62fF
C15651 a_2959_47113# a_16385_51183# 0.59fF
C15652 a_13669_39605# a_12473_37429# 2.12fF
C15653 a_1761_39215# a_1761_37039# 1.09fF
C15654 a_22291_29415# a_33839_28309# 0.45fF
C15655 a_7598_36103# VDD 2.11fF
C15656 a_1761_44111# a_20899_44211# 0.78fF
C15657 a_11067_46823# a_18703_29199# 1.28fF
C15658 a_5755_14709# VDD 1.00fF
C15659 a_27406_71230# a_28410_71230# 0.97fF
C15660 vcm_commonmode a_32426_69222# 0.87fF
C15661 a_2143_15271# a_1586_9991# 0.43fF
C15662 a_3339_43023# a_4500_45289# 0.39fF
C15663 a_46390_23914# a_46482_23548# 0.32fF
C15664 a_24959_30503# a_32367_28309# 1.36fF
C15665 a_39454_11500# a_40458_11500# 0.97fF
C15666 a_12947_56817# ctopp 1.43fF
C15667 a_13183_52047# a_17366_59182# 0.38fF
C15668 a_43378_66210# a_43470_66210# 0.32fF
C15669 vcm_commonmode a_39454_22544# 0.87fF
C15670 a_10531_31055# a_14361_29967# 0.47fF
C15671 a_21479_42405# VDD 0.84fF
C15672 vcm_commonmode a_30418_65206# 0.87fF
C15673 a_43362_28879# a_10975_66407# 0.40fF
C15674 a_32426_18528# VDD 0.51fF
C15675 a_30947_51157# VDD 0.40fF
C15676 a_7203_24527# VDD 0.33fF
C15677 ctopn a_30418_8488# 3.40fF
C15678 a_43470_24552# a_44474_24552# 0.97fF
C15679 a_20286_12870# a_20378_12504# 0.32fF
C15680 vcm_commonmode a_39362_18894# 0.31fF
C15681 a_32426_66210# ctopp 3.59fF
C15682 vcm_commonmode a_19282_24918# 0.31fF
C15683 a_4495_35925# a_6649_25615# 0.86fF
C15684 a_23390_55166# VDD 0.60fF
C15685 a_24959_30503# a_26523_29199# 0.34fF
C15686 a_40458_62194# a_41462_62194# 0.97fF
C15687 a_1770_14441# config_2_in[10] 0.48fF
C15688 vcm_commonmode a_35438_14512# 0.87fF
C15689 a_4191_33449# a_5915_30287# 0.40fF
C15690 vcm_commonmode a_30326_55166# 0.30fF
C15691 a_41462_10496# VDD 0.51fF
C15692 a_13576_40413# VDD 2.53fF
C15693 vcm_commonmode a_21290_57174# 0.31fF
C15694 a_1761_52815# a_2952_46805# 0.42fF
C15695 a_41261_28335# a_12901_66665# 0.40fF
C15696 a_39362_20902# a_39454_20536# 0.32fF
C15697 vcm_commonmode a_48398_10862# 0.31fF
C15698 a_16362_58178# ctopp 1.35fF
C15699 a_28318_63198# a_28410_63198# 0.32fF
C15700 a_33798_31145# VDD 0.50fF
C15701 a_45478_57174# a_46482_57174# 0.97fF
C15702 a_19374_57174# a_19374_56170# 1.00fF
C15703 a_48490_15516# a_49494_15516# 0.97fF
C15704 vcm_commonmode a_40458_23548# 0.87fF
C15705 a_1761_11471# VDD 0.31fF
C15706 vcm_commonmode a_37446_66210# 0.87fF
C15707 a_19576_51701# VDD 1.10fF
C15708 a_6559_59663# a_6775_53877# 0.74fF
C15709 a_25744_7638# a_12899_11471# 0.41fF
C15710 a_26748_7638# a_26402_16520# 0.38fF
C15711 a_28410_62194# VDD 0.51fF
C15712 a_10055_58791# a_29760_7638# 0.41fF
C15713 a_11710_58487# a_11521_58951# 0.56fF
C15714 vcm_commonmode a_49494_19532# 0.96fF
C15715 ctopn a_31422_16520# 3.59fF
C15716 a_41261_28335# a_42466_55166# 0.45fF
C15717 a_31768_55394# a_31422_63198# 0.42fF
C15718 vcm_commonmode a_35346_62194# 0.31fF
C15719 a_36442_15516# VDD 0.51fF
C15720 a_46482_71230# a_47486_71230# 0.97fF
C15721 a_22294_59182# a_22386_59182# 0.32fF
C15722 a_75794_38962# a_76346_38962# 0.57fF
C15723 a_2124_64507# VDD 0.69fF
C15724 a_5831_39189# a_16917_31573# 0.67fF
C15725 vcm_commonmode a_43378_15882# 0.31fF
C15726 a_36442_63198# ctopp 3.64fF
C15727 a_1761_41935# a_13909_39747# 1.05fF
C15728 a_34434_71230# VDD 0.58fF
C15729 a_1761_52815# a_1761_35407# 3.13fF
C15730 a_38557_32143# a_12901_58799# 0.40fF
C15731 a_38101_38565# VDD 1.62fF
C15732 a_46482_11500# VDD 0.51fF
C15733 a_20286_17890# a_20378_17524# 0.32fF
C15734 a_1761_31055# a_12663_35431# 2.16fF
C15735 a_7571_16917# VDD 0.44fF
C15736 a_33338_72234# a_33430_72234# 0.32fF
C15737 vcm_commonmode a_41370_71230# 0.31fF
C15738 a_36629_27791# a_12877_14441# 0.41fF
C15739 a_15607_46805# a_17712_7638# 0.52fF
C15740 a_6467_55527# a_4674_57685# 0.35fF
C15741 a_30418_59182# ctopp 3.59fF
C15742 a_42718_27497# a_11067_21583# 0.41fF
C15743 a_25419_50959# a_26523_29199# 1.31fF
C15744 a_27535_30503# a_35815_31751# 0.42fF
C15745 a_26402_64202# a_26402_63198# 1.23fF
C15746 a_39362_12870# a_39454_12504# 0.32fF
C15747 a_12663_40871# a_12343_42333# 0.58fF
C15748 a_12257_56623# a_16362_57174# 19.89fF
C15749 a_9227_12015# VDD 0.67fF
C15750 a_10883_18543# a_11049_18543# 0.69fF
C15751 a_34434_59182# a_34434_58178# 1.00fF
C15752 ctopn m2_48260_24282# 1.16fF
C15753 a_2124_54715# VDD 0.67fF
C15754 a_18370_22544# a_18370_21540# 1.00fF
C15755 a_1761_39215# a_13557_37999# 0.42fF
C15756 vcm_commonmode a_20286_13874# 0.31fF
C15757 a_5085_23047# a_5531_22895# 0.48fF
C15758 a_1761_50639# a_1761_35407# 1.43fF
C15759 a_25398_13508# a_26402_13508# 0.97fF
C15760 a_7381_35407# VDD 0.40fF
C15761 a_7841_12167# a_5671_21495# 0.39fF
C15762 a_1761_27791# VDD 8.31fF
C15763 a_30418_68218# a_31422_68218# 0.97fF
C15764 vcm_commonmode a_41462_63198# 0.92fF
C15765 a_41427_52263# a_12355_15055# 0.40fF
C15766 a_13183_52047# a_17366_57174# 0.38fF
C15767 a_16746_71232# a_12901_66665# 0.41fF
C15768 a_29760_55394# a_12516_7093# 0.40fF
C15769 m3_49396_72146# VDD 0.50fF
C15770 a_22843_29415# a_26523_29199# 0.39fF
C15771 a_42466_56170# a_42466_55166# 1.00fF
C15772 a_43470_24552# m3_43372_24414# 2.81fF
C15773 a_47394_63198# a_47486_63198# 0.32fF
C15774 a_39223_32463# a_12546_22351# 0.41fF
C15775 a_7841_12167# a_2292_17179# 1.04fF
C15776 a_38450_57174# a_38450_56170# 1.00fF
C15777 a_38358_72234# VDD 0.61fF
C15778 vcm_commonmode a_35438_59182# 0.87fF
C15779 a_23395_32463# a_26523_29199# 0.45fF
C15780 a_19004_40413# VDD 2.71fF
C15781 a_21371_52263# a_15548_30761# 0.34fF
C15782 a_34342_21906# a_34434_21540# 0.32fF
C15783 a_9751_25071# VDD 2.84fF
C15784 a_34434_60186# ctopp 3.59fF
C15785 a_5085_23047# a_7187_20719# 0.33fF
C15786 a_37446_68218# VDD 0.51fF
C15787 a_18811_34789# VDD 0.83fF
C15788 a_37354_7850# VDD 0.63fF
C15789 a_11803_55311# a_12981_62313# 1.07fF
C15790 a_22386_16520# a_22386_15516# 1.00fF
C15791 ctopn a_33430_22544# 3.59fF
C15792 vcm_commonmode a_44382_68218# 0.31fF
C15793 a_5190_59575# a_4482_57863# 0.81fF
C15794 a_41370_59182# a_41462_59182# 0.32fF
C15795 a_4758_45369# a_12755_53030# 0.66fF
C15796 a_4191_33449# a_5915_35943# 0.33fF
C15797 vcm_commonmode a_47486_21540# 0.87fF
C15798 a_18627_40767# VDD 0.89fF
C15799 a_5682_69367# a_7803_55509# 0.42fF
C15800 a_1950_59887# a_4339_64521# 0.34fF
C15801 a_39362_17890# a_39454_17524# 0.32fF
C15802 a_6725_49557# VDD 0.65fF
C15803 a_2419_48783# a_2872_44111# 0.94fF
C15804 a_26310_60186# a_26402_60186# 0.32fF
C15805 vcm_commonmode a_24394_10496# 0.87fF
C15806 a_4798_23759# a_8933_22583# 0.36fF
C15807 a_40675_27791# a_12985_7663# 0.41fF
C15808 a_15439_49525# a_16362_63198# 1.13fF
C15809 a_45478_64202# a_45478_63198# 1.23fF
C15810 ctopn a_29414_14512# 3.59fF
C15811 vcm_commonmode a_39454_60186# 0.87fF
C15812 vcm_commonmode a_16746_23546# 5.35fF
C15813 a_16362_7484# m3_16264_7346# 2.81fF
C15814 a_8583_33551# a_42165_36367# 1.19fF
C15815 a_21290_18894# a_21382_18528# 0.32fF
C15816 a_6559_59879# a_14983_51157# 0.77fF
C15817 a_37446_22544# a_37446_21540# 1.00fF
C15818 a_30023_41959# a_1761_32143# 0.37fF
C15819 a_27250_27791# VDD 0.70fF
C15820 a_37446_56170# VDD 0.52fF
C15821 a_44474_13508# a_45478_13508# 0.97fF
C15822 a_2099_59861# a_2011_34837# 1.79fF
C15823 a_20378_8488# VDD 0.58fF
C15824 a_12727_67753# a_12983_63151# 23.55fF
C15825 vcm_commonmode a_36629_27791# 10.35fF
C15826 vcm_commonmode a_44382_56170# 0.31fF
C15827 a_39222_48169# a_12257_56623# 0.40fF
C15828 ctopn a_34434_23548# 3.44fF
C15829 a_4491_47893# VDD 0.40fF
C15830 vcm_commonmode a_27314_8854# 0.31fF
C15831 vcm_commonmode a_19374_15516# 0.87fF
C15832 a_30418_56170# a_31422_56170# 0.97fF
C15833 a_30418_57174# ctopp 3.58fF
C15834 a_34251_52263# a_10515_22671# 0.40fF
C15835 ctopn a_43470_19532# 3.59fF
C15836 a_32970_31145# a_32823_29397# 0.31fF
C15837 a_18370_72234# m3_18272_72146# 2.80fF
C15838 a_3247_20495# a_5535_18012# 0.61fF
C15839 a_3987_19623# a_4839_21495# 0.37fF
C15840 a_12473_36341# a_32327_35839# 0.60fF
C15841 a_2479_50899# VDD 0.45fF
C15842 vcm_commonmode a_17366_71230# 1.82fF
C15843 a_18611_52047# a_21371_52263# 8.31fF
C15844 a_36442_61190# VDD 0.51fF
C15845 a_6559_22671# a_5085_23047# 1.85fF
C15846 vcm_commonmode a_29414_11500# 0.87fF
C15847 a_34434_58178# a_34434_57174# 1.00fF
C15848 a_12447_29199# a_5915_35943# 1.15fF
C15849 a_9529_28335# a_10873_27497# 0.39fF
C15850 vcm_commonmode a_43378_61190# 0.31fF
C15851 a_41462_16520# a_41462_15516# 1.00fF
C15852 vcm_commonmode a_33430_24552# 0.84fF
C15853 a_17599_52263# a_22386_68218# 0.38fF
C15854 a_26402_19532# a_26402_18528# 1.00fF
C15855 a_4685_37583# a_5691_36727# 0.77fF
C15856 a_7571_26151# a_10899_28879# 0.59fF
C15857 a_30326_10862# a_30418_10496# 0.32fF
C15858 a_44474_62194# ctopp 3.59fF
C15859 a_40458_70226# VDD 0.51fF
C15860 a_18351_37503# VDD 0.87fF
C15861 vcm_commonmode a_43470_55166# 0.84fF
C15862 vcm_commonmode a_35438_57174# 0.87fF
C15863 a_21382_16520# VDD 0.51fF
C15864 vcm_commonmode a_47394_70226# 0.31fF
C15865 a_36613_48169# a_37446_71230# 0.38fF
C15866 a_11115_59317# VDD 0.64fF
C15867 a_45386_60186# a_45478_60186# 0.32fF
C15868 a_3949_41935# a_5631_38127# 0.96fF
C15869 a_15851_27791# VDD 1.04fF
C15870 vcm_commonmode a_28318_16886# 0.31fF
C15871 a_21371_50959# a_26321_50095# 0.61fF
C15872 a_20378_72234# VDD 1.24fF
C15873 a_18611_52047# a_12727_58255# 0.40fF
C15874 a_42985_46831# a_48490_61190# 0.38fF
C15875 a_16955_52047# a_20378_60186# 0.38fF
C15876 a_21382_15516# a_21382_14512# 1.00fF
C15877 ctopn a_46482_20536# 3.59fF
C15878 a_4674_40277# a_5831_39189# 2.11fF
C15879 a_36717_47375# a_36442_67214# 0.38fF
C15880 a_40366_18894# a_40458_18528# 0.32fF
C15881 vcm_commonmode a_25398_72234# 0.69fF
C15882 a_2959_47113# a_3295_54421# 0.50fF
C15883 a_29414_61190# a_30418_61190# 0.97fF
C15884 a_20286_24918# a_20378_24552# 0.32fF
C15885 a_41967_31375# a_42466_20536# 0.38fF
C15886 a_1586_21959# a_2223_28617# 0.56fF
C15887 a_41597_29967# a_43269_29967# 0.36fF
C15888 vcm_commonmode a_49494_62194# 0.92fF
C15889 a_35438_68218# a_35438_67214# 1.00fF
C15890 a_17599_52263# a_22386_56170# 0.38fF
C15891 a_21187_29415# a_7295_44647# 1.13fF
C15892 vcm_commonmode a_20378_68218# 0.87fF
C15893 a_29414_58178# VDD 0.51fF
C15894 a_4792_52539# a_4831_52413# 0.73fF
C15895 a_12355_15055# a_4191_33449# 0.52fF
C15896 a_1591_21807# a_1757_21807# 0.63fF
C15897 a_17274_62194# a_17366_62194# 0.32fF
C15898 a_35615_30199# VDD 0.48fF
C15899 a_10515_63143# a_8569_24527# 0.38fF
C15900 ctopn a_46482_12504# 3.59fF
C15901 a_17507_52047# a_26465_48463# 0.52fF
C15902 a_1761_52815# a_24194_35823# 0.33fF
C15903 vcm_commonmode a_36350_58178# 0.31fF
C15904 a_13669_38517# VDD 4.69fF
C15905 a_20378_69222# a_20378_68218# 1.00fF
C15906 a_6863_49722# VDD 0.47fF
C15907 a_31768_7638# a_31422_14512# 0.38fF
C15908 a_41967_31375# a_42466_12504# 0.38fF
C15909 a_2099_59861# VDD 9.43fF
C15910 a_31330_55166# a_31422_55166# 0.32fF
C15911 a_32426_8488# a_33430_8488# 0.97fF
C15912 a_46482_67214# VDD 0.51fF
C15913 a_8491_41383# ctopn 0.32fF
C15914 a_22294_57174# a_22386_57174# 0.32fF
C15915 a_2021_17973# config_2_in[0] 0.48fF
C15916 a_25306_15882# a_25398_15516# 0.32fF
C15917 vcm_commonmode a_49494_24552# 0.87fF
C15918 ctopn a_41462_21540# 3.59fF
C15919 a_24331_44581# VDD 0.92fF
C15920 a_33430_70226# a_34434_70226# 0.97fF
C15921 a_45478_19532# a_45478_18528# 1.00fF
C15922 a_3339_43023# a_3949_41935# 0.32fF
C15923 a_12473_37429# a_16152_37601# 2.16fF
C15924 a_11067_47695# a_7000_43541# 1.96fF
C15925 a_49402_63198# VDD 0.31fF
C15926 a_30023_41959# a_12663_35431# 0.41fF
C15927 a_49402_10862# a_49494_10496# 0.32fF
C15928 vcm_commonmode a_34434_13508# 0.87fF
C15929 a_44474_59182# a_44474_58178# 1.00fF
C15930 ctopn a_18370_10496# 3.58fF
C15931 a_12901_66959# VDD 6.94fF
C15932 ctopn a_46482_17524# 3.59fF
C15933 a_6752_29941# a_6649_25615# 0.95fF
C15934 a_43470_9492# VDD 0.51fF
C15935 vcm_commonmode a_20378_56170# 0.87fF
C15936 a_17488_48731# VDD 2.84fF
C15937 vcm_commonmode a_23298_69222# 0.31fF
C15938 a_23298_71230# a_23390_71230# 0.32fF
C15939 a_31422_60186# a_31422_59182# 1.00fF
C15940 a_23390_22544# VDD 0.51fF
C15941 a_6831_63303# a_4215_51157# 0.54fF
C15942 a_41967_31375# a_42466_17524# 0.38fF
C15943 a_12355_15055# a_12981_59343# 23.65fF
C15944 a_20378_63198# a_20378_62194# 1.00fF
C15945 a_35346_11866# a_35438_11500# 0.32fF
C15946 a_49402_72234# VDD 0.74fF
C15947 a_40458_15516# a_40458_14512# 1.00fF
C15948 vcm_commonmode a_30326_22910# 0.31fF
C15949 a_18370_70226# ctopp 3.57fF
C15950 a_2004_42453# a_3023_16341# 0.49fF
C15951 a_1761_41935# VDD 10.28fF
C15952 a_39222_48169# a_10975_66407# 0.40fF
C15953 vcm_commonmode a_21290_65206# 0.31fF
C15954 a_17039_51157# VDD 5.61fF
C15955 a_2775_46025# a_2292_43291# 2.09fF
C15956 a_48490_61190# a_49494_61190# 0.97fF
C15957 a_12981_59343# a_16746_60188# 2.28fF
C15958 a_25398_9492# a_25398_8488# 1.00fF
C15959 a_5190_59575# a_11141_55535# 0.45fF
C15960 a_39362_24918# a_39454_24552# 0.32fF
C15961 a_11067_23759# a_12877_16911# 0.34fF
C15962 a_35601_27497# a_35438_23548# 0.38fF
C15963 a_1867_32839# VDD 0.37fF
C15964 VDD result_out[4] 0.82fF
C15965 a_37446_58178# a_36442_58178# 0.97fF
C15966 vcm_commonmode a_19374_61190# 0.87fF
C15967 a_20378_67214# a_21382_67214# 0.97fF
C15968 a_19374_14512# VDD 0.51fF
C15969 a_45478_64202# VDD 0.51fF
C15970 a_20267_30503# a_41842_27221# 0.33fF
C15971 a_36350_62194# a_36442_62194# 0.32fF
C15972 a_6467_55527# a_2959_47113# 3.02fF
C15973 vcm_commonmode a_26310_14878# 0.31fF
C15974 ctopn a_23390_11500# 3.59fF
C15975 a_18007_27441# a_17712_7638# 0.59fF
C15976 a_16362_70226# VDD 2.48fF
C15977 a_26753_37981# VDD 0.99fF
C15978 ctopn a_47486_18528# 3.58fF
C15979 VDD result_out[13] 0.60fF
C15980 a_76971_38925# VDD 46.80fF
C15981 a_39454_69222# a_39454_68218# 1.00fF
C15982 a_21187_29415# a_11067_46823# 0.64fF
C15983 vcm_commonmode a_23390_70226# 0.87fF
C15984 a_34251_52263# a_12901_66665# 0.40fF
C15985 a_40458_58178# vcm_commonmode 0.87fF
C15986 a_43470_58178# a_44474_58178# 0.97fF
C15987 a_1586_51335# a_1923_54591# 1.88fF
C15988 a_29414_8488# a_29414_7484# 1.00fF
C15989 a_24394_23548# VDD 0.52fF
C15990 a_21382_66210# VDD 0.51fF
C15991 a_11902_27497# a_17222_27247# 0.38fF
C15992 a_16510_8760# a_12985_7663# 1.07fF
C15993 a_12473_42869# a_26433_39631# 0.31fF
C15994 a_41370_57174# a_41462_57174# 0.32fF
C15995 a_2747_72007# VDD 1.08fF
C15996 a_12877_16911# a_16362_12504# 19.89fF
C15997 a_44382_15882# a_44474_15516# 0.32fF
C15998 a_12516_7093# a_11619_3303# 2.03fF
C15999 vcm_commonmode a_31330_23914# 0.31fF
C16000 vcm_commonmode a_28318_66210# 0.31fF
C16001 a_22386_58178# a_23390_58178# 0.97fF
C16002 a_33430_19532# VDD 0.51fF
C16003 vcm_commonmode a_16270_72234# 0.33fF
C16004 a_17366_9492# a_18370_9492# 0.97fF
C16005 a_7841_12167# a_3327_9308# 0.54fF
C16006 a_18370_13508# a_18370_12504# 1.00fF
C16007 vcm_commonmode a_40366_19898# 0.31fF
C16008 a_24394_67214# ctopp 3.59fF
C16009 a_38557_32143# a_38450_55166# 0.46fF
C16010 a_12381_43957# a_13067_38517# 0.56fF
C16011 a_23395_52047# a_27406_63198# 0.42fF
C16012 a_33430_16520# a_34434_16520# 0.97fF
C16013 a_13643_28327# a_15607_46805# 7.72fF
C16014 a_42374_71230# a_42466_71230# 0.32fF
C16015 vcm_commonmode a_41462_8488# 0.86fF
C16016 a_39454_63198# a_39454_62194# 1.00fF
C16017 a_5085_23047# a_4571_26677# 1.87fF
C16018 a_31768_55394# a_12901_58799# 0.40fF
C16019 a_24800_41953# VDD 1.66fF
C16020 a_13183_52047# a_17366_65206# 0.38fF
C16021 a_19720_7638# a_19374_8488# 0.38fF
C16022 ctopn a_36797_27497# 2.62fF
C16023 a_8583_33551# a_12641_37684# 0.38fF
C16024 a_5535_18012# a_2143_15271# 1.99fF
C16025 a_44474_9492# a_44474_8488# 1.00fF
C16026 a_41370_24918# VDD 0.36fF
C16027 a_42718_27497# a_12546_22351# 0.41fF
C16028 a_12341_3311# a_22386_23548# 0.38fF
C16029 a_39299_48783# a_38115_52263# 0.65fF
C16030 a_39223_32463# a_39454_24552# 0.46fF
C16031 a_2021_22325# a_4314_40821# 0.96fF
C16032 a_44474_58178# a_44474_57174# 1.00fF
C16033 a_39454_67214# a_40458_67214# 0.97fF
C16034 a_15607_46805# a_34062_47607# 0.49fF
C16035 a_2292_43291# a_2927_39733# 0.39fF
C16036 a_1761_25071# VDD 8.29fF
C16037 vcm_commonmode a_29414_67214# 0.87fF
C16038 a_1586_18695# a_7737_16917# 0.60fF
C16039 a_36442_20536# VDD 0.51fF
C16040 a_25398_63198# VDD 0.57fF
C16041 a_1591_26159# a_1757_26159# 0.69fF
C16042 a_26550_40871# a_24029_39355# 1.10fF
C16043 a_6515_62037# a_2840_53511# 0.48fF
C16044 a_21290_13874# a_21382_13508# 0.32fF
C16045 vcm_commonmode a_43378_20902# 0.31fF
C16046 a_13183_52047# a_17366_55166# 0.47fF
C16047 a_49494_71230# m3_49396_71142# 2.78fF
C16048 a_12725_44527# a_12621_44099# 3.50fF
C16049 vcm_commonmode a_32334_63198# 0.31fF
C16050 a_34780_56398# a_12355_15055# 0.40fF
C16051 a_26310_68218# a_26402_68218# 0.32fF
C16052 a_30005_48463# VDD 0.82fF
C16053 a_17599_52263# a_12516_7093# 0.40fF
C16054 a_19374_59182# VDD 0.51fF
C16055 a_25398_7484# a_26402_7484# 0.97fF
C16056 a_48490_8488# a_48490_7484# 1.00fF
C16057 vcm_commonmode a_26402_9492# 0.87fF
C16058 m3_21284_72146# VDD 0.39fF
C16059 a_2787_32679# a_2011_34837# 0.66fF
C16060 a_7571_29199# a_7862_34025# 0.43fF
C16061 a_36442_24552# m3_36344_24414# 2.81fF
C16062 a_43378_58178# a_43470_58178# 0.32fF
C16063 vcm_commonmode a_42466_16520# 0.87fF
C16064 a_23390_64202# ctopp 3.59fF
C16065 ctopn a_28410_13508# 3.59fF
C16066 a_31330_72234# VDD 0.61fF
C16067 vcm_commonmode a_26310_59182# 0.31fF
C16068 a_36442_12504# VDD 0.51fF
C16069 a_8273_42479# VDD 3.30fF
C16070 a_36442_9492# a_37446_9492# 0.97fF
C16071 vcm_commonmode a_43378_12870# 0.31fF
C16072 a_19374_64202# a_20378_64202# 0.97fF
C16073 a_33903_35561# VDD 0.61fF
C16074 a_37446_13508# a_37446_12504# 1.00fF
C16075 a_7803_55509# a_8453_51727# 0.55fF
C16076 a_10379_66389# a_11619_63151# 0.33fF
C16077 a_11067_46823# a_26523_28111# 0.74fF
C16078 a_10995_14333# VDD 0.44fF
C16079 a_20853_47375# VDD 0.39fF
C16080 a_10515_22671# a_15009_47919# 0.32fF
C16081 a_3325_49551# a_5135_50069# 0.53fF
C16082 a_31422_21540# VDD 0.51fF
C16083 vcm_commonmode a_34434_7484# 0.69fF
C16084 a_27752_7638# a_12877_16911# 0.41fF
C16085 a_49494_58178# VDD 1.12fF
C16086 a_5085_23047# a_5085_24759# 0.48fF
C16087 a_1591_40303# a_1757_40303# 0.69fF
C16088 vcm_commonmode a_38358_21906# 0.31fF
C16089 a_32426_69222# ctopp 3.59fF
C16090 a_4578_40455# VDD 1.55fF
C16091 vcm_commonmode a_28410_64202# 0.87fF
C16092 a_2283_15797# a_2899_16367# 0.38fF
C16093 a_12473_36341# a_1761_34319# 0.30fF
C16094 a_36442_17524# VDD 0.51fF
C16095 a_34145_49007# VDD 1.44fF
C16096 a_29760_7638# a_12877_14441# 0.41fF
C16097 a_11067_21583# a_12899_10927# 0.81fF
C16098 a_23390_60186# VDD 0.51fF
C16099 a_8491_57487# a_10680_52245# 3.16fF
C16100 a_11067_67279# a_4482_57863# 0.45fF
C16101 vcm_commonmode a_43378_17890# 0.31fF
C16102 a_30418_65206# ctopp 3.59fF
C16103 a_30565_30199# a_17712_7638# 0.41fF
C16104 a_27406_67214# a_27406_66210# 1.00fF
C16105 vcm_commonmode a_30326_60186# 0.31fF
C16106 a_10791_15529# a_10956_14459# 0.43fF
C16107 a_14646_29423# a_23626_31573# 0.44fF
C16108 a_16746_18526# a_12899_10927# 2.28fF
C16109 a_49494_15516# m3_49396_15378# 2.78fF
C16110 a_36629_27791# a_12899_11471# 0.41fF
C16111 a_7199_62839# VDD 0.60fF
C16112 a_2339_38129# a_1915_35015# 0.41fF
C16113 a_3247_20495# a_5547_31599# 0.42fF
C16114 a_10055_58791# a_19720_7638# 0.41fF
C16115 a_23390_65206# a_23390_64202# 1.00fF
C16116 a_16928_36391# VDD 1.98fF
C16117 a_40366_13874# a_40458_13508# 0.32fF
C16118 vcm_commonmode a_16746_19530# 5.36fF
C16119 a_45386_68218# a_45478_68218# 0.32fF
C16120 a_25787_28327# a_12257_56623# 0.40fF
C16121 a_2847_15039# VDD 0.37fF
C16122 vcm_commonmode a_37446_69222# 0.87fF
C16123 a_4891_47388# a_22989_48437# 2.57fF
C16124 a_44474_7484# a_45478_7484# 0.97fF
C16125 a_17366_23548# a_17366_22544# 1.00fF
C16126 a_29927_29199# a_33694_30761# 0.99fF
C16127 a_4563_32900# a_4425_32687# 0.70fF
C16128 a_2959_47113# a_8132_53511# 0.31fF
C16129 a_26310_56170# a_26402_56170# 0.32fF
C16130 a_10975_66407# a_16362_65206# 1.15fF
C16131 a_28756_55394# a_10515_22671# 0.40fF
C16132 vcm_commonmode a_44474_22544# 0.87fF
C16133 a_3339_43023# a_1761_37039# 0.57fF
C16134 a_8556_10357# VDD 0.39fF
C16135 a_28410_69222# a_29414_69222# 0.97fF
C16136 vcm_commonmode a_35438_65206# 0.87fF
C16137 a_1770_14441# a_2012_33927# 3.03fF
C16138 a_12869_2741# a_10407_47607# 0.65fF
C16139 a_37446_18528# VDD 0.51fF
C16140 a_14287_51175# a_18151_52263# 1.27fF
C16141 a_16955_52047# a_17599_52263# 0.81fF
C16142 a_20378_72234# a_21382_72234# 0.97fF
C16143 a_7479_54439# a_23763_47381# 0.62fF
C16144 a_23390_61190# a_23390_60186# 1.00fF
C16145 a_17366_24552# VDD 0.65fF
C16146 vcm_commonmode a_20286_11866# 0.31fF
C16147 ctopn a_35438_8488# 3.40fF
C16148 a_6515_67477# VDD 1.10fF
C16149 a_5831_39189# a_6883_37019# 0.71fF
C16150 a_38450_64202# a_39454_64202# 0.97fF
C16151 vcm_commonmode a_44382_18894# 0.31fF
C16152 a_37446_66210# ctopp 3.59fF
C16153 a_23395_52047# a_28881_52271# 1.24fF
C16154 a_41967_31375# a_40675_27791# 1.14fF
C16155 a_5755_14709# a_4629_13647# 0.83fF
C16156 vcm_commonmode a_24302_24918# 0.31fF
C16157 a_11067_23759# a_31659_31751# 0.35fF
C16158 a_10515_32143# a_9765_32143# 0.72fF
C16159 a_5039_42167# a_5831_39189# 0.34fF
C16160 a_2787_32679# VDD 11.54fF
C16161 a_14287_51175# a_18370_68218# 0.38fF
C16162 a_13909_38659# a_13669_37429# 4.17fF
C16163 a_28410_55166# VDD 0.60fF
C16164 a_35438_22544# a_36442_22544# 0.97fF
C16165 a_1823_53885# config_2_in[15] 0.33fF
C16166 a_2021_22325# a_6243_30662# 1.03fF
C16167 a_11067_46823# a_39727_27765# 0.68fF
C16168 a_10873_27497# VDD 3.40fF
C16169 a_19374_57174# VDD 0.51fF
C16170 vcm_commonmode a_40458_14512# 0.87fF
C16171 a_26402_65206# a_27406_65206# 0.97fF
C16172 vcm_commonmode a_19374_20536# 0.87fF
C16173 vcm_commonmode a_34342_55166# 0.31fF
C16174 a_30790_30663# a_30891_28309# 0.34fF
C16175 a_1689_10396# a_3247_20495# 0.43fF
C16176 a_3339_43023# a_1761_32143# 0.81fF
C16177 a_46482_10496# VDD 0.51fF
C16178 a_28152_40517# VDD 1.58fF
C16179 a_22386_17524# a_22386_16520# 1.00fF
C16180 vcm_commonmode a_26310_57174# 0.31fF
C16181 a_7387_46831# VDD 0.58fF
C16182 a_25787_28327# a_33430_71230# 0.38fF
C16183 a_4119_70741# a_5682_69367# 0.42fF
C16184 a_39223_32463# a_12985_16367# 0.41fF
C16185 a_25744_7638# a_12985_7663# 0.41fF
C16186 a_17366_23548# a_18370_23548# 0.97fF
C16187 a_26402_56170# a_26402_55166# 1.00fF
C16188 a_1761_52815# a_27652_38237# 0.42fF
C16189 a_46482_67214# a_46482_66210# 1.00fF
C16190 a_39299_48783# a_44474_61190# 0.38fF
C16191 a_12877_14441# a_16746_14510# 0.41fF
C16192 vcm_commonmode a_45478_23548# 0.87fF
C16193 a_14859_43447# VDD 0.60fF
C16194 vcm_commonmode a_42466_66210# 0.87fF
C16195 a_39299_48783# a_12983_63151# 0.40fF
C16196 a_28547_51175# a_32426_67214# 0.38fF
C16197 a_27752_7638# a_27406_8488# 0.38fF
C16198 vcm_commonmode a_18370_72234# 0.69fF
C16199 a_8491_27023# a_12877_16911# 0.41fF
C16200 a_33430_62194# VDD 0.51fF
C16201 a_2411_26133# a_4259_32687# 0.70fF
C16202 a_25306_61190# a_25398_61190# 0.32fF
C16203 a_19889_27497# VDD 1.02fF
C16204 a_10975_55535# VDD 0.43fF
C16205 a_10055_58791# a_40491_27247# 0.41fF
C16206 vcm_commonmode a_19374_12504# 0.87fF
C16207 ctopn a_20378_9492# 3.58fF
C16208 a_24740_7638# a_24394_23548# 0.38fF
C16209 a_5160_68315# VDD 1.25fF
C16210 a_4191_33449# a_4811_34855# 1.38fF
C16211 a_42466_65206# a_42466_64202# 1.00fF
C16212 a_31243_35831# VDD 0.64fF
C16213 ctopn a_36442_16520# 3.59fF
C16214 a_49402_8854# VDD 0.30fF
C16215 a_43267_31055# a_12981_62313# 0.40fF
C16216 vcm_commonmode a_40366_62194# 0.31fF
C16217 vcm_commonmode a_29760_7638# 10.35fF
C16218 a_14287_51175# a_18370_56170# 0.36fF
C16219 a_4811_34855# a_31964_30485# 0.52fF
C16220 a_22015_28111# a_22291_29415# 1.02fF
C16221 a_41462_15516# VDD 0.51fF
C16222 a_30764_7638# a_30418_13508# 0.38fF
C16223 a_26402_19532# a_27406_19532# 0.97fF
C16224 a_36442_23548# a_36442_22544# 1.00fF
C16225 a_7295_44647# a_35815_31751# 0.37fF
C16226 a_12263_4391# VDD 2.49fF
C16227 vcm_commonmode a_48398_15882# 0.31fF
C16228 a_41462_63198# ctopp 3.64fF
C16229 a_45386_56170# a_45478_56170# 0.32fF
C16230 a_39454_71230# VDD 0.58fF
C16231 a_30418_66210# a_30418_65206# 1.00fF
C16232 a_31422_14512# a_32426_14512# 0.97fF
C16233 a_2952_46805# a_2927_39733# 0.31fF
C16234 a_5831_39189# a_3987_19623# 1.55fF
C16235 a_1895_40516# VDD 0.85fF
C16236 a_47486_69222# a_48490_69222# 0.97fF
C16237 a_12381_35836# a_1761_35407# 0.43fF
C16238 a_30928_49007# VDD 3.48fF
C16239 vcm_commonmode a_46390_71230# 0.31fF
C16240 a_34251_52263# a_35438_72234# 0.34fF
C16241 a_12447_29199# a_28305_28879# 0.88fF
C16242 a_42466_61190# a_42466_60186# 1.00fF
C16243 a_28318_8854# a_28410_8488# 0.32fF
C16244 a_5531_22895# VDD 0.90fF
C16245 a_35438_59182# ctopp 3.59fF
C16246 vcm_commonmode a_19374_17524# 0.87fF
C16247 a_5449_25071# a_4417_22671# 0.38fF
C16248 a_18370_13508# VDD 0.52fF
C16249 a_15193_44005# VDD 1.47fF
C16250 a_42985_46831# a_12727_67753# 0.40fF
C16251 a_29322_70226# a_29414_70226# 0.32fF
C16252 a_13484_39325# a_12381_35836# 2.40fF
C16253 a_19576_51701# a_26397_51183# 1.12fF
C16254 a_6236_54421# VDD 0.55fF
C16255 a_2959_47113# a_35568_49525# 0.32fF
C16256 a_1799_29556# a_13123_38231# 0.51fF
C16257 a_28410_62194# a_28410_61190# 1.00fF
C16258 a_19374_10496# a_19374_9492# 1.00fF
C16259 vcm_commonmode a_25306_13874# 0.31fF
C16260 a_45478_65206# a_46482_65206# 0.97fF
C16261 a_12283_36919# VDD 0.61fF
C16262 a_12725_44527# a_2021_17973# 0.97fF
C16263 vcm_commonmode a_46482_63198# 0.92fF
C16264 a_41462_17524# a_41462_16520# 1.00fF
C16265 a_23395_52047# a_4351_67279# 0.70fF
C16266 a_28410_20536# a_28410_19532# 1.00fF
C16267 a_2021_22325# a_5085_23047# 0.63fF
C16268 a_7187_20719# VDD 0.57fF
C16269 m3_16264_64114# VDD 0.35fF
C16270 a_36442_23548# a_37446_23548# 0.97fF
C16271 a_12447_29199# a_4811_34855# 0.73fF
C16272 a_41261_28335# VDD 9.42fF
C16273 vcm_commonmode a_40458_59182# 0.87fF
C16274 a_33430_66210# a_34434_66210# 0.97fF
C16275 a_16510_8760# a_12899_3855# 1.81fF
C16276 a_8583_33551# a_5915_35943# 1.79fF
C16277 a_33856_42693# VDD 1.65fF
C16278 a_25787_28327# a_10975_66407# 0.40fF
C16279 a_43175_28335# a_46482_9492# 0.38fF
C16280 a_9707_51325# VDD 0.46fF
C16281 vcm_commonmode a_43362_28879# 10.09fF
C16282 a_44382_61190# a_44474_61190# 0.32fF
C16283 a_9670_24527# VDD 1.46fF
C16284 a_39454_60186# ctopp 3.59fF
C16285 a_42466_68218# VDD 0.51fF
C16286 vcm_commonmode a_20378_18528# 0.87fF
C16287 a_42374_7850# VDD 0.62fF
C16288 a_16746_67216# a_12983_63151# 0.41fF
C16289 a_10975_66407# a_2235_30503# 0.32fF
C16290 ctopn a_38450_22544# 3.58fF
C16291 a_33430_71230# a_33430_70226# 1.00fF
C16292 vcm_commonmode a_49402_68218# 0.30fF
C16293 a_45478_19532# a_46482_19532# 0.97fF
C16294 a_30991_29397# VDD 0.52fF
C16295 a_6835_46823# VDD 8.88fF
C16296 vcm_commonmode a_16746_14510# 5.36fF
C16297 a_43270_27791# a_42718_27497# 2.00fF
C16298 a_12907_56399# a_12901_58799# 0.34fF
C16299 a_49494_66210# a_49494_65206# 1.00fF
C16300 a_5993_37039# VDD 0.39fF
C16301 a_25263_41001# VDD 0.62fF
C16302 a_27535_30503# a_16863_29415# 1.57fF
C16303 a_28756_55394# a_12901_66665# 0.40fF
C16304 a_29414_20536# a_30418_20536# 0.97fF
C16305 a_47394_8854# a_47486_8488# 0.32fF
C16306 a_11522_23145# VDD 0.44fF
C16307 vcm_commonmode a_29414_10496# 0.87fF
C16308 a_18370_63198# a_19374_63198# 0.97fF
C16309 a_23119_31599# VDD 1.24fF
C16310 ctopn a_34434_14512# 3.59fF
C16311 a_2686_70223# VDD 4.27fF
C16312 vcm_commonmode a_44474_60186# 0.87fF
C16313 a_17366_71230# ctopp 3.24fF
C16314 a_11067_23759# a_34759_31029# 0.58fF
C16315 a_14354_32117# a_14361_29967# 0.30fF
C16316 a_21233_44220# VDD 0.86fF
C16317 a_48398_70226# a_48490_70226# 0.32fF
C16318 a_18278_58178# a_18370_58178# 0.32fF
C16319 a_13123_38231# a_19096_36513# 2.75fF
C16320 a_5612_52520# VDD 0.67fF
C16321 a_11299_62215# VDD 0.37fF
C16322 a_47486_62194# a_47486_61190# 1.00fF
C16323 a_38450_10496# a_38450_9492# 1.00fF
C16324 a_42466_56170# VDD 0.52fF
C16325 a_13097_39631# a_13669_39605# 0.42fF
C16326 a_4191_33449# a_5079_35639# 0.68fF
C16327 a_34780_56398# a_34434_55166# 0.43fF
C16328 a_1761_44111# a_1803_19087# 0.50fF
C16329 a_25398_8488# VDD 0.58fF
C16330 vcm_commonmode a_16746_62196# 5.36fF
C16331 a_18611_52047# a_23390_63198# 0.42fF
C16332 a_29322_16886# a_29414_16520# 0.32fF
C16333 vcm_commonmode a_49402_56170# 0.30fF
C16334 ctopn a_39454_23548# 3.40fF
C16335 a_6559_22671# VDD 8.08fF
C16336 a_47486_20536# a_47486_19532# 1.00fF
C16337 a_9135_27239# a_21382_13508# 0.38fF
C16338 a_2411_26133# a_2317_28892# 0.90fF
C16339 vcm_commonmode a_32334_8854# 0.31fF
C16340 m3_16264_11362# VDD 0.34fF
C16341 a_1952_60431# a_2952_53333# 1.28fF
C16342 a_18979_30287# a_3339_30503# 0.55fF
C16343 vcm_commonmode a_24394_15516# 0.87fF
C16344 a_35438_57174# ctopp 3.58fF
C16345 a_16746_71232# VDD 33.49fF
C16346 a_18151_52263# a_12901_58799# 0.40fF
C16347 a_8583_33551# inp_analog 1.83fF
C16348 ctopn a_48490_19532# 3.43fF
C16349 a_21382_72234# m3_21284_72146# 2.80fF
C16350 a_14293_41807# VDD 2.47fF
C16351 a_5963_36585# a_1761_32143# 0.58fF
C16352 vcm_commonmode a_22386_71230# 0.86fF
C16353 a_26310_72234# a_26402_72234# 0.32fF
C16354 a_27406_21540# a_27406_20536# 1.00fF
C16355 a_41462_61190# VDD 0.51fF
C16356 VDD config_2_in[12] 0.84fF
C16357 vcm_commonmode a_34434_11500# 0.87fF
C16358 a_33864_28111# a_34434_22544# 0.38fF
C16359 a_11619_63151# VDD 0.84fF
C16360 a_29414_12504# a_30418_12504# 0.97fF
C16361 a_35346_67214# a_35438_67214# 0.32fF
C16362 vcm_commonmode a_48398_61190# 0.31fF
C16363 a_12727_15529# a_12877_14441# 23.87fF
C16364 vcm_commonmode a_38450_24552# 0.84fF
C16365 a_2473_34293# a_1586_21959# 0.73fF
C16366 vcm_commonmode a_20286_67214# 0.31fF
C16367 a_1586_51335# a_4215_51157# 0.62fF
C16368 a_9135_27239# a_12899_10927# 0.41fF
C16369 a_15439_49525# VDD 5.55fF
C16370 a_7295_44647# a_33641_29967# 1.16fF
C16371 a_43495_28487# VDD 0.63fF
C16372 a_11067_23759# a_12895_13967# 0.36fF
C16373 a_45478_70226# VDD 0.51fF
C16374 a_16362_13508# a_16746_13506# 2.28fF
C16375 a_20378_68218# ctopp 3.59fF
C16376 vcm_commonmode a_49494_55166# 0.87fF
C16377 a_7948_38377# VDD 0.90fF
C16378 a_23395_52047# a_12355_15055# 0.40fF
C16379 a_30764_7638# a_30418_7484# 0.34fF
C16380 vcm_commonmode a_40458_57174# 0.87fF
C16381 a_5915_30287# a_8117_30287# 0.67fF
C16382 a_17039_51157# a_21095_47919# 0.37fF
C16383 a_26402_16520# VDD 0.51fF
C16384 a_48490_20536# a_49494_20536# 0.97fF
C16385 a_21290_7850# a_21382_7484# 0.32fF
C16386 vcm_commonmode a_17274_9858# 0.33fF
C16387 a_10975_66407# a_13809_48463# 0.49fF
C16388 a_29414_24552# m3_29316_24414# 2.81fF
C16389 a_37446_63198# a_38450_63198# 0.97fF
C16390 vcm_commonmode a_33338_16886# 0.31fF
C16391 a_8531_70543# a_29361_51727# 0.37fF
C16392 a_24302_72234# VDD 0.62fF
C16393 vcm_commonmode a_16362_59182# 4.47fF
C16394 a_41289_43421# VDD 1.08fF
C16395 a_28756_7638# a_28410_9492# 0.38fF
C16396 ctopn a_26748_7638# 2.62fF
C16397 a_30757_37455# a_12473_36341# 0.49fF
C16398 a_24394_21540# a_25398_21540# 0.97fF
C16399 a_32334_9858# a_32426_9492# 0.32fF
C16400 a_10472_26159# a_11574_22869# 0.51fF
C16401 a_21663_35327# VDD 0.97fF
C16402 a_8583_33551# a_31659_31751# 0.31fF
C16403 a_18370_7484# VDD 1.42fF
C16404 a_48398_16886# a_48490_16520# 0.32fF
C16405 vcm_commonmode a_25398_68218# 0.87fF
C16406 a_34434_58178# VDD 0.51fF
C16407 a_31422_59182# a_32426_59182# 0.97fF
C16408 a_41597_29967# VDD 1.91fF
C16409 a_7461_27247# a_8491_27023# 0.57fF
C16410 a_20378_56170# ctopp 3.40fF
C16411 a_1929_12131# a_7999_13083# 0.32fF
C16412 vcm_commonmode a_19282_64202# 0.31fF
C16413 a_29414_17524# a_30418_17524# 0.97fF
C16414 a_46482_21540# a_46482_20536# 1.00fF
C16415 a_33430_24552# a_33430_23548# 1.00fF
C16416 a_2021_17973# a_2012_33927# 1.83fF
C16417 a_48490_12504# a_49494_12504# 0.97fF
C16418 a_18370_12504# a_18370_11500# 1.00fF
C16419 a_33694_30761# VDD 3.24fF
C16420 a_3978_74183# VDD 0.66fF
C16421 ctopn a_46482_21540# 3.59fF
C16422 a_32887_44581# VDD 0.87fF
C16423 a_13183_52047# a_12983_63151# 0.40fF
C16424 a_11067_63143# a_7000_43541# 0.39fF
C16425 a_1952_60431# a_3295_54421# 0.76fF
C16426 vcm_commonmode a_39454_13508# 0.87fF
C16427 a_19374_61190# ctopp 3.59fF
C16428 ctopn a_23390_10496# 3.59fF
C16429 a_41967_31375# a_42466_21540# 0.38fF
C16430 a_21382_69222# VDD 0.51fF
C16431 a_48490_9492# VDD 0.54fF
C16432 a_21371_52263# a_12257_56623# 0.40fF
C16433 vcm_commonmode a_25398_56170# 0.87fF
C16434 a_19807_28111# a_28108_48463# 0.34fF
C16435 vcm_commonmode a_28318_69222# 0.31fF
C16436 a_35601_27497# a_35438_14512# 0.38fF
C16437 a_40366_7850# a_40458_7484# 0.32fF
C16438 a_28410_22544# VDD 0.51fF
C16439 a_19374_65206# VDD 0.51fF
C16440 a_40691_30511# VDD 0.44fF
C16441 vcm_commonmode a_12727_15529# 6.31fF
C16442 a_15681_27497# a_11430_26159# 0.34fF
C16443 a_8935_27791# a_7369_24233# 0.45fF
C16444 a_17507_52047# a_10515_22671# 0.40fF
C16445 vcm_commonmode a_35346_22910# 0.31fF
C16446 a_23390_70226# ctopp 3.58fF
C16447 a_36507_31573# a_34759_31029# 0.49fF
C16448 a_40458_58178# ctopp 3.59fF
C16449 a_24302_69222# a_24394_69222# 0.32fF
C16450 vcm_commonmode a_26310_65206# 0.31fF
C16451 a_30418_18528# a_30418_17524# 1.00fF
C16452 a_43470_21540# a_44474_21540# 0.97fF
C16453 a_42718_27497# a_12985_16367# 0.41fF
C16454 a_1761_27791# a_12549_35836# 0.31fF
C16455 a_12447_29199# a_13239_29575# 0.49fF
C16456 a_2411_26133# a_1683_31599# 0.34fF
C16457 a_34342_64202# a_34434_64202# 0.32fF
C16458 a_21479_34239# VDD 0.77fF
C16459 ctopn a_18370_15516# 3.58fF
C16460 vcm_commonmode a_24394_61190# 0.87fF
C16461 a_1761_50639# a_1761_44111# 1.10fF
C16462 a_24394_14512# VDD 0.51fF
C16463 a_49494_16520# m3_49396_16382# 2.78fF
C16464 a_19282_55166# VDD 0.35fF
C16465 a_31330_22910# a_31422_22544# 0.32fF
C16466 a_20378_10496# a_21382_10496# 0.97fF
C16467 vcm_commonmode a_31330_14878# 0.31fF
C16468 ctopn a_28410_11500# 3.59fF
C16469 a_22294_65206# a_22386_65206# 0.32fF
C16470 a_31422_14512# a_31422_13508# 1.00fF
C16471 a_33727_38007# VDD 0.65fF
C16472 a_3143_66972# a_7213_62215# 0.52fF
C16473 a_9135_27239# a_21382_7484# 0.34fF
C16474 a_48490_17524# a_49494_17524# 0.97fF
C16475 vcm_commonmode a_16362_57174# 4.47fF
C16476 ctopn a_32426_24552# 1.02fF
C16477 a_29760_55394# a_29414_71230# 0.38fF
C16478 vcm_commonmode a_28410_70226# 0.87fF
C16479 a_35438_60186# a_36442_60186# 0.97fF
C16480 a_29414_23548# VDD 0.52fF
C16481 a_27752_7638# a_12895_13967# 0.41fF
C16482 a_26402_66210# VDD 0.51fF
C16483 a_9219_11471# a_9455_11079# 0.37fF
C16484 a_37446_12504# a_37446_11500# 1.00fF
C16485 a_39222_48169# a_40458_61190# 0.38fF
C16486 vcm_commonmode a_36350_23914# 0.31fF
C16487 a_2235_30503# a_8739_28879# 0.40fF
C16488 a_28756_55394# a_28410_67214# 0.38fF
C16489 a_24394_70226# a_24394_69222# 1.00fF
C16490 vcm_commonmode a_33338_66210# 0.31fF
C16491 a_36613_48169# a_12983_63151# 0.40fF
C16492 a_30418_18528# a_31422_18528# 0.97fF
C16493 a_38450_19532# VDD 0.51fF
C16494 a_29760_7638# a_12899_11471# 0.41fF
C16495 a_8273_42479# a_9307_30663# 0.38fF
C16496 a_20267_30503# a_28670_30663# 0.33fF
C16497 a_4571_26677# VDD 4.40fF
C16498 a_31768_7638# a_11067_21583# 0.41fF
C16499 vcm_commonmode a_45386_19898# 0.31fF
C16500 a_29414_67214# ctopp 3.59fF
C16501 a_1761_46287# a_6473_40277# 0.62fF
C16502 a_39389_52271# a_12981_62313# 0.40fF
C16503 a_7000_43541# a_15607_46805# 0.63fF
C16504 a_35539_47919# VDD 0.55fF
C16505 a_22294_19898# a_22386_19532# 0.32fF
C16506 a_12341_3311# a_22386_14512# 0.38fF
C16507 a_10791_57711# VDD 0.42fF
C16508 vcm_commonmode a_46482_8488# 0.86fF
C16509 a_23390_11500# a_23390_10496# 1.00fF
C16510 a_6782_29967# VDD 0.32fF
C16511 vcm_commonmode a_17366_58178# 1.83fF
C16512 a_30912_39429# VDD 1.67fF
C16513 a_27314_14878# a_27406_14512# 0.32fF
C16514 a_8753_31055# a_6459_30511# 0.30fF
C16515 a_3339_43023# a_4495_35925# 0.32fF
C16516 a_32795_41855# VDD 0.87fF
C16517 a_43378_69222# a_43470_69222# 0.32fF
C16518 a_49494_18528# a_49494_17524# 1.00fF
C16519 a_19720_7638# a_12877_14441# 0.41fF
C16520 a_7571_29199# a_7369_24233# 0.62fF
C16521 a_21382_55166# a_22386_55166# 0.97fF
C16522 a_46390_24918# VDD 0.36fF
C16523 a_30764_7638# a_11067_21583# 0.41fF
C16524 a_7155_55509# a_6095_44807# 0.39fF
C16525 a_11067_63143# a_5915_35943# 0.71fF
C16526 vcm_commonmode a_34434_67214# 0.87fF
C16527 a_41427_52263# a_12727_67753# 0.40fF
C16528 a_2099_59861# a_3247_20495# 0.34fF
C16529 ctopn a_43269_29967# 2.61fF
C16530 a_41462_20536# VDD 0.51fF
C16531 a_32951_27247# a_12899_10927# 0.41fF
C16532 a_30418_63198# VDD 0.57fF
C16533 a_1761_40847# a_1761_30511# 2.25fF
C16534 a_39454_10496# a_40458_10496# 0.97fF
C16535 a_10055_58791# a_32772_7638# 0.41fF
C16536 a_41370_65206# a_41462_65206# 0.32fF
C16537 vcm_commonmode a_48398_20902# 0.31fF
C16538 a_30052_32117# a_28756_7638# 0.44fF
C16539 vcm_commonmode a_37354_63198# 0.31fF
C16540 a_10239_16367# a_10405_16367# 0.69fF
C16541 a_45478_72234# a_45478_71230# 1.00fF
C16542 a_24394_59182# VDD 0.51fF
C16543 a_5963_20149# VDD 0.95fF
C16544 vcm_commonmode a_31422_9492# 0.87fF
C16545 a_32334_23914# a_32426_23548# 0.32fF
C16546 a_6519_65301# VDD 0.38fF
C16547 a_25398_11500# a_26402_11500# 0.97fF
C16548 vcm_commonmode a_47486_16520# 0.87fF
C16549 a_11067_13095# a_6451_22895# 0.37fF
C16550 a_28410_64202# ctopp 3.59fF
C16551 ctopn a_33430_13508# 3.59fF
C16552 a_49494_67214# m3_49396_67126# 2.78fF
C16553 a_8273_42479# a_5363_30503# 1.92fF
C16554 a_34251_52263# VDD 15.19fF
C16555 a_1761_52815# a_25133_37571# 0.45fF
C16556 a_29322_66210# a_29414_66210# 0.32fF
C16557 vcm_commonmode a_31330_59182# 0.31fF
C16558 a_4811_34855# a_27752_7638# 0.48fF
C16559 vcm_commonmode m3_16264_68130# 3.21fF
C16560 a_3339_43023# a_13123_38231# 0.83fF
C16561 a_2292_43291# a_6559_42479# 0.70fF
C16562 a_41462_12504# VDD 0.51fF
C16563 a_43470_70226# a_43470_69222# 1.00fF
C16564 a_21371_52263# a_10975_66407# 0.44fF
C16565 vcm_commonmode a_39222_48169# 10.02fF
C16566 a_40675_27791# a_12727_13353# 0.41fF
C16567 a_5085_24759# VDD 1.94fF
C16568 vcm_commonmode a_48398_12870# 0.31fF
C16569 a_49494_63198# m3_49396_63110# 2.78fF
C16570 a_29414_24552# a_30418_24552# 0.97fF
C16571 a_11416_12283# a_11455_12157# 0.57fF
C16572 a_12516_7093# a_12355_15055# 0.53fF
C16573 a_9989_46831# a_7571_26151# 0.76fF
C16574 a_41872_29423# a_12901_66959# 0.40fF
C16575 a_41370_19898# a_41462_19532# 0.32fF
C16576 a_36442_21540# VDD 0.51fF
C16577 vcm_commonmode a_39454_7484# 0.69fF
C16578 a_42709_29199# a_48490_18528# 0.38fF
C16579 a_43175_28335# a_12899_10927# 0.41fF
C16580 a_8491_27023# a_12895_13967# 0.41fF
C16581 a_26402_62194# a_27406_62194# 0.97fF
C16582 a_42466_11500# a_42466_10496# 1.00fF
C16583 a_19442_28585# VDD 0.60fF
C16584 a_1761_50639# a_25133_37571# 2.65fF
C16585 a_46390_14878# a_46482_14512# 0.32fF
C16586 a_34639_38825# VDD 0.59fF
C16587 vcm_commonmode a_43378_21906# 0.31fF
C16588 a_37446_69222# ctopp 3.59fF
C16589 a_1591_45205# a_1757_45205# 0.42fF
C16590 vcm_commonmode a_33430_64202# 0.87fF
C16591 a_29760_7638# a_29414_8488# 0.38fF
C16592 a_41462_17524# VDD 0.51fF
C16593 a_45478_72234# a_46482_72234# 0.97fF
C16594 a_17507_52047# a_12901_66665# 0.40fF
C16595 a_40491_27247# a_12877_14441# 0.41fF
C16596 a_25306_20902# a_25398_20536# 0.32fF
C16597 a_28410_60186# VDD 0.51fF
C16598 a_39454_55166# a_40458_55166# 0.97fF
C16599 vcm_commonmode a_20286_10862# 0.31fF
C16600 a_36629_27791# a_12985_7663# 0.41fF
C16601 vcm_commonmode a_48398_17890# 0.31fF
C16602 a_35438_65206# ctopp 3.59fF
C16603 a_31422_57174# a_32426_57174# 0.97fF
C16604 vcm_commonmode a_35346_60186# 0.31fF
C16605 a_1591_66415# a_1757_66415# 0.39fF
C16606 a_34434_15516# a_35438_15516# 0.97fF
C16607 a_30764_7638# a_30418_11500# 0.38fF
C16608 a_10055_58791# a_37919_28111# 0.41fF
C16609 a_40675_27791# a_10515_23975# 0.41fF
C16610 vcm_commonmode a_21382_19532# 0.87fF
C16611 a_12579_44310# a_12381_43957# 0.30fF
C16612 a_19720_55394# a_19374_63198# 0.42fF
C16613 a_1591_64239# a_3295_62083# 0.42fF
C16614 vcm_commonmode a_19720_7638# 10.36fF
C16615 a_22015_28111# a_12907_27023# 0.79fF
C16616 a_27869_50095# a_31753_47919# 0.32fF
C16617 a_11067_46823# a_4443_46607# 1.49fF
C16618 vcm_commonmode a_42466_69222# 0.87fF
C16619 a_32426_71230# a_33430_71230# 0.97fF
C16620 a_6559_59663# a_26218_48981# 0.54fF
C16621 a_8491_57487# VDD 6.13fF
C16622 a_43269_29967# a_47486_18528# 0.38fF
C16623 a_32772_7638# a_32426_19532# 0.38fF
C16624 a_44474_11500# a_45478_11500# 0.97fF
C16625 a_4351_67279# a_16385_51183# 0.50fF
C16626 a_48398_66210# a_48490_66210# 0.32fF
C16627 vcm_commonmode a_49494_22544# 0.89fF
C16628 vcm_commonmode m3_16264_15378# 3.21fF
C16629 a_18370_11500# VDD 0.52fF
C16630 a_41351_42405# VDD 0.90fF
C16631 vcm_commonmode a_40458_65206# 0.87fF
C16632 a_43362_28879# a_12355_65103# 0.40fF
C16633 a_42466_18528# VDD 0.51fF
C16634 vcm_commonmode a_12947_71576# 4.77fF
C16635 a_22386_24552# VDD 0.60fF
C16636 vcm_commonmode a_25306_11866# 0.31fF
C16637 ctopn a_40458_8488# 3.40fF
C16638 a_12355_15055# a_11067_63143# 0.86fF
C16639 a_25306_12870# a_25398_12504# 0.32fF
C16640 vcm_commonmode a_49402_18894# 0.31fF
C16641 a_42466_66210# ctopp 3.59fF
C16642 a_2927_68565# a_1768_13103# 0.72fF
C16643 a_11067_67279# a_23736_7638# 0.41fF
C16644 vcm_commonmode a_29322_24918# 0.31fF
C16645 a_12907_27023# a_37557_32463# 2.58fF
C16646 a_2539_42106# VDD 0.94fF
C16647 a_20378_59182# a_20378_58178# 1.00fF
C16648 a_12869_2741# VDD 16.90fF
C16649 a_43270_27791# a_12899_10927# 0.41fF
C16650 a_45478_62194# a_46482_62194# 0.97fF
C16651 a_24394_57174# VDD 0.51fF
C16652 vcm_commonmode a_45478_14512# 0.87fF
C16653 a_9731_22895# a_11130_22869# 0.38fF
C16654 a_1761_50639# a_12473_36341# 0.37fF
C16655 a_13669_37429# VDD 6.11fF
C16656 vcm_commonmode a_24394_20536# 0.87fF
C16657 vcm_commonmode a_39362_55166# 0.30fF
C16658 a_24029_39355# VDD 1.81fF
C16659 a_16955_52047# a_12355_15055# 0.40fF
C16660 vcm_commonmode a_31330_57174# 0.31fF
C16661 a_24740_7638# a_24394_14512# 0.38fF
C16662 a_44382_20902# a_44474_20536# 0.32fF
C16663 a_10515_22671# a_10073_23439# 0.50fF
C16664 a_11067_13095# a_6646_50639# 0.39fF
C16665 VDD config_1_in[3] 1.23fF
C16666 a_22386_24552# m3_22288_24414# 2.81fF
C16667 a_33338_63198# a_33430_63198# 0.32fF
C16668 a_1761_41935# a_15189_39889# 1.32fF
C16669 a_24394_57174# a_24394_56170# 1.00fF
C16670 a_11067_13095# a_6243_30662# 0.32fF
C16671 a_4674_40277# a_8080_47607# 0.30fF
C16672 a_25447_43447# VDD 0.63fF
C16673 vcm_commonmode a_47486_66210# 0.87fF
C16674 a_20286_21906# a_20378_21540# 0.32fF
C16675 a_2411_19605# a_10883_18543# 0.70fF
C16676 a_38450_62194# VDD 0.51fF
C16677 a_18979_30287# a_20505_29967# 1.54fF
C16678 vcm_commonmode a_24394_12504# 0.87fF
C16679 ctopn a_25398_9492# 3.58fF
C16680 a_7155_55509# VDD 3.60fF
C16681 ctopn a_41462_16520# 3.59fF
C16682 a_16510_8760# a_12947_23413# 1.04fF
C16683 vcm_commonmode a_45386_62194# 0.31fF
C16684 a_7580_61751# a_7803_55509# 1.15fF
C16685 vcm_commonmode a_40491_27247# 10.40fF
C16686 a_46482_15516# VDD 0.51fF
C16687 a_1941_47381# VDD 0.30fF
C16688 vcm_commonmode a_16746_68220# 5.36fF
C16689 a_1586_18695# a_2411_18517# 1.25fF
C16690 a_27314_59182# a_27406_59182# 0.32fF
C16691 a_13837_38772# a_13909_38659# 0.78fF
C16692 a_12659_54965# a_6775_53877# 0.33fF
C16693 a_11067_13095# a_4298_58951# 0.35fF
C16694 a_46482_63198# ctopp 3.64fF
C16695 a_7847_40847# a_8017_40847# 0.42fF
C16696 a_44474_71230# VDD 0.58fF
C16697 a_12985_16367# a_16362_11500# 1.27fF
C16698 a_75111_39506# VDD 0.45fF
C16699 vcm_commonmode a_19374_21540# 0.87fF
C16700 a_16228_28335# a_17651_30485# 0.43fF
C16701 a_4706_40847# VDD 0.40fF
C16702 a_25306_17890# a_25398_17524# 0.32fF
C16703 a_40458_59182# ctopp 3.59fF
C16704 a_31422_64202# a_31422_63198# 1.23fF
C16705 a_44382_12870# a_44474_12504# 0.32fF
C16706 vcm_commonmode a_24394_17524# 0.87fF
C16707 a_5475_74895# VDD 0.40fF
C16708 a_28547_51175# a_2775_46025# 0.91fF
C16709 a_43362_28879# ctopp 2.61fF
C16710 a_23390_13508# VDD 0.51fF
C16711 a_2021_22325# VDD 7.81fF
C16712 a_9135_27239# a_21382_11500# 0.38fF
C16713 a_23390_22544# a_23390_21540# 1.00fF
C16714 vcm_commonmode a_30326_13874# 0.31fF
C16715 a_25971_52263# a_20267_30503# 0.38fF
C16716 a_30418_13508# a_31422_13508# 0.97fF
C16717 a_24515_36965# VDD 1.03fF
C16718 m2_48260_54946# m3_48392_55078# 0.85fF
C16719 a_35438_68218# a_36442_68218# 0.97fF
C16720 a_12546_22351# a_16362_10496# 1.27fF
C16721 a_19720_55394# a_12257_56623# 0.40fF
C16722 a_16510_8760# a_3339_30503# 0.36fF
C16723 a_2419_48783# a_1761_50639# 0.81fF
C16724 a_1768_16367# a_1761_27791# 0.31fF
C16725 a_4075_64239# VDD 0.59fF
C16726 a_47486_56170# a_47486_55166# 1.00fF
C16727 a_6459_30511# VDD 2.78fF
C16728 a_43470_57174# a_43470_56170# 1.00fF
C16729 vcm_commonmode a_45478_59182# 0.87fF
C16730 ctopn a_12985_19087# 2.95fF
C16731 vcm_commonmode a_16362_65206# 4.47fF
C16732 a_14983_51157# VDD 1.23fF
C16733 a_6559_59663# a_19478_51959# 0.40fF
C16734 a_39362_21906# a_39454_21540# 0.32fF
C16735 a_6382_61127# VDD 0.48fF
C16736 a_11067_63143# a_11887_19087# 0.86fF
C16737 a_44474_60186# ctopp 3.59fF
C16738 a_20378_58178# a_20378_57174# 1.00fF
C16739 ctopn a_16746_8486# 1.36fF
C16740 a_16510_8760# a_12727_13353# 1.08fF
C16741 a_47486_68218# VDD 0.51fF
C16742 vcm_commonmode a_25398_18528# 0.87fF
C16743 a_47394_7850# VDD 0.62fF
C16744 a_27406_16520# a_27406_15516# 1.00fF
C16745 ctopn a_43470_22544# 3.58fF
C16746 a_2012_33927# a_2347_28918# 0.31fF
C16747 a_7939_30503# a_8117_30287# 0.34fF
C16748 a_5993_32687# a_7281_29423# 0.62fF
C16749 a_12907_27023# a_22291_29415# 0.90fF
C16750 a_2656_45895# VDD 1.67fF
C16751 a_4482_57863# a_21003_49007# 0.63fF
C16752 a_46390_59182# a_46482_59182# 0.32fF
C16753 a_12869_2741# a_29055_49525# 0.33fF
C16754 a_6372_38279# a_5691_36727# 0.57fF
C16755 a_2124_56891# VDD 0.62fF
C16756 a_16746_62196# ctopp 1.68fF
C16757 a_11955_69653# VDD 0.35fF
C16758 a_33819_41001# VDD 0.65fF
C16759 a_12516_7093# a_11067_66191# 1.39fF
C16760 a_44382_17890# a_44474_17524# 0.32fF
C16761 a_17095_49525# VDD 0.55fF
C16762 a_21371_50959# a_25398_71230# 0.38fF
C16763 vcm_commonmode a_19282_70226# 0.31fF
C16764 a_31330_60186# a_31422_60186# 0.32fF
C16765 vcm_commonmode a_34434_10496# 0.87fF
C16766 ctopn a_39454_14512# 3.59fF
C16767 a_2223_28617# a_2315_24540# 1.22fF
C16768 a_2317_28892# a_3301_27791# 0.43fF
C16769 a_6607_42167# a_6579_42255# 0.38fF
C16770 a_1823_66941# a_1768_13103# 0.54fF
C16771 vcm_commonmode a_49494_60186# 0.91fF
C16772 a_36717_47375# a_36442_61190# 0.38fF
C16773 a_22386_71230# ctopp 3.40fF
C16774 ctopn a_18370_20536# 3.58fF
C16775 a_1761_49007# a_12725_44527# 2.25fF
C16776 a_1757_12565# VDD 0.64fF
C16777 a_30323_44265# VDD 0.64fF
C16778 a_25971_52263# a_12983_63151# 0.40fF
C16779 a_18151_52263# a_24394_67214# 0.38fF
C16780 a_26310_18894# a_26402_18528# 0.32fF
C16781 a_17039_51157# a_24683_51183# 0.35fF
C16782 a_1849_52271# VDD 0.62fF
C16783 a_6224_73095# a_7707_70741# 1.53fF
C16784 a_12341_3311# a_12899_10927# 1.38fF
C16785 a_42466_22544# a_42466_21540# 1.00fF
C16786 a_3983_20719# a_4149_20719# 0.39fF
C16787 a_47486_56170# VDD 0.52fF
C16788 a_42718_27497# a_44474_24552# 0.54fF
C16789 a_31768_7638# a_12546_22351# 0.41fF
C16790 a_16510_8760# a_10515_23975# 1.11fF
C16791 a_30418_8488# VDD 0.58fF
C16792 a_21382_68218# a_21382_67214# 1.00fF
C16793 vcm_commonmode a_21382_62194# 0.87fF
C16794 a_28547_51175# a_12981_62313# 0.40fF
C16795 ctopn a_44474_23548# 3.40fF
C16796 a_2292_43291# a_5179_47919# 0.31fF
C16797 a_15009_47919# VDD 0.35fF
C16798 vcm_commonmode a_37354_8854# 0.31fF
C16799 vcm_commonmode a_29414_15516# 0.87fF
C16800 ctopn a_18370_12504# 3.58fF
C16801 a_35438_56170# a_36442_56170# 0.97fF
C16802 a_40458_57174# ctopp 3.58fF
C16803 a_12191_39095# VDD 0.59fF
C16804 a_19626_31751# a_26523_29199# 0.32fF
C16805 a_24394_72234# m3_24296_72146# 2.80fF
C16806 a_2216_28309# a_3607_34639# 0.57fF
C16807 a_30928_49007# a_22843_29415# 0.50fF
C16808 vcm_commonmode a_27406_71230# 0.86fF
C16809 a_28756_55394# a_28410_72234# 0.35fF
C16810 a_46482_61190# VDD 0.51fF
C16811 a_18370_8488# a_19374_8488# 0.97fF
C16812 vcm_commonmode a_39454_11500# 0.87fF
C16813 a_16362_59182# ctopp 1.35fF
C16814 a_30764_7638# a_12546_22351# 0.41fF
C16815 a_18370_67214# VDD 0.52fF
C16816 a_8531_70543# a_6831_63303# 3.62fF
C16817 a_46482_16520# a_46482_15516# 1.00fF
C16818 a_11067_67279# a_11155_30663# 0.38fF
C16819 vcm_commonmode a_43470_24552# 0.84fF
C16820 a_6361_44655# VDD 0.74fF
C16821 vcm_commonmode a_25306_67214# 0.31fF
C16822 a_34780_56398# a_12727_67753# 0.40fF
C16823 a_19374_70226# a_20378_70226# 0.97fF
C16824 a_31422_19532# a_31422_18528# 1.00fF
C16825 a_1923_54591# a_4831_58497# 0.32fF
C16826 a_35346_10862# a_35438_10496# 0.32fF
C16827 a_14912_27497# VDD 0.74fF
C16828 a_10515_63143# a_8105_21263# 0.34fF
C16829 a_3663_39991# a_3759_39991# 0.31fF
C16830 a_25787_28327# a_33430_58178# 0.38fF
C16831 a_32365_37692# VDD 0.85fF
C16832 a_25398_68218# ctopp 3.59fF
C16833 ctopn a_18370_17524# 3.58fF
C16834 a_14293_39631# VDD 1.03fF
C16835 vcm_commonmode a_45478_57174# 0.87fF
C16836 a_11067_46823# a_16863_29415# 1.66fF
C16837 a_26662_48981# a_26218_48981# 0.73fF
C16838 a_31422_16520# VDD 0.51fF
C16839 a_28108_48463# VDD 1.00fF
C16840 a_41462_72234# a_41462_71230# 1.00fF
C16841 a_17366_60186# a_17366_59182# 1.00fF
C16842 vcm_commonmode a_22294_9858# 0.31fF
C16843 a_1770_14441# a_1923_54591# 1.19fF
C16844 a_21290_11866# a_21382_11500# 0.32fF
C16845 vcm_commonmode a_38358_16886# 0.31fF
C16846 a_11902_27497# a_12707_26159# 0.55fF
C16847 a_15459_41781# a_16012_41959# 0.31fF
C16848 a_28756_55394# VDD 6.81fF
C16849 a_26402_15516# a_26402_14512# 1.00fF
C16850 a_7862_34025# a_8485_29673# 1.02fF
C16851 a_19720_55394# a_10975_66407# 0.40fF
C16852 a_45386_18894# a_45478_18528# 0.32fF
C16853 vcm_commonmode a_25787_28327# 10.04fF
C16854 a_18979_30287# a_33839_28309# 0.30fF
C16855 a_34434_61190# a_35438_61190# 0.97fF
C16856 a_25306_24918# a_25398_24552# 0.32fF
C16857 a_13005_43983# a_13835_43177# 0.63fF
C16858 a_23390_7484# VDD 1.23fF
C16859 a_40458_68218# a_40458_67214# 1.00fF
C16860 a_1823_66941# a_1770_14441# 0.59fF
C16861 a_2606_41079# a_4563_32900# 0.40fF
C16862 vcm_commonmode a_30418_68218# 0.87fF
C16863 a_36717_47375# a_12901_66959# 0.40fF
C16864 a_15285_52245# a_15557_52245# 0.49fF
C16865 a_36797_27497# a_12985_19087# 0.41fF
C16866 a_17366_64202# VDD 0.58fF
C16867 a_22294_62194# a_22386_62194# 0.32fF
C16868 a_5087_29423# VDD 0.80fF
C16869 m2_48260_24282# VDD 0.39fF
C16870 a_25398_56170# ctopp 3.40fF
C16871 a_17033_38565# VDD 1.24fF
C16872 a_11067_67279# a_39673_28111# 0.41fF
C16873 ctopn a_19374_18528# 3.59fF
C16874 a_36579_41271# VDD 0.64fF
C16875 a_25398_69222# a_25398_68218# 1.00fF
C16876 vcm_commonmode a_24302_64202# 0.31fF
C16877 a_12381_35836# a_13669_35253# 0.79fF
C16878 a_28639_49551# VDD 0.34fF
C16879 a_41261_28335# a_41872_29423# 1.21fF
C16880 a_35346_55166# a_35438_55166# 0.32fF
C16881 a_37446_8488# a_38450_8488# 0.97fF
C16882 a_27314_57174# a_27406_57174# 0.32fF
C16883 a_30326_15882# a_30418_15516# 0.32fF
C16884 a_2787_30503# a_23747_31055# 0.85fF
C16885 a_38450_70226# a_39454_70226# 0.97fF
C16886 a_19720_7638# a_12899_11471# 0.41fF
C16887 a_5671_21495# a_4792_20443# 0.91fF
C16888 vcm_commonmode a_44474_13508# 0.87fF
C16889 a_49494_59182# a_49494_58178# 1.00fF
C16890 a_24394_61190# ctopp 3.59fF
C16891 ctopn a_28410_10496# 3.59fF
C16892 a_1586_21959# a_3983_20719# 0.83fF
C16893 a_26402_69222# VDD 0.51fF
C16894 a_12725_44527# a_27359_43985# 0.41fF
C16895 a_19374_16520# a_20378_16520# 0.97fF
C16896 vcm_commonmode a_30418_56170# 0.87fF
C16897 a_8361_15529# VDD 0.43fF
C16898 a_26465_48463# VDD 1.04fF
C16899 a_28318_71230# a_28410_71230# 0.32fF
C16900 vcm_commonmode a_33338_69222# 0.31fF
C16901 a_36442_60186# a_36442_59182# 1.00fF
C16902 a_33430_22544# VDD 0.51fF
C16903 a_24394_65206# VDD 0.51fF
C16904 a_24959_30503# a_33694_30761# 1.40fF
C16905 a_25398_63198# a_25398_62194# 1.00fF
C16906 a_40366_11866# a_40458_11500# 0.32fF
C16907 a_2223_28617# a_3355_25071# 0.46fF
C16908 a_16362_57174# ctopp 1.33fF
C16909 a_4191_33449# a_7841_12167# 2.91fF
C16910 a_45478_15516# a_45478_14512# 1.00fF
C16911 vcm_commonmode a_40366_22910# 0.31fF
C16912 a_28410_70226# ctopp 3.58fF
C16913 a_8583_33551# a_12473_37429# 0.74fF
C16914 vcm_commonmode a_31330_65206# 0.31fF
C16915 a_39222_48169# a_12355_65103# 0.40fF
C16916 a_7598_36103# a_7215_36201# 0.32fF
C16917 a_32091_51157# VDD 0.32fF
C16918 a_19282_72234# a_19374_72234# 0.32fF
C16919 a_25744_7638# a_12727_13353# 0.41fF
C16920 a_32772_7638# a_12877_14441# 0.41fF
C16921 a_7571_29199# a_17222_27247# 1.27fF
C16922 a_8583_33551# a_20635_29415# 0.61fF
C16923 a_30418_9492# a_30418_8488# 1.00fF
C16924 a_44382_24918# a_44474_24552# 0.32fF
C16925 ctopn a_23390_15516# 3.59fF
C16926 a_32038_29575# a_28305_28879# 0.46fF
C16927 a_49494_69222# m3_49396_69134# 2.78fF
C16928 a_1761_43567# a_3949_41935# 0.41fF
C16929 vcm_commonmode a_29414_61190# 0.87fF
C16930 a_25398_67214# a_26402_67214# 0.97fF
C16931 a_29414_14512# VDD 0.51fF
C16932 a_24302_55166# VDD 0.35fF
C16933 a_18979_30287# a_14926_31849# 0.57fF
C16934 a_41370_62194# a_41462_62194# 0.32fF
C16935 a_15661_29199# VDD 1.65fF
C16936 a_7479_54439# VDD 7.94fF
C16937 vcm_commonmode a_36350_14878# 0.31fF
C16938 ctopn a_33430_11500# 3.59fF
C16939 a_28547_51175# a_37557_32463# 5.95fF
C16940 a_32951_27247# a_30764_7638# 0.35fF
C16941 a_6372_38279# a_4685_37583# 2.88fF
C16942 a_3668_56311# a_3780_56347# 0.62fF
C16943 a_16744_40517# VDD 1.81fF
C16944 a_44474_69222# a_44474_68218# 1.00fF
C16945 vcm_commonmode a_33430_70226# 0.87fF
C16946 a_34434_8488# a_34434_7484# 1.00fF
C16947 a_34434_23548# VDD 0.52fF
C16948 a_17366_58178# ctopp 3.42fF
C16949 a_29760_7638# a_12985_7663# 0.41fF
C16950 a_31422_66210# VDD 0.51fF
C16951 a_13576_42589# a_23567_42035# 0.87fF
C16952 a_46390_57174# a_46482_57174# 0.32fF
C16953 a_4719_71855# VDD 0.39fF
C16954 a_49402_15882# a_49494_15516# 0.32fF
C16955 vcm_commonmode a_41370_23914# 0.31fF
C16956 vcm_commonmode a_38358_66210# 0.31fF
C16957 a_27406_58178# a_28410_58178# 0.97fF
C16958 a_43470_19532# VDD 0.51fF
C16959 a_19877_52245# VDD 0.67fF
C16960 a_5190_59575# a_9240_53877# 0.66fF
C16961 a_40491_27247# a_12899_11471# 0.41fF
C16962 a_22386_9492# a_23390_9492# 0.97fF
C16963 a_25744_7638# a_10515_23975# 0.41fF
C16964 a_12447_29199# a_7841_12167# 2.26fF
C16965 a_23390_13508# a_23390_12504# 1.00fF
C16966 a_34434_67214# ctopp 3.59fF
C16967 a_38450_16520# a_39454_16520# 0.97fF
C16968 a_32672_49007# a_32856_48463# 0.31fF
C16969 a_47394_71230# a_47486_71230# 0.32fF
C16970 a_8295_47388# a_17039_51157# 0.33fF
C16971 a_6417_62215# a_9424_60949# 0.57fF
C16972 a_44474_63198# a_44474_62194# 1.00fF
C16973 vcm_commonmode a_22386_58178# 0.87fF
C16974 a_41820_41501# VDD 1.86fF
C16975 a_4351_67279# a_11521_66567# 0.34fF
C16976 a_12381_35836# a_12621_36091# 0.84fF
C16977 a_37919_28111# a_12877_14441# 0.41fF
C16978 a_49494_9492# a_49494_8488# 1.00fF
C16979 a_15607_46805# a_4811_34855# 1.64fF
C16980 a_49494_58178# a_49494_57174# 1.00fF
C16981 a_44474_67214# a_45478_67214# 0.97fF
C16982 a_21371_50959# a_2775_46025# 0.54fF
C16983 a_39222_48169# ctopp 2.62fF
C16984 a_23395_32463# a_33694_30761# 0.84fF
C16985 a_1586_45431# a_6559_45205# 0.82fF
C16986 a_13510_44759# VDD 0.63fF
C16987 vcm_commonmode a_39454_67214# 0.87fF
C16988 a_46482_20536# VDD 0.51fF
C16989 a_43270_27791# a_45478_18528# 0.38fF
C16990 a_35438_63198# VDD 0.57fF
C16991 a_5924_69135# VDD 0.61fF
C16992 a_26310_13874# a_26402_13508# 0.32fF
C16993 a_2223_28617# config_1_in[15] 0.52fF
C16994 a_2021_22325# a_23567_44211# 1.28fF
C16995 ctopn VDD 94.48fF
C16996 a_31330_68218# a_31422_68218# 0.32fF
C16997 vcm_commonmode a_42374_63198# 0.31fF
C16998 vcm_commonmode a_32772_7638# 10.34fF
C16999 a_29414_59182# VDD 0.51fF
C17000 a_30418_7484# a_31422_7484# 0.97fF
C17001 a_1867_21263# VDD 0.32fF
C17002 vcm_commonmode a_36442_9492# 0.87fF
C17003 a_33430_64202# ctopp 3.59fF
C17004 ctopn a_38450_13508# 3.59fF
C17005 a_16955_52047# a_20156_49667# 0.61fF
C17006 vcm_commonmode a_36350_59182# 0.31fF
C17007 vcm_commonmode a_16746_22542# 5.36fF
C17008 a_46482_12504# VDD 0.51fF
C17009 a_27271_37455# VDD 0.76fF
C17010 a_30764_7638# a_30418_10496# 0.38fF
C17011 a_13576_37149# a_12473_36341# 2.53fF
C17012 a_4719_71855# a_4885_71855# 0.43fF
C17013 a_9526_61751# VDD 0.52fF
C17014 a_41462_9492# a_42466_9492# 0.97fF
C17015 a_24394_64202# a_25398_64202# 0.97fF
C17016 a_42466_13508# a_42466_12504# 1.00fF
C17017 a_20715_34717# VDD 1.72fF
C17018 vcm_commonmode a_16362_18528# 4.47fF
C17019 a_14258_44527# a_13576_42589# 0.67fF
C17020 a_7797_13885# VDD 0.36fF
C17021 a_8491_41383# VDD 10.01fF
C17022 a_6559_59663# a_4482_57863# 0.39fF
C17023 a_41462_21540# VDD 0.51fF
C17024 vcm_commonmode a_44474_7484# 0.68fF
C17025 a_21382_22544# a_22386_22544# 0.97fF
C17026 a_40050_48463# a_45478_59182# 0.38fF
C17027 a_6095_44807# a_11067_13095# 0.48fF
C17028 a_3137_37589# VDD 0.46fF
C17029 vcm_commonmode a_48398_21906# 0.31fF
C17030 a_42466_69222# ctopp 3.59fF
C17031 a_18370_10496# VDD 0.52fF
C17032 a_15397_39631# VDD 2.09fF
C17033 vcm_commonmode a_38450_64202# 0.87fF
C17034 a_32951_27247# a_33430_8488# 0.38fF
C17035 a_46482_17524# VDD 0.51fF
C17036 a_1923_73087# a_3325_69135# 0.40fF
C17037 a_17507_52047# a_21382_71230# 0.38fF
C17038 a_4758_45369# a_5831_39189# 0.71fF
C17039 a_4298_58951# a_6646_50639# 0.87fF
C17040 a_33430_60186# VDD 0.51fF
C17041 vcm_commonmode a_25306_10862# 0.31fF
C17042 a_6095_44807# a_6559_59879# 1.96fF
C17043 a_12215_31573# VDD 1.12fF
C17044 a_40458_65206# ctopp 3.59fF
C17045 a_32426_67214# a_32426_66210# 1.00fF
C17046 vcm_commonmode a_40366_60186# 0.31fF
C17047 a_39299_48783# a_12981_59343# 0.40fF
C17048 a_28547_51175# a_32426_61190# 0.38fF
C17049 a_2689_65103# a_2794_62697# 0.92fF
C17050 vcm_commonmode a_17366_23548# 1.82fF
C17051 a_12947_71576# ctopp 1.23fF
C17052 a_16510_8760# a_20505_29967# 0.36fF
C17053 a_16955_52047# a_20378_67214# 0.38fF
C17054 a_18611_52047# a_12983_63151# 0.40fF
C17055 a_1987_52484# VDD 0.79fF
C17056 a_1591_59343# VDD 1.66fF
C17057 a_36797_27497# a_37446_24552# 0.46fF
C17058 a_28410_65206# a_28410_64202# 1.00fF
C17059 a_45386_13874# a_45478_13508# 0.32fF
C17060 a_31223_36369# VDD 0.79fF
C17061 vcm_commonmode a_26402_19532# 0.87fF
C17062 a_21371_50959# a_12981_62313# 0.40fF
C17063 a_43267_31055# a_46482_64202# 0.38fF
C17064 vcm_commonmode a_37919_28111# 10.35fF
C17065 a_2079_47546# VDD 0.42fF
C17066 vcm_commonmode a_47486_69222# 0.87fF
C17067 a_33864_28111# a_34434_13508# 0.38fF
C17068 a_9215_58487# VDD 0.53fF
C17069 a_41462_58178# a_41427_52263# 0.38fF
C17070 a_22386_23548# a_22386_22544# 1.00fF
C17071 vcm_commonmode a_20286_15882# 0.31fF
C17072 a_31330_56170# a_31422_56170# 0.32fF
C17073 a_12355_65103# a_16362_65206# 19.89fF
C17074 a_17366_14512# a_18370_14512# 0.97fF
C17075 a_77664_40024# VDD 0.40fF
C17076 a_23390_11500# VDD 0.51fF
C17077 a_12713_41923# VDD 0.78fF
C17078 vcm_commonmode a_45478_65206# 0.87fF
C17079 a_33430_69222# a_34434_69222# 0.97fF
C17080 a_3987_19623# a_4792_20443# 1.08fF
C17081 a_47486_18528# VDD 0.51fF
C17082 a_3891_50645# VDD 0.43fF
C17083 vcm_commonmode a_18278_71230# 0.31fF
C17084 a_28410_61190# a_28410_60186# 1.00fF
C17085 a_27406_24552# VDD 0.60fF
C17086 vcm_commonmode a_30326_11866# 0.31fF
C17087 ctopn a_45478_8488# 3.40fF
C17088 a_7833_66415# VDD 0.88fF
C17089 a_43470_64202# a_44474_64202# 0.97fF
C17090 a_47486_66210# ctopp 3.58fF
C17091 a_5254_67503# a_7803_55509# 1.33fF
C17092 vcm_commonmode a_34342_24918# 0.31fF
C17093 a_23395_52047# a_12727_67753# 0.40fF
C17094 a_28881_52271# a_35568_49525# 0.78fF
C17095 a_37446_55166# VDD 0.60fF
C17096 a_40458_22544# a_41462_22544# 0.97fF
C17097 a_29414_57174# VDD 0.51fF
C17098 a_7210_55081# a_6646_54135# 0.31fF
C17099 a_25787_28327# a_7295_44647# 0.51fF
C17100 a_42709_29199# a_49494_24552# 0.30fF
C17101 a_29760_55394# a_29414_58178# 0.38fF
C17102 a_31422_65206# a_32426_65206# 0.97fF
C17103 a_12985_16367# a_16362_10496# 19.89fF
C17104 a_10317_13647# a_9491_12297# 0.63fF
C17105 a_17585_37477# VDD 1.49fF
C17106 vcm_commonmode a_29414_20536# 0.87fF
C17107 a_16746_68220# ctopp 1.68fF
C17108 vcm_commonmode a_44382_55166# 0.30fF
C17109 vcm_commonmode a_18370_63198# 0.93fF
C17110 a_27406_17524# a_27406_16520# 1.00fF
C17111 vcm_commonmode a_36350_57174# 0.31fF
C17112 a_17668_49007# VDD 0.30fF
C17113 a_37446_72234# a_37446_71230# 1.00fF
C17114 a_3339_43023# a_4674_40277# 0.88fF
C17115 a_2775_46025# a_2419_48783# 0.65fF
C17116 a_22386_23548# a_23390_23548# 0.97fF
C17117 a_6607_42167# a_5631_38127# 0.35fF
C17118 a_31422_56170# a_31422_55166# 1.00fF
C17119 a_16362_11500# a_16746_11498# 2.28fF
C17120 a_14625_30761# VDD 1.44fF
C17121 a_36717_47375# a_30928_49007# 0.31fF
C17122 a_12889_40977# a_13097_40719# 0.41fF
C17123 a_17507_52047# VDD 9.35fF
C17124 a_19374_66210# a_20378_66210# 0.97fF
C17125 a_45478_7484# m3_45380_7346# 2.80fF
C17126 a_5682_69367# a_8772_63927# 0.76fF
C17127 a_9135_27239# a_21382_10496# 0.38fF
C17128 a_7841_12167# a_11067_23759# 1.31fF
C17129 a_7050_53333# a_17843_48981# 0.31fF
C17130 a_11855_51959# VDD 0.58fF
C17131 vcm_commonmode a_21371_52263# 10.02fF
C17132 a_43470_62194# VDD 0.51fF
C17133 a_30326_61190# a_30418_61190# 0.32fF
C17134 a_36797_27497# VDD 6.22fF
C17135 a_42466_55166# m3_42368_55078# 2.81fF
C17136 vcm_commonmode a_29414_12504# 0.87fF
C17137 ctopn a_30418_9492# 3.58fF
C17138 a_2840_66103# a_19478_51959# 0.59fF
C17139 a_47486_65206# a_47486_64202# 1.00fF
C17140 a_13909_35395# VDD 3.14fF
C17141 ctopn a_46482_16520# 3.59fF
C17142 a_11067_47695# a_7841_12167# 1.69fF
C17143 a_13183_52047# a_4758_45369# 0.54fF
C17144 a_40050_48463# a_45478_57174# 0.38fF
C17145 a_4191_33449# a_5831_39189# 2.42fF
C17146 a_19374_71230# a_19374_70226# 1.00fF
C17147 vcm_commonmode a_21290_68218# 0.31fF
C17148 a_29760_55394# a_12901_66959# 0.40fF
C17149 a_31422_19532# a_32426_19532# 0.97fF
C17150 a_3247_20495# a_5085_24759# 0.39fF
C17151 a_41462_23548# a_41462_22544# 1.00fF
C17152 a_41967_31375# a_42466_16520# 0.38fF
C17153 a_5428_63669# VDD 0.54fF
C17154 a_17507_52047# a_26514_47375# 0.39fF
C17155 a_5885_39759# a_6559_39759# 0.36fF
C17156 a_49494_71230# VDD 1.18fF
C17157 a_1761_52815# a_16510_8760# 0.47fF
C17158 a_35438_66210# a_35438_65206# 1.00fF
C17159 a_5254_67503# a_6831_63303# 0.65fF
C17160 a_36442_14512# a_37446_14512# 0.97fF
C17161 a_13837_38772# VDD 1.02fF
C17162 vcm_commonmode a_24394_21540# 0.87fF
C17163 a_1761_9295# VDD 0.32fF
C17164 a_12801_38517# VDD 3.04fF
C17165 a_38450_72234# a_39454_72234# 0.97fF
C17166 a_35601_27497# a_12727_15529# 0.41fF
C17167 a_47486_61190# a_47486_60186# 1.00fF
C17168 a_33338_8854# a_33430_8488# 0.32fF
C17169 a_45478_59182# ctopp 3.59fF
C17170 ctopp m3_32328_55078# 0.38fF
C17171 a_10055_58791# a_39223_32463# 0.41fF
C17172 vcm_commonmode a_29414_17524# 0.87fF
C17173 a_16362_65206# ctopp 1.35fF
C17174 a_12357_37999# a_18127_35797# 0.50fF
C17175 vcm_commonmode a_12727_58255# 6.23fF
C17176 a_5682_69367# a_7265_56053# 0.37fF
C17177 a_30788_28487# a_34267_31599# 0.53fF
C17178 a_34482_29941# a_8491_41383# 1.20fF
C17179 a_28410_13508# VDD 0.51fF
C17180 a_22411_44535# VDD 0.60fF
C17181 a_34342_70226# a_34434_70226# 0.32fF
C17182 a_28881_52271# a_35676_49525# 0.84fF
C17183 a_9031_54135# VDD 0.54fF
C17184 a_31768_7638# a_12985_16367# 0.41fF
C17185 a_33430_62194# a_33430_61190# 1.00fF
C17186 a_24394_10496# a_24394_9492# 1.00fF
C17187 vcm_commonmode a_35346_13874# 0.31fF
C17188 a_17712_7638# a_17366_24552# 0.46fF
C17189 a_40675_27791# a_41462_24552# 0.47fF
C17190 a_31787_36919# VDD 0.61fF
C17191 a_46482_17524# a_46482_16520# 1.00fF
C17192 a_34251_52263# a_41334_29575# 0.31fF
C17193 vcm_commonmode a_21290_56170# 0.31fF
C17194 a_33430_20536# a_33430_19532# 1.00fF
C17195 a_26748_7638# a_12985_19087# 0.41fF
C17196 a_41462_23548# a_42466_23548# 0.97fF
C17197 a_11067_13095# VDD 18.28fF
C17198 a_13643_28327# a_15851_27791# 0.96fF
C17199 a_22151_29941# VDD 0.72fF
C17200 a_25787_28327# a_11067_46823# 1.47fF
C17201 a_16955_52047# a_20635_29415# 0.77fF
C17202 a_12899_2767# a_8491_27023# 1.37fF
C17203 a_38450_66210# a_39454_66210# 0.97fF
C17204 config_1_in[12] config_1_in[11] 0.34fF
C17205 ctopn a_20378_19532# 3.59fF
C17206 a_2473_34293# a_2315_24540# 0.34fF
C17207 a_25787_28327# a_12355_65103# 0.40fF
C17208 ctopn a_24740_7638# 2.62fF
C17209 a_12671_36694# a_12473_36341# 0.30fF
C17210 a_17475_51157# VDD 0.51fF
C17211 a_30764_7638# a_12985_16367# 0.41fF
C17212 a_6559_59879# VDD 6.89fF
C17213 a_49402_61190# a_49494_61190# 0.32fF
C17214 a_12981_59343# a_16362_60186# 1.15fF
C17215 a_7295_25321# VDD 0.41fF
C17216 a_2840_53511# a_6831_63303# 2.09fF
C17217 VDD dummypin[4] 0.96fF
C17218 vcm_commonmode a_30418_18528# 0.87fF
C17219 a_12355_15055# a_8132_53511# 0.91fF
C17220 a_26191_29397# a_26221_29423# 0.31fF
C17221 a_5831_39189# a_3305_38671# 0.46fF
C17222 vcm_commonmode a_20286_61190# 0.31fF
C17223 a_21290_67214# a_21382_67214# 0.32fF
C17224 ctopn a_48490_22544# 3.43fF
C17225 a_3339_30503# a_2787_30503# 0.93fF
C17226 a_13183_52047# a_17366_68218# 0.38fF
C17227 a_38450_71230# a_38450_70226# 1.00fF
C17228 a_16362_55166# VDD 1.22fF
C17229 a_3295_62083# a_7210_55081# 0.38fF
C17230 a_21382_62194# ctopp 3.59fF
C17231 a_19596_40743# a_19245_39747# 0.43fF
C17232 a_17366_70226# VDD 0.58fF
C17233 a_26359_38007# VDD 0.59fF
C17234 vcm_commonmode a_21382_55166# 0.84fF
C17235 VDD result_out[11] 0.80fF
C17236 a_33864_28111# a_34434_7484# 0.34fF
C17237 a_23830_49525# VDD 0.92fF
C17238 vcm_commonmode a_24302_70226# 0.31fF
C17239 a_2686_70223# a_5208_70063# 0.31fF
C17240 a_34434_20536# a_35438_20536# 0.97fF
C17241 a_41370_58178# vcm_commonmode 0.31fF
C17242 vcm_commonmode a_39454_10496# 0.87fF
C17243 a_12947_23413# a_16746_23546# 0.37fF
C17244 a_20635_29415# a_30052_32117# 1.34fF
C17245 a_23390_63198# a_24394_63198# 0.97fF
C17246 ctopn a_44474_14512# 3.59fF
C17247 a_11067_23759# a_11067_21583# 0.36fF
C17248 a_12257_56623# a_16362_56170# 1.15fF
C17249 a_2191_68565# a_3016_60949# 0.54fF
C17250 a_7580_61751# a_7773_63927# 0.71fF
C17251 a_27406_71230# ctopp 3.40fF
C17252 ctopn a_23390_20536# 3.59fF
C17253 a_9491_12297# VDD 1.00fF
C17254 a_23298_58178# a_23390_58178# 0.32fF
C17255 a_8003_72917# a_6921_72943# 0.30fF
C17256 a_1923_73087# a_1950_59887# 2.08fF
C17257 a_18278_9858# a_18370_9492# 0.32fF
C17258 a_43470_10496# a_43470_9492# 1.00fF
C17259 a_3972_25615# VDD 1.98fF
C17260 a_25398_55166# m3_25300_55078# 2.81fF
C17261 a_3295_54421# a_4555_55233# 0.45fF
C17262 a_13005_35823# VDD 6.06fF
C17263 a_35438_8488# VDD 0.58fF
C17264 vcm_commonmode a_26402_62194# 0.87fF
C17265 a_34342_16886# a_34434_16520# 0.32fF
C17266 a_13183_52047# a_17366_56170# 0.38fF
C17267 a_20635_29415# a_15607_46805# 1.35fF
C17268 a_4191_33449# a_7571_29199# 0.47fF
C17269 a_17366_59182# a_18370_59182# 0.97fF
C17270 vcm_commonmode a_42374_8854# 0.31fF
C17271 m3_38352_7346# VDD 0.33fF
C17272 a_43175_28335# a_46482_19532# 0.38fF
C17273 a_3339_32463# a_4903_31849# 0.49fF
C17274 vcm_commonmode a_34434_15516# 0.87fF
C17275 ctopn a_23390_12504# 3.59fF
C17276 a_12707_26159# a_10964_25615# 0.39fF
C17277 a_7464_39215# a_7987_40821# 0.50fF
C17278 a_45478_57174# ctopp 3.58fF
C17279 a_19743_39095# VDD 0.62fF
C17280 a_27406_72234# m3_27308_72146# 2.80fF
C17281 a_1586_66567# a_1770_14441# 0.80fF
C17282 a_4307_67477# a_4211_67655# 0.64fF
C17283 a_49494_13508# m3_49396_13370# 2.78fF
C17284 a_1761_50639# a_1586_45431# 0.82fF
C17285 vcm_commonmode a_32426_71230# 0.86fF
C17286 a_32426_21540# a_32426_20536# 1.00fF
C17287 vcm_commonmode a_44474_11500# 0.87fF
C17288 a_19374_24552# a_19374_23548# 1.00fF
C17289 a_23390_67214# VDD 0.51fF
C17290 a_34434_12504# a_35438_12504# 0.97fF
C17291 a_11619_56615# a_11067_13095# 1.59fF
C17292 a_40366_67214# a_40458_67214# 0.32fF
C17293 a_14287_51175# a_2775_46025# 0.37fF
C17294 a_13183_52047# a_12981_59343# 0.40fF
C17295 a_25787_28327# ctopp 2.67fF
C17296 ctopn a_18370_21540# 3.58fF
C17297 a_2292_43291# a_4842_45467# 0.79fF
C17298 a_1591_44655# VDD 0.42fF
C17299 vcm_commonmode a_30326_67214# 0.31fF
C17300 a_8491_57487# a_4674_57685# 0.34fF
C17301 a_32772_7638# a_12899_11471# 0.41fF
C17302 a_19245_39747# a_14963_39783# 0.43fF
C17303 a_30418_68218# ctopp 3.59fF
C17304 ctopn a_23390_17524# 3.59fF
C17305 a_13183_52047# a_18602_55312# 0.41fF
C17306 a_20378_9492# VDD 0.51fF
C17307 a_24331_39679# VDD 1.18fF
C17308 a_36442_16520# VDD 0.51fF
C17309 a_30609_49159# VDD 0.38fF
C17310 a_26310_7850# a_26402_7484# 0.32fF
C17311 vcm_commonmode a_27314_9858# 0.31fF
C17312 a_42466_63198# a_43470_63198# 0.97fF
C17313 a_7213_62215# a_6559_59663# 0.40fF
C17314 vcm_commonmode a_43378_16886# 0.31fF
C17315 a_4811_34855# a_28841_29575# 0.74fF
C17316 a_7571_29199# a_12447_29199# 4.38fF
C17317 a_1586_66567# a_8772_63927# 1.10fF
C17318 a_12899_10927# a_16362_17524# 19.89fF
C17319 a_8295_47388# a_6559_22671# 0.38fF
C17320 a_3891_50645# a_4057_50645# 0.72fF
C17321 a_33360_51701# VDD 0.76fF
C17322 a_36629_27791# a_12727_13353# 0.41fF
C17323 a_29414_21540# a_30418_21540# 0.97fF
C17324 a_2787_32679# a_4248_29967# 0.58fF
C17325 a_37354_9858# a_37446_9492# 0.32fF
C17326 a_20286_64202# a_20378_64202# 0.32fF
C17327 a_28410_7484# VDD 1.24fF
C17328 a_47486_58178# a_48490_58178# 0.97fF
C17329 a_23763_47381# VDD 0.38fF
C17330 vcm_commonmode a_35438_68218# 0.87fF
C17331 a_36442_59182# a_37446_59182# 0.97fF
C17332 a_17274_22910# a_17366_22544# 0.32fF
C17333 a_22386_64202# VDD 0.51fF
C17334 a_7369_24233# a_10286_26311# 0.39fF
C17335 a_30418_56170# ctopp 3.40fF
C17336 a_3372_70197# VDD 0.31fF
C17337 a_41427_52263# a_41462_59182# 0.38fF
C17338 a_17366_14512# a_17366_13508# 1.00fF
C17339 a_24892_38237# VDD 1.31fF
C17340 ctopn a_24394_18528# 3.59fF
C17341 a_2847_9813# VDD 0.44fF
C17342 a_7097_40303# VDD 0.42fF
C17343 vcm_commonmode a_29322_64202# 0.31fF
C17344 a_34434_17524# a_35438_17524# 0.97fF
C17345 a_44382_72234# a_44474_72234# 0.32fF
C17346 a_23395_52047# a_7841_12167# 0.49fF
C17347 a_21382_60186# a_22386_60186# 0.97fF
C17348 a_10073_23439# VDD 0.89fF
C17349 a_38450_24552# a_38450_23548# 1.00fF
C17350 a_10515_23975# a_16746_23546# 2.28fF
C17351 a_43269_29967# a_12985_19087# 0.41fF
C17352 a_19720_7638# a_12985_7663# 0.41fF
C17353 a_1895_66628# VDD 0.46fF
C17354 a_23390_12504# a_23390_11500# 1.00fF
C17355 a_36199_32143# VDD 0.36fF
C17356 a_28756_55394# a_26397_51183# 0.95fF
C17357 a_28756_55394# a_28410_61190# 0.38fF
C17358 a_36613_48169# a_12981_59343# 0.40fF
C17359 a_2216_28309# a_2223_28617# 1.26fF
C17360 a_8583_33551# a_7841_12167# 3.22fF
C17361 a_12355_15055# a_9865_14441# 0.34fF
C17362 a_8933_22583# a_10394_19605# 0.60fF
C17363 a_37919_28111# a_12899_11471# 0.41fF
C17364 a_7619_62581# VDD 0.46fF
C17365 a_12447_29199# a_32823_29397# 1.60fF
C17366 vcm_commonmode a_49494_13508# 0.89fF
C17367 a_29414_61190# ctopp 3.59fF
C17368 ctopn a_33430_10496# 3.59fF
C17369 a_36629_27791# a_10515_23975# 0.41fF
C17370 a_4528_26159# a_4417_22671# 0.76fF
C17371 a_27752_7638# a_11067_21583# 0.41fF
C17372 a_31422_69222# VDD 0.51fF
C17373 vcm_commonmode a_17274_19898# 0.33fF
C17374 a_38210_30199# a_12899_2767# 0.68fF
C17375 a_11710_58487# a_11521_66567# 1.97fF
C17376 a_14287_51175# a_12981_62313# 0.40fF
C17377 a_41261_28335# a_42466_64202# 0.38fF
C17378 vcm_commonmode a_35438_56170# 0.87fF
C17379 a_5052_14709# VDD 0.41fF
C17380 vcm_commonmode a_38358_69222# 0.31fF
C17381 a_37446_58178# a_36613_48169# 0.38fF
C17382 a_45386_7850# a_45478_7484# 0.32fF
C17383 a_38450_22544# VDD 0.51fF
C17384 vcm_commonmode a_18370_8488# 0.87fF
C17385 a_28756_7638# a_28410_19532# 0.38fF
C17386 a_29414_65206# VDD 0.51fF
C17387 a_1823_62589# a_2794_62697# 0.44fF
C17388 a_21012_30761# VDD 0.78fF
C17389 a_12473_42869# a_30115_38695# 0.74fF
C17390 a_1761_52815# a_1761_30511# 5.00fF
C17391 vcm_commonmode a_45386_22910# 0.31fF
C17392 a_33430_70226# ctopp 3.58fF
C17393 a_15548_30761# a_17554_30663# 0.36fF
C17394 a_10883_11177# VDD 0.71fF
C17395 a_29322_69222# a_29414_69222# 0.32fF
C17396 vcm_commonmode a_36350_65206# 0.31fF
C17397 a_35438_18528# a_35438_17524# 1.00fF
C17398 a_17507_52047# a_21382_72234# 0.34fF
C17399 a_48490_21540# a_49494_21540# 0.97fF
C17400 a_18278_24918# VDD 0.36fF
C17401 a_3987_19623# a_5631_38127# 0.47fF
C17402 a_39362_64202# a_39454_64202# 0.32fF
C17403 ctopn a_28410_15516# 3.59fF
C17404 a_32695_43455# a_30412_42589# 1.22fF
C17405 vcm_commonmode a_34434_61190# 0.87fF
C17406 a_7939_30503# a_25263_29981# 0.31fF
C17407 a_22015_28111# a_18979_30287# 0.43fF
C17408 a_34434_14512# VDD 0.51fF
C17409 a_16955_52047# a_12727_67753# 0.40fF
C17410 config_2_in[12] config_2_in[11] 0.51fF
C17411 a_29322_55166# VDD 0.35fF
C17412 a_36350_22910# a_36442_22544# 0.32fF
C17413 a_3339_43023# a_38115_52263# 0.54fF
C17414 a_25398_10496# a_26402_10496# 0.97fF
C17415 vcm_commonmode a_41370_14878# 0.31fF
C17416 ctopn a_38450_11500# 3.59fF
C17417 a_12202_54599# a_12755_53030# 1.51fF
C17418 a_1761_50639# a_1761_30511# 1.77fF
C17419 a_21371_50959# a_25398_58178# 0.38fF
C17420 a_27314_65206# a_27406_65206# 0.32fF
C17421 a_36442_14512# a_36442_13508# 1.00fF
C17422 a_5547_36495# VDD 0.30fF
C17423 vcm_commonmode a_20286_20902# 0.31fF
C17424 a_2411_26133# config_2_in[7] 0.46fF
C17425 a_40050_48463# a_45478_65206# 0.38fF
C17426 a_3872_15939# VDD 0.62fF
C17427 a_8399_49159# VDD 0.50fF
C17428 a_33430_72234# a_33430_71230# 1.00fF
C17429 vcm_commonmode a_38450_70226# 0.87fF
C17430 a_10515_22671# VDD 11.81fF
C17431 a_6559_22671# a_9260_25045# 0.74fF
C17432 a_40458_60186# a_41462_60186# 0.97fF
C17433 a_39454_23548# VDD 0.52fF
C17434 a_22386_58178# ctopp 3.59fF
C17435 a_40491_27247# a_12985_7663# 0.41fF
C17436 a_18278_23914# a_18370_23548# 0.32fF
C17437 a_36442_66210# VDD 0.51fF
C17438 a_42466_12504# a_42466_11500# 1.00fF
C17439 vcm_commonmode a_19374_16520# 0.87fF
C17440 a_12663_40871# a_12801_38517# 0.47fF
C17441 vcm_commonmode a_46390_23914# 0.31fF
C17442 a_38450_7484# m3_38352_7346# 2.80fF
C17443 a_17711_43439# VDD 1.54fF
C17444 vcm_commonmode a_43378_66210# 0.31fF
C17445 a_29414_70226# a_29414_69222# 1.00fF
C17446 a_35438_18528# a_36442_18528# 0.97fF
C17447 a_48490_19532# VDD 0.54fF
C17448 vcm_commonmode a_19720_55394# 10.02fF
C17449 a_24768_27247# VDD 0.31fF
C17450 a_35438_55166# m3_35340_55078# 2.81fF
C17451 vcm_commonmode a_20286_12870# 0.31fF
C17452 a_10055_58791# a_42718_27497# 0.41fF
C17453 a_39454_67214# ctopp 3.59fF
C17454 a_26523_29199# a_28305_28879# 1.03fF
C17455 a_41427_52263# a_41462_57174# 0.38fF
C17456 a_19807_28111# a_29927_29199# 2.06fF
C17457 a_17599_52263# a_12901_66959# 0.40fF
C17458 a_43267_31055# a_46482_70226# 0.38fF
C17459 a_2419_48783# a_2292_43291# 1.01fF
C17460 a_27314_19898# a_27406_19532# 0.32fF
C17461 a_3339_43023# a_3987_19623# 1.24fF
C17462 a_3969_20175# VDD 0.42fF
C17463 a_2840_66103# a_4482_57863# 0.44fF
C17464 a_28410_11500# a_28410_10496# 1.00fF
C17465 a_18151_52263# a_4443_46607# 0.38fF
C17466 a_1923_59583# a_2163_64381# 0.31fF
C17467 vcm_commonmode a_27406_58178# 0.87fF
C17468 a_32334_14878# a_32426_14512# 0.32fF
C17469 a_4314_40821# VDD 1.86fF
C17470 a_42985_46831# a_48490_66210# 0.38fF
C17471 a_48398_69222# a_48490_69222# 0.32fF
C17472 a_5915_35943# a_8461_32937# 0.67fF
C17473 a_34251_52263# a_36717_47375# 0.87fF
C17474 a_7377_18012# a_12985_19087# 0.32fF
C17475 a_3295_62083# a_4482_57863# 1.22fF
C17476 a_26402_55166# a_27406_55166# 0.97fF
C17477 a_6451_22895# VDD 0.62fF
C17478 a_8491_27023# a_11067_21583# 0.41fF
C17479 vcm_commonmode a_20286_17890# 0.31fF
C17480 a_17507_52047# a_19502_51157# 0.63fF
C17481 a_23567_43123# a_13576_42589# 0.95fF
C17482 a_17366_57174# a_18370_57174# 0.97fF
C17483 a_34251_52263# a_2959_47113# 0.48fF
C17484 a_43362_28879# a_47486_62194# 0.38fF
C17485 a_20378_15516# a_21382_15516# 0.97fF
C17486 a_2339_38129# a_5135_19061# 0.38fF
C17487 a_4811_34855# a_26523_29199# 0.59fF
C17488 a_37427_47893# a_37557_32463# 0.58fF
C17489 vcm_commonmode a_44474_67214# 0.87fF
C17490 a_33864_28111# a_34434_11500# 0.38fF
C17491 a_11619_56615# a_10883_11177# 0.44fF
C17492 a_6743_54447# VDD 0.31fF
C17493 a_5441_72399# a_1923_73087# 0.42fF
C17494 a_9503_26151# a_20378_18528# 0.38fF
C17495 a_40458_63198# VDD 0.57fF
C17496 a_16863_29415# a_12899_3855# 0.37fF
C17497 a_19807_28111# a_28817_29111# 0.38fF
C17498 a_44474_10496# a_45478_10496# 0.97fF
C17499 a_26748_7638# VDD 7.17fF
C17500 a_36629_27791# a_36442_24552# 0.47fF
C17501 a_46390_65206# a_46482_65206# 0.32fF
C17502 a_15775_36965# VDD 0.97fF
C17503 a_12725_44527# a_13716_43047# 0.47fF
C17504 vcm_commonmode a_47394_63198# 0.31fF
C17505 a_2473_34293# a_2787_30503# 0.36fF
C17506 a_18370_71230# a_19374_71230# 0.97fF
C17507 a_34434_59182# VDD 0.51fF
C17508 a_3339_43023# a_20267_30503# 6.26fF
C17509 vcm_commonmode a_41462_9492# 0.87fF
C17510 a_37354_23914# a_37446_23548# 0.32fF
C17511 a_30418_11500# a_31422_11500# 0.97fF
C17512 a_43680_29941# VDD 0.69fF
C17513 a_38450_64202# ctopp 3.59fF
C17514 ctopn a_43470_13508# 3.59fF
C17515 a_42466_72234# VDD 1.36fF
C17516 a_40050_48463# a_12727_58255# 0.40fF
C17517 vcm_commonmode a_41370_59182# 0.31fF
C17518 a_34342_66210# a_34434_66210# 0.32fF
C17519 vcm_commonmode a_21382_22544# 0.87fF
C17520 a_1644_76181# VDD 0.32fF
C17521 a_36395_43177# VDD 0.64fF
C17522 a_48490_70226# a_48490_69222# 1.00fF
C17523 a_21371_52263# a_12355_65103# 0.43fF
C17524 a_19720_7638# a_19374_9492# 0.38fF
C17525 a_25133_37571# a_1761_35407# 1.34fF
C17526 a_11067_47695# a_7571_29199# 0.44fF
C17527 vcm_commonmode a_47486_72234# 0.69fF
C17528 a_32772_7638# a_32426_22544# 0.38fF
C17529 a_34434_24552# a_35438_24552# 0.97fF
C17530 a_28115_34743# VDD 0.59fF
C17531 vcm_commonmode a_21290_18894# 0.31fF
C17532 a_4339_64521# a_7479_54439# 0.59fF
C17533 a_8491_41383# a_5363_30503# 1.02fF
C17534 a_12983_63151# a_16362_67214# 19.89fF
C17535 a_9821_46831# VDD 0.41fF
C17536 a_46390_19898# a_46482_19532# 0.32fF
C17537 a_10515_22671# a_16746_58180# 0.41fF
C17538 a_46482_21540# VDD 0.51fF
C17539 vcm_commonmode a_49494_7484# 0.72fF
C17540 a_41967_31375# a_12727_15529# 0.41fF
C17541 a_31422_62194# a_32426_62194# 0.97fF
C17542 a_47486_11500# a_47486_10496# 1.00fF
C17543 a_32167_29611# VDD 0.69fF
C17544 a_9123_57399# VDD 0.51fF
C17545 vcm_commonmode a_17366_14512# 1.82fF
C17546 a_11803_55311# a_12901_58799# 1.07fF
C17547 a_6559_37583# VDD 0.52fF
C17548 a_47486_69222# ctopp 3.58fF
C17549 a_30052_32117# a_12899_2767# 0.52fF
C17550 a_23390_10496# VDD 0.51fF
C17551 a_26550_40871# VDD 3.36fF
C17552 vcm_commonmode a_43470_64202# 0.87fF
C17553 a_30764_7638# a_30418_15516# 0.38fF
C17554 a_30326_20902# a_30418_20536# 0.32fF
C17555 a_38450_60186# VDD 0.51fF
C17556 a_44474_55166# a_45478_55166# 0.97fF
C17557 vcm_commonmode a_30326_10862# 0.31fF
C17558 a_7987_64213# VDD 0.58fF
C17559 a_27535_30503# a_32970_31145# 0.47fF
C17560 a_7479_54439# a_9547_54421# 0.32fF
C17561 a_19282_63198# a_19374_63198# 0.32fF
C17562 a_24746_31849# VDD 0.49fF
C17563 a_45478_65206# ctopp 3.59fF
C17564 a_11067_23759# a_12546_22351# 0.36fF
C17565 a_23736_7638# a_23390_24552# 0.46fF
C17566 a_12473_42869# a_19967_41781# 1.77fF
C17567 a_36442_57174# a_37446_57174# 0.97fF
C17568 a_6453_71855# VDD 1.69fF
C17569 a_5682_69367# a_4758_45369# 0.31fF
C17570 vcm_commonmode a_45386_60186# 0.31fF
C17571 a_39454_15516# a_40458_15516# 0.97fF
C17572 vcm_commonmode a_22386_23548# 0.87fF
C17573 a_22291_29415# a_18979_30287# 0.47fF
C17574 vcm_commonmode a_19374_66210# 0.87fF
C17575 a_6559_59879# a_19502_51157# 0.52fF
C17576 a_18370_55166# m3_18272_55078# 2.45fF
C17577 vcm_commonmode a_31422_19532# 0.87fF
C17578 a_39454_58178# a_39454_59182# 1.00fF
C17579 vcm_commonmode a_17274_62194# 0.33fF
C17580 a_18370_15516# VDD 0.52fF
C17581 a_6863_42692# VDD 1.52fF
C17582 a_37446_71230# a_38450_71230# 0.97fF
C17583 a_39223_32463# a_12877_14441# 0.41fF
C17584 vcm_commonmode a_25306_15882# 0.31fF
C17585 a_18370_63198# ctopp 3.63fF
C17586 a_12901_66665# VDD 8.03fF
C17587 a_1761_52815# a_17863_36595# 1.21fF
C17588 a_12985_19087# a_16746_8486# 0.41fF
C17589 a_2847_38975# VDD 0.69fF
C17590 a_10515_63143# a_2235_30503# 0.44fF
C17591 a_28410_11500# VDD 0.51fF
C17592 a_6646_50639# VDD 2.08fF
C17593 vcm_commonmode a_23298_71230# 0.31fF
C17594 a_33864_28111# a_12727_15529# 0.41fF
C17595 VDD dummypin[6] 0.93fF
C17596 a_3016_60949# a_1923_54591# 0.38fF
C17597 a_32426_24552# VDD 0.60fF
C17598 vcm_commonmode a_35346_11866# 0.31fF
C17599 a_17366_64202# a_17366_63198# 1.23fF
C17600 a_30326_12870# a_30418_12504# 0.32fF
C17601 a_6243_30662# VDD 2.05fF
C17602 a_12549_44212# a_12473_41781# 1.79fF
C17603 vcm_commonmode a_39362_24918# 0.31fF
C17604 a_21371_52263# ctopp 2.62fF
C17605 a_25398_59182# a_25398_58178# 1.00fF
C17606 a_4215_51157# a_7073_51433# 0.41fF
C17607 a_42466_55166# VDD 0.60fF
C17608 a_16362_63198# VDD 2.48fF
C17609 a_11067_47695# a_11130_22869# 0.55fF
C17610 a_12641_37684# a_13669_38517# 3.40fF
C17611 a_3339_32463# a_13353_30511# 0.66fF
C17612 a_34434_57174# VDD 0.51fF
C17613 vcm_commonmode a_34434_20536# 0.87fF
C17614 vcm_commonmode a_23390_63198# 0.92fF
C17615 a_21382_68218# a_22386_68218# 0.97fF
C17616 vcm_commonmode a_41370_57174# 0.31fF
C17617 a_3607_34639# a_2235_30503# 0.37fF
C17618 a_25419_50959# a_8491_41383# 7.37fF
C17619 a_49402_20902# a_49494_20536# 0.32fF
C17620 a_4298_58951# VDD 2.81fF
C17621 a_38358_63198# a_38450_63198# 0.32fF
C17622 a_29414_57174# a_29414_56170# 1.00fF
C17623 vcm_commonmode a_17366_59182# 1.83fF
C17624 a_6559_22671# a_1761_46287# 2.37fF
C17625 a_40895_43447# VDD 0.61fF
C17626 a_25306_21906# a_25398_21540# 0.32fF
C17627 a_42709_29199# a_12727_15529# 0.40fF
C17628 a_48490_62194# VDD 0.54fF
C17629 a_10680_52245# VDD 8.17fF
C17630 vcm_commonmode a_34434_12504# 0.87fF
C17631 a_12727_58255# ctopp 3.23fF
C17632 ctopn a_35438_9492# 3.58fF
C17633 a_19374_68218# VDD 0.51fF
C17634 a_49494_57174# m3_49396_57086# 2.78fF
C17635 a_22595_35561# VDD 0.63fF
C17636 a_1689_10396# a_3063_9295# 0.32fF
C17637 a_2787_32679# a_5490_41365# 1.36fF
C17638 a_13005_43983# a_16152_43677# 0.49fF
C17639 a_19282_7850# VDD 0.62fF
C17640 a_11803_55311# a_12947_56817# 1.06fF
C17641 a_10407_47607# VDD 0.50fF
C17642 vcm_commonmode a_26310_68218# 0.31fF
C17643 a_32334_59182# a_32426_59182# 0.32fF
C17644 a_11759_63927# VDD 0.38fF
C17645 a_8491_41383# a_23395_32463# 1.52fF
C17646 a_43269_29967# VDD 6.52fF
C17647 a_36613_48169# a_37446_59182# 0.38fF
C17648 a_13909_38659# VDD 1.94fF
C17649 vcm_commonmode a_29414_21540# 0.87fF
C17650 a_2787_30503# a_26191_29397# 0.35fF
C17651 a_29943_41317# VDD 0.90fF
C17652 a_30326_17890# a_30418_17524# 0.32fF
C17653 vcm_commonmode a_47486_58178# 0.87fF
C17654 a_27411_50069# VDD 0.62fF
C17655 a_9503_26151# a_12727_15529# 0.41fF
C17656 a_9135_27239# a_21382_15516# 0.38fF
C17657 a_17274_60186# a_17366_60186# 0.32fF
C17658 a_12869_2741# a_8295_47388# 7.57fF
C17659 a_4443_46607# a_1761_34319# 0.49fF
C17660 a_7773_63927# a_2794_62697# 0.36fF
C17661 a_1823_63677# a_3016_60949# 0.34fF
C17662 a_36442_64202# a_36442_63198# 1.23fF
C17663 a_49402_12870# a_49494_12504# 0.32fF
C17664 vcm_commonmode a_34434_17524# 0.87fF
C17665 a_25971_52263# a_12981_59343# 0.40fF
C17666 vcm_commonmode a_21382_60186# 0.87fF
C17667 a_18151_52263# a_24394_61190# 0.38fF
C17668 a_33430_13508# VDD 0.51fF
C17669 a_39454_58178# a_39454_57174# 1.00fF
C17670 a_30967_44535# VDD 0.59fF
C17671 a_27752_7638# a_27406_9492# 0.38fF
C17672 vcm_commonmode a_39223_32463# 10.35fF
C17673 a_28410_22544# a_28410_21540# 1.00fF
C17674 a_5085_23047# VDD 3.55fF
C17675 a_19374_56170# VDD 0.52fF
C17676 vcm_commonmode a_40366_13874# 0.31fF
C17677 a_25971_52263# a_12447_29199# 0.45fF
C17678 a_27752_7638# a_12546_22351# 0.41fF
C17679 a_35438_13508# a_36442_13508# 0.97fF
C17680 a_12516_7093# a_11067_21583# 0.68fF
C17681 a_40458_68218# a_41462_68218# 0.97fF
C17682 a_38557_32143# a_38450_64202# 0.38fF
C17683 vcm_commonmode a_26310_56170# 0.31fF
C17684 ctopn a_16362_23548# 1.09fF
C17685 a_39299_48783# a_12516_7093# 0.40fF
C17686 a_1761_22895# a_1761_31055# 2.12fF
C17687 a_3325_29967# VDD 1.40fF
C17688 a_48490_57174# a_48490_56170# 1.00fF
C17689 a_21382_56170# a_22386_56170# 0.97fF
C17690 a_5254_67503# a_7773_63927# 0.65fF
C17691 ctopn a_25398_19532# 3.59fF
C17692 a_10055_58791# a_16362_11500# 19.89fF
C17693 a_44382_21906# a_44474_21540# 0.32fF
C17694 a_29760_7638# a_12727_13353# 0.41fF
C17695 a_18370_61190# VDD 0.52fF
C17696 a_25398_58178# a_25398_57174# 1.00fF
C17697 a_2840_66103# a_2775_46025# 1.42fF
C17698 a_1823_63677# a_2944_63400# 0.59fF
C17699 a_22411_34473# VDD 0.61fF
C17700 vcm_commonmode a_35438_18528# 0.87fF
C17701 a_8383_27247# a_6162_28487# 0.70fF
C17702 vcm_commonmode a_25306_61190# 0.31fF
C17703 a_32426_16520# a_32426_15516# 1.00fF
C17704 a_5682_69367# a_8123_56399# 0.54fF
C17705 a_9367_29397# a_10515_32143# 0.62fF
C17706 a_3143_66972# a_6008_69679# 0.38fF
C17707 a_17366_19532# a_17366_18528# 1.00fF
C17708 a_21290_10862# a_21382_10496# 0.32fF
C17709 a_6162_28487# VDD 2.48fF
C17710 a_26402_62194# ctopp 3.59fF
C17711 a_2191_68565# a_2606_41079# 1.63fF
C17712 a_22386_70226# VDD 0.51fF
C17713 a_17507_52047# a_21382_58178# 0.38fF
C17714 a_37076_37253# VDD 1.80fF
C17715 a_39454_58178# VDD 0.51fF
C17716 vcm_commonmode a_26402_55166# 0.84fF
C17717 a_1591_44655# a_1757_44655# 0.72fF
C17718 a_7244_39189# VDD 0.99fF
C17719 a_41427_52263# a_41462_65206# 0.38fF
C17720 a_49402_17890# a_49494_17524# 0.32fF
C17721 vcm_commonmode a_17366_57174# 1.83fF
C17722 a_19807_28111# VDD 15.77fF
C17723 a_29414_72234# a_29414_71230# 1.00fF
C17724 vcm_commonmode a_29322_70226# 0.31fF
C17725 a_39222_48169# a_12907_56399# 0.83fF
C17726 a_2021_17973# a_2317_28892# 0.61fF
C17727 a_2099_59861# a_2124_59459# 0.37fF
C17728 a_36350_60186# a_36442_60186# 0.32fF
C17729 vcm_commonmode a_44474_10496# 0.87fF
C17730 a_21187_29415# a_14926_31849# 0.50fF
C17731 a_4443_46607# a_3339_30503# 0.31fF
C17732 a_13643_28327# a_33694_30761# 0.54fF
C17733 a_2099_59861# a_5449_25071# 0.36fF
C17734 a_28817_29111# a_37699_27221# 0.69fF
C17735 a_10949_72719# VDD 0.39fF
C17736 a_32426_71230# ctopp 3.40fF
C17737 ctopn a_28410_20536# 3.59fF
C17738 a_31422_7484# m3_31324_7346# 2.80fF
C17739 a_15548_30761# a_20881_28111# 0.90fF
C17740 a_7571_29199# a_18539_47617# 0.63fF
C17741 a_31330_18894# a_31422_18528# 0.32fF
C17742 a_47486_22544# a_47486_21540# 1.00fF
C17743 a_20378_61190# a_21382_61190# 0.97fF
C17744 a_29760_7638# a_10515_23975# 0.41fF
C17745 a_7213_62215# a_3295_62083# 0.52fF
C17746 a_37527_29397# a_28841_29575# 0.63fF
C17747 a_2539_42106# a_2235_41941# 0.32fF
C17748 a_40458_8488# VDD 0.58fF
C17749 vcm_commonmode a_31422_62194# 0.87fF
C17750 a_26402_68218# a_26402_67214# 1.00fF
C17751 a_36613_48169# a_37446_57174# 0.38fF
C17752 a_7000_43541# a_17488_48731# 0.51fF
C17753 a_40599_47919# VDD 0.43fF
C17754 a_41261_28335# a_42466_70226# 0.38fF
C17755 a_7377_18012# VDD 3.48fF
C17756 vcm_commonmode a_47394_8854# 0.31fF
C17757 a_20635_29415# a_26523_29199# 0.57fF
C17758 a_2339_38129# a_2012_33927# 0.52fF
C17759 vcm_commonmode a_39454_15516# 0.87fF
C17760 ctopn a_28410_12504# 3.59fF
C17761 a_12473_42869# a_1761_27791# 1.15fF
C17762 a_40458_56170# a_41462_56170# 0.97fF
C17763 config_2_in[3] config_2_in[4] 0.31fF
C17764 vcm_commonmode a_18278_58178# 0.31fF
C17765 a_47486_24552# m2_48260_24282# 0.92fF
C17766 a_30418_72234# m3_30320_72146# 2.80fF
C17767 a_32029_41829# VDD 1.86fF
C17768 a_11803_55311# a_2840_66103# 1.80fF
C17769 a_39299_48783# a_44474_66210# 0.38fF
C17770 a_22181_50645# VDD 0.38fF
C17771 vcm_commonmode a_37446_71230# 0.86fF
C17772 a_31422_72234# a_32426_72234# 0.97fF
C17773 a_23390_8488# a_24394_8488# 0.97fF
C17774 a_22294_55166# a_22386_55166# 0.32fF
C17775 vcm_commonmode a_49494_11500# 0.90fF
C17776 a_8491_27023# a_12546_22351# 0.46fF
C17777 a_32772_7638# a_12985_7663# 0.41fF
C17778 a_28410_67214# VDD 0.51fF
C17779 a_20905_32143# VDD 1.28fF
C17780 a_9731_22895# a_12631_28585# 0.30fF
C17781 a_41967_31375# a_40491_27247# 1.18fF
C17782 a_12473_42869# a_19004_40413# 1.89fF
C17783 a_8583_33551# a_32823_29397# 0.78fF
C17784 a_41872_29423# a_43470_62194# 0.38fF
C17785 a_12983_63151# a_10975_66407# 23.50fF
C17786 a_16362_15516# a_16746_15514# 2.28fF
C17787 ctopn a_23390_21540# 3.59fF
C17788 a_1586_45431# a_2927_39733# 0.48fF
C17789 a_2313_12015# VDD 0.69fF
C17790 a_24394_70226# a_25398_70226# 0.97fF
C17791 vcm_commonmode a_35346_67214# 0.31fF
C17792 a_36442_19532# a_36442_18528# 1.00fF
C17793 a_41462_58178# a_42466_58178# 0.97fF
C17794 a_11067_21583# a_16746_21538# 0.41fF
C17795 a_40366_10862# a_40458_10496# 0.32fF
C17796 vcm_commonmode a_16362_13508# 4.47fF
C17797 a_3143_22364# a_2411_19605# 0.44fF
C17798 a_11067_13095# a_4339_64521# 0.75fF
C17799 a_35438_68218# ctopp 3.59fF
C17800 ctopn a_28410_17524# 3.59fF
C17801 a_25398_9492# VDD 0.51fF
C17802 a_41462_16520# VDD 0.51fF
C17803 a_12947_71576# a_12907_56399# 0.31fF
C17804 a_22386_60186# a_22386_59182# 1.00fF
C17805 vcm_commonmode a_32334_9858# 0.31fF
C17806 m3_38352_72146# VDD 0.33fF
C17807 a_7000_65595# VDD 0.63fF
C17808 a_8123_56399# a_4215_51157# 0.50fF
C17809 a_4339_64521# a_6559_59879# 1.69fF
C17810 a_26310_11866# a_26402_11500# 0.32fF
C17811 vcm_commonmode a_48398_16886# 0.31fF
C17812 a_35438_72234# VDD 1.23fF
C17813 a_38557_32143# a_12727_58255# 0.40fF
C17814 a_31422_15516# a_31422_14512# 1.00fF
C17815 vcm_commonmode m3_16264_67126# 3.21fF
C17816 a_21663_42943# VDD 0.92fF
C17817 a_19720_55394# a_12355_65103# 0.40fF
C17818 a_2216_28309# a_2473_34293# 1.18fF
C17819 a_33748_51727# VDD 0.45fF
C17820 vcm_commonmode a_40458_72234# 0.69fF
C17821 a_11067_13095# a_3247_20495# 0.79fF
C17822 a_2775_46025# a_14831_50095# 0.53fF
C17823 a_39454_61190# a_40458_61190# 0.97fF
C17824 a_30326_24918# a_30418_24552# 0.32fF
C17825 a_7061_34319# VDD 0.60fF
C17826 a_33430_7484# VDD 1.62fF
C17827 a_45478_68218# a_45478_67214# 1.00fF
C17828 a_4259_32687# a_4425_32687# 0.43fF
C17829 vcm_commonmode a_40458_68218# 0.87fF
C17830 a_27406_64202# VDD 0.51fF
C17831 a_27314_62194# a_27406_62194# 0.32fF
C17832 a_9529_28335# VDD 5.72fF
C17833 a_19720_7638# a_9503_26151# 3.17fF
C17834 a_35438_56170# ctopp 3.40fF
C17835 ctopn a_29414_18528# 3.59fF
C17836 vcm_commonmode a_34342_64202# 0.31fF
C17837 a_30418_69222# a_30418_68218# 1.00fF
C17838 a_13097_36367# a_1761_34319# 3.49fF
C17839 a_43267_31055# a_46482_72234# 0.34fF
C17840 a_42718_27497# a_12877_14441# 0.41fF
C17841 a_42466_8488# a_43470_8488# 0.97fF
C17842 a_20378_8488# a_20378_7484# 1.00fF
C17843 a_40366_55166# a_40458_55166# 0.32fF
C17844 a_37919_28111# a_12985_7663# 0.41fF
C17845 a_11067_67279# a_2419_48783# 3.13fF
C17846 a_32334_57174# a_32426_57174# 0.32fF
C17847 a_1591_66415# a_1923_59583# 0.33fF
C17848 a_35346_15882# a_35438_15516# 0.32fF
C17849 a_4674_40277# config_2_in[7] 0.31fF
C17850 a_5791_43541# VDD 0.36fF
C17851 a_43470_70226# a_44474_70226# 0.97fF
C17852 a_12985_19087# VDD 8.02fF
C17853 a_34434_61190# ctopp 3.59fF
C17854 ctopn a_38450_10496# 3.59fF
C17855 a_36442_69222# VDD 0.51fF
C17856 a_17488_48731# a_5915_35943# 0.65fF
C17857 vcm_commonmode a_22294_19898# 0.31fF
C17858 a_16746_8486# VDD 33.50fF
C17859 a_24394_16520# a_25398_16520# 0.97fF
C17860 vcm_commonmode a_40458_56170# 0.87fF
C17861 a_2339_38129# a_4839_21495# 0.75fF
C17862 a_22015_28111# a_18703_29199# 0.82fF
C17863 a_19807_28111# a_34482_29941# 0.43fF
C17864 a_29927_29199# VDD 7.42fF
C17865 a_33338_71230# a_33430_71230# 0.32fF
C17866 vcm_commonmode a_43378_69222# 0.31fF
C17867 a_41462_60186# a_41462_59182# 1.00fF
C17868 a_43470_22544# VDD 0.51fF
C17869 vcm_commonmode a_23390_8488# 0.86fF
C17870 a_30764_7638# a_30418_20536# 0.38fF
C17871 a_2411_19605# a_4792_20443# 0.30fF
C17872 a_34434_65206# VDD 0.51fF
C17873 a_30418_63198# a_30418_62194# 1.00fF
C17874 a_45386_11866# a_45478_11500# 0.32fF
C17875 a_4351_67279# a_17039_51157# 0.89fF
C17876 a_38450_70226# ctopp 3.58fF
C17877 vcm_commonmode m3_16264_14374# 3.21fF
C17878 a_14625_30761# a_18162_31055# 0.63fF
C17879 a_42283_42359# VDD 0.67fF
C17880 vcm_commonmode a_41370_65206# 0.31fF
C17881 a_1761_27791# a_15968_36061# 2.45fF
C17882 a_2021_22325# a_4248_29967# 0.46fF
C17883 a_35438_9492# a_35438_8488# 1.00fF
C17884 a_23298_24918# VDD 0.36fF
C17885 a_10379_66389# VDD 0.70fF
C17886 a_1683_33237# VDD 0.45fF
C17887 ctopn a_33430_15516# 3.59fF
C17888 a_1689_10396# config_2_in[0] 0.39fF
C17889 a_30418_67214# a_31422_67214# 0.97fF
C17890 vcm_commonmode a_39454_61190# 0.87fF
C17891 a_19720_55394# ctopp 2.62fF
C17892 a_39454_14512# VDD 0.51fF
C17893 a_42985_46831# a_48490_69222# 0.38fF
C17894 a_30764_7638# a_30418_12504# 0.38fF
C17895 a_18370_20536# VDD 0.52fF
C17896 a_33430_55166# VDD 0.60fF
C17897 a_46390_62194# a_46482_62194# 0.32fF
C17898 a_28817_29111# VDD 3.40fF
C17899 vcm_commonmode a_46390_14878# 0.31fF
C17900 ctopn a_43470_11500# 3.59fF
C17901 vcm_commonmode a_25306_20902# 0.31fF
C17902 a_2787_30503# a_26350_28585# 1.05fF
C17903 a_13909_39747# VDD 8.96fF
C17904 a_17274_68218# a_17366_68218# 0.32fF
C17905 a_49494_69222# a_49494_68218# 1.00fF
C17906 ctopn a_47486_24552# 0.30fF
C17907 a_9392_48981# VDD 0.56fF
C17908 a_13183_52047# a_12516_7093# 0.41fF
C17909 vcm_commonmode a_43470_70226# 0.87fF
C17910 a_5535_18012# a_8539_18231# 0.37fF
C17911 a_39454_8488# a_39454_7484# 1.00fF
C17912 a_16362_7484# a_17366_7484# 0.97fF
C17913 a_44474_23548# VDD 0.52fF
C17914 a_27406_58178# ctopp 3.59fF
C17915 a_11067_13095# a_9963_50959# 0.65fF
C17916 a_41462_66210# VDD 0.51fF
C17917 VDD config_1_in[2] 1.04fF
C17918 a_8753_31055# VDD 1.39fF
C17919 vcm_commonmode a_24394_16520# 0.87fF
C17920 a_12899_3311# a_33864_28111# 0.51fF
C17921 a_13576_42589# a_12473_41781# 1.36fF
C17922 a_2004_42453# config_2_in[0] 1.54fF
C17923 a_3339_43023# m2_48260_54946# 0.36fF
C17924 a_18370_12504# VDD 0.52fF
C17925 a_27999_41495# VDD 0.96fF
C17926 vcm_commonmode a_48398_66210# 0.31fF
C17927 a_2689_65103# a_3024_67191# 0.47fF
C17928 a_33864_28111# a_34434_10496# 0.38fF
C17929 a_32426_58178# a_33430_58178# 0.97fF
C17930 a_30764_7638# a_30418_17524# 0.38fF
C17931 a_27406_9492# a_28410_9492# 0.97fF
C17932 a_1823_54973# VDD 1.67fF
C17933 vcm_commonmode a_25306_12870# 0.31fF
C17934 a_9914_68279# VDD 0.77fF
C17935 a_28410_13508# a_28410_12504# 1.00fF
C17936 a_44474_67214# ctopp 3.59fF
C17937 a_43470_16520# a_44474_16520# 0.97fF
C17938 vcm_commonmode a_42718_27497# 10.41fF
C17939 vcm_commonmode a_16362_68218# 4.47fF
C17940 a_3339_43023# a_12621_44099# 0.37fF
C17941 vcm_commonmode a_16362_7484# 1.71fF
C17942 a_31768_7638# a_31422_18528# 0.38fF
C17943 a_49494_63198# a_49494_62194# 1.00fF
C17944 vcm_commonmode a_32426_58178# 0.87fF
C17945 a_43267_31055# a_12901_58799# 0.40fF
C17946 a_25787_28327# a_33430_59182# 0.38fF
C17947 vcm_commonmode a_20286_21906# 0.31fF
C17948 VDD config_2_in[5] 0.75fF
C17949 a_18370_17524# VDD 0.52fF
C17950 a_4031_50247# VDD 0.41fF
C17951 a_37354_72234# a_37446_72234# 0.32fF
C17952 a_39223_32463# a_12899_11471# 0.41fF
C17953 a_11067_23759# a_12985_16367# 0.36fF
C17954 a_26413_31055# VDD 0.41fF
C17955 vcm_commonmode a_25306_17890# 0.31fF
C17956 a_7755_74581# VDD 0.50fF
C17957 a_16955_52047# a_20378_61190# 0.38fF
C17958 a_18611_52047# a_12981_59343# 0.40fF
C17959 a_18370_67214# a_18370_66210# 1.00fF
C17960 a_16928_44007# VDD 1.62fF
C17961 vcm_commonmode a_49494_67214# 0.91fF
C17962 a_76971_38925# inp_analog 1.02fF
C17963 a_45478_63198# VDD 0.57fF
C17964 a_37699_27221# VDD 0.73fF
C17965 a_3005_56079# VDD 0.49fF
C17966 a_31330_13874# a_31422_13508# 0.32fF
C17967 a_22411_36919# VDD 0.60fF
C17968 a_3987_19623# a_1803_20719# 0.36fF
C17969 a_34780_56398# a_34434_64202# 0.38fF
C17970 a_36350_68218# a_36442_68218# 0.32fF
C17971 a_2283_15797# a_3019_13621# 0.49fF
C17972 vcm_commonmode a_16362_56170# 4.45fF
C17973 a_3247_20495# a_6608_19319# 0.31fF
C17974 vcm_commonmode a_19374_69222# 0.87fF
C17975 a_36613_48169# a_12516_7093# 0.40fF
C17976 a_10515_23975# a_12727_15529# 0.32fF
C17977 a_39454_59182# VDD 0.51fF
C17978 a_35438_7484# a_36442_7484# 0.97fF
C17979 vcm_commonmode a_46482_9492# 0.87fF
C17980 a_9135_27239# a_21382_20536# 0.38fF
C17981 a_6095_44807# VDD 7.48fF
C17982 a_8273_42479# a_5915_35943# 1.26fF
C17983 a_43470_64202# ctopp 3.59fF
C17984 ctopn a_48490_13508# 3.43fF
C17985 a_41427_52263# a_20359_29199# 0.50fF
C17986 a_3301_27791# a_3325_18543# 0.44fF
C17987 a_17274_56170# a_17366_56170# 0.32fF
C17988 a_46390_72234# VDD 0.61fF
C17989 vcm_commonmode a_46390_59182# 0.31fF
C17990 vcm_commonmode a_26402_22544# 0.87fF
C17991 ctopn a_16362_19532# 1.35fF
C17992 a_19374_69222# a_20378_69222# 0.97fF
C17993 vcm_commonmode a_17366_65206# 1.83fF
C17994 a_19374_18528# VDD 0.51fF
C17995 a_11067_63143# a_7571_29199# 5.86fF
C17996 a_46482_9492# a_47486_9492# 0.97fF
C17997 a_4149_24527# VDD 0.80fF
C17998 ctopn a_17366_8488# 3.24fF
C17999 a_29414_64202# a_30418_64202# 0.97fF
C18000 a_1923_59583# a_2775_46025# 0.49fF
C18001 a_7580_61751# a_7107_58487# 0.36fF
C18002 a_47486_13508# a_47486_12504# 1.00fF
C18003 vcm_commonmode a_26310_18894# 0.31fF
C18004 a_19374_66210# ctopp 3.59fF
C18005 a_34482_29941# a_29927_29199# 0.68fF
C18006 a_10317_13647# VDD 0.69fF
C18007 ctopn m3_17268_23410# 0.46fF
C18008 a_4482_57863# a_21169_49007# 0.60fF
C18009 a_9135_27239# a_21382_12504# 0.38fF
C18010 a_26402_22544# a_27406_22544# 0.97fF
C18011 a_7295_44647# a_32970_31145# 0.93fF
C18012 a_16362_10496# a_16746_10494# 2.28fF
C18013 vcm_commonmode a_22386_14512# 0.87fF
C18014 a_17366_65206# a_18370_65206# 0.97fF
C18015 a_18811_38053# VDD 0.89fF
.ends

