VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_top
  CLASS BLOCK ;
  FOREIGN adc_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 423.500 BY 403.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 399.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 425.280 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 397.680 425.280 399.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.680 3.280 425.280 399.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.720 -0.020 18.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.720 -0.020 42.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 -0.020 66.320 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.720 134.310 90.320 176.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.720 225.845 90.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.720 134.310 114.320 176.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.720 225.845 114.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.720 134.310 138.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 160.720 134.310 162.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 134.310 186.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 134.310 210.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.720 134.310 234.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.720 134.310 258.320 181.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.720 216.190 258.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 280.720 134.310 282.320 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.720 196.960 306.320 225.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.720 196.960 330.320 225.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 352.720 196.960 354.320 225.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 376.720 174.300 378.320 204.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.720 -0.020 402.320 402.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 34.080 79.800 35.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 58.080 79.800 59.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 82.080 79.800 83.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 106.080 79.800 107.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 130.080 79.800 131.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 154.080 428.580 155.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 178.080 428.580 179.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 202.080 428.580 203.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 226.080 428.580 227.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 250.080 428.580 251.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 274.080 79.800 275.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 298.080 79.800 299.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 322.080 79.800 323.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 346.080 79.800 347.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 370.080 79.800 371.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 34.080 428.580 35.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 58.080 428.580 59.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 82.080 428.580 83.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 106.080 428.580 107.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 130.080 428.580 131.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 274.080 428.580 275.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 298.080 428.580 299.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 322.080 428.580 323.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 346.080 428.580 347.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 370.080 428.580 371.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 409.060 10.640 410.660 391.920 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 402.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 428.580 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 400.980 428.580 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.980 -0.020 428.580 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.020 -0.020 21.620 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.020 -0.020 45.620 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.020 -0.020 69.620 176.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.020 225.845 69.620 402.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.020 134.310 93.620 176.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.020 225.845 93.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.020 134.310 117.620 176.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.020 225.845 117.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 140.020 134.310 141.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.020 134.310 165.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 134.310 189.620 166.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 229.660 189.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.020 134.310 213.620 166.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.020 229.660 213.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 236.020 134.310 237.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.020 134.310 261.620 181.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.020 216.190 261.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.020 134.310 285.620 266.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.020 196.960 309.620 225.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.020 196.960 333.620 225.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 356.020 196.960 357.620 225.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 -0.020 405.620 402.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 37.380 79.800 38.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 61.380 79.800 62.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 85.380 79.800 86.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 109.380 79.800 110.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 133.380 428.580 134.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 157.380 428.580 158.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 181.380 428.580 182.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 205.380 428.580 206.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 229.380 428.580 230.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 253.380 428.580 254.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 277.380 79.800 278.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 301.380 79.800 302.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 325.380 79.800 326.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 349.380 79.800 350.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 373.380 428.580 374.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 37.380 428.580 38.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 61.380 428.580 62.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 85.380 428.580 86.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 109.380 428.580 110.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 277.380 428.580 278.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 301.380 428.580 302.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 325.380 428.580 326.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.560 349.380 428.580 350.980 ;
    END
  END VSS
  PIN clk_vcm
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 179.560 423.500 180.160 ;
    END
  END clk_vcm
  PIN config_1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END config_1_in[0]
  PIN config_1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END config_1_in[10]
  PIN config_1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END config_1_in[11]
  PIN config_1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END config_1_in[12]
  PIN config_1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END config_1_in[13]
  PIN config_1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END config_1_in[14]
  PIN config_1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END config_1_in[15]
  PIN config_1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END config_1_in[1]
  PIN config_1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END config_1_in[2]
  PIN config_1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END config_1_in[3]
  PIN config_1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END config_1_in[4]
  PIN config_1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END config_1_in[5]
  PIN config_1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END config_1_in[6]
  PIN config_1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END config_1_in[7]
  PIN config_1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END config_1_in[8]
  PIN config_1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END config_1_in[9]
  PIN config_2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END config_2_in[0]
  PIN config_2_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END config_2_in[10]
  PIN config_2_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END config_2_in[11]
  PIN config_2_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END config_2_in[12]
  PIN config_2_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END config_2_in[13]
  PIN config_2_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END config_2_in[14]
  PIN config_2_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END config_2_in[15]
  PIN config_2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END config_2_in[1]
  PIN config_2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END config_2_in[2]
  PIN config_2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END config_2_in[3]
  PIN config_2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END config_2_in[4]
  PIN config_2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END config_2_in[5]
  PIN config_2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END config_2_in[6]
  PIN config_2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END config_2_in[7]
  PIN config_2_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END config_2_in[8]
  PIN config_2_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END config_2_in[9]
  PIN conversion_finished_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END conversion_finished_out
  PIN dummypin[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 390.360 423.500 390.960 ;
    END
  END dummypin[0]
  PIN dummypin[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 116.320 423.500 116.920 ;
    END
  END dummypin[10]
  PIN dummypin[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 95.240 423.500 95.840 ;
    END
  END dummypin[11]
  PIN dummypin[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 74.160 423.500 74.760 ;
    END
  END dummypin[12]
  PIN dummypin[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 53.080 423.500 53.680 ;
    END
  END dummypin[13]
  PIN dummypin[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 32.000 423.500 32.600 ;
    END
  END dummypin[14]
  PIN dummypin[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 10.920 423.500 11.520 ;
    END
  END dummypin[15]
  PIN dummypin[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 369.280 423.500 369.880 ;
    END
  END dummypin[1]
  PIN dummypin[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 348.200 423.500 348.800 ;
    END
  END dummypin[2]
  PIN dummypin[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 327.120 423.500 327.720 ;
    END
  END dummypin[3]
  PIN dummypin[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 306.040 423.500 306.640 ;
    END
  END dummypin[4]
  PIN dummypin[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 284.960 423.500 285.560 ;
    END
  END dummypin[5]
  PIN dummypin[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 263.880 423.500 264.480 ;
    END
  END dummypin[6]
  PIN dummypin[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 242.800 423.500 243.400 ;
    END
  END dummypin[7]
  PIN dummypin[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 158.480 423.500 159.080 ;
    END
  END dummypin[8]
  PIN dummypin[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 137.400 423.500 138.000 ;
    END
  END dummypin[9]
  PIN inn_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 200.640 423.500 201.240 ;
    END
  END inn_analog
  PIN inp_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.500 221.720 423.500 222.320 ;
    END
  END inp_analog
  PIN result_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END result_out[0]
  PIN result_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END result_out[10]
  PIN result_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END result_out[11]
  PIN result_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END result_out[12]
  PIN result_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END result_out[13]
  PIN result_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END result_out[14]
  PIN result_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END result_out[15]
  PIN result_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END result_out[1]
  PIN result_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END result_out[2]
  PIN result_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END result_out[3]
  PIN result_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END result_out[4]
  PIN result_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END result_out[5]
  PIN result_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END result_out[6]
  PIN result_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END result_out[7]
  PIN result_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END result_out[8]
  PIN result_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END result_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END rst_n
  PIN start_conversion_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END start_conversion_in
  OBS
      LAYER li1 ;
        RECT 5.520 10.000 417.680 391.765 ;
      LAYER met1 ;
        RECT 5.520 8.880 417.680 391.920 ;
      LAYER met2 ;
        RECT 6.530 8.850 415.290 391.865 ;
      LAYER met3 ;
        RECT 4.000 391.360 419.500 391.845 ;
        RECT 4.000 389.960 419.100 391.360 ;
        RECT 4.000 388.640 419.500 389.960 ;
        RECT 4.400 387.240 419.500 388.640 ;
        RECT 4.000 381.160 419.500 387.240 ;
        RECT 4.400 379.760 419.500 381.160 ;
        RECT 4.000 373.680 419.500 379.760 ;
        RECT 4.400 372.280 419.500 373.680 ;
        RECT 4.000 370.280 419.500 372.280 ;
        RECT 4.000 368.880 419.100 370.280 ;
        RECT 4.000 366.200 419.500 368.880 ;
        RECT 4.400 364.800 419.500 366.200 ;
        RECT 4.000 358.720 419.500 364.800 ;
        RECT 4.400 357.320 419.500 358.720 ;
        RECT 4.000 351.240 419.500 357.320 ;
        RECT 4.400 349.840 419.500 351.240 ;
        RECT 4.000 349.200 419.500 349.840 ;
        RECT 4.000 347.800 419.100 349.200 ;
        RECT 4.000 343.760 419.500 347.800 ;
        RECT 4.400 342.360 419.500 343.760 ;
        RECT 4.000 336.280 419.500 342.360 ;
        RECT 4.400 334.880 419.500 336.280 ;
        RECT 4.000 328.800 419.500 334.880 ;
        RECT 4.400 328.120 419.500 328.800 ;
        RECT 4.400 327.400 419.100 328.120 ;
        RECT 4.000 326.720 419.100 327.400 ;
        RECT 4.000 321.320 419.500 326.720 ;
        RECT 4.400 319.920 419.500 321.320 ;
        RECT 4.000 313.840 419.500 319.920 ;
        RECT 4.400 312.440 419.500 313.840 ;
        RECT 4.000 307.040 419.500 312.440 ;
        RECT 4.000 306.360 419.100 307.040 ;
        RECT 4.400 305.640 419.100 306.360 ;
        RECT 4.400 304.960 419.500 305.640 ;
        RECT 4.000 298.880 419.500 304.960 ;
        RECT 4.400 297.480 419.500 298.880 ;
        RECT 4.000 291.400 419.500 297.480 ;
        RECT 4.400 290.000 419.500 291.400 ;
        RECT 4.000 285.960 419.500 290.000 ;
        RECT 4.000 284.560 419.100 285.960 ;
        RECT 4.000 283.920 419.500 284.560 ;
        RECT 4.400 282.520 419.500 283.920 ;
        RECT 4.000 276.440 419.500 282.520 ;
        RECT 4.400 275.040 419.500 276.440 ;
        RECT 4.000 268.960 419.500 275.040 ;
        RECT 4.400 267.560 419.500 268.960 ;
        RECT 4.000 264.880 419.500 267.560 ;
        RECT 4.000 263.480 419.100 264.880 ;
        RECT 4.000 261.480 419.500 263.480 ;
        RECT 4.400 260.080 419.500 261.480 ;
        RECT 4.000 254.000 419.500 260.080 ;
        RECT 4.400 252.600 419.500 254.000 ;
        RECT 4.000 246.520 419.500 252.600 ;
        RECT 4.400 245.120 419.500 246.520 ;
        RECT 4.000 243.800 419.500 245.120 ;
        RECT 4.000 242.400 419.100 243.800 ;
        RECT 4.000 239.040 419.500 242.400 ;
        RECT 4.400 237.640 419.500 239.040 ;
        RECT 4.000 231.560 419.500 237.640 ;
        RECT 4.400 230.160 419.500 231.560 ;
        RECT 4.000 224.080 419.500 230.160 ;
        RECT 4.400 222.720 419.500 224.080 ;
        RECT 4.400 222.680 419.100 222.720 ;
        RECT 4.000 221.320 419.100 222.680 ;
        RECT 4.000 216.600 419.500 221.320 ;
        RECT 4.400 215.200 419.500 216.600 ;
        RECT 4.000 209.120 419.500 215.200 ;
        RECT 4.400 207.720 419.500 209.120 ;
        RECT 4.000 201.640 419.500 207.720 ;
        RECT 4.400 200.240 419.100 201.640 ;
        RECT 4.000 194.160 419.500 200.240 ;
        RECT 4.400 192.760 419.500 194.160 ;
        RECT 4.000 186.680 419.500 192.760 ;
        RECT 4.400 185.280 419.500 186.680 ;
        RECT 4.000 180.560 419.500 185.280 ;
        RECT 4.000 179.200 419.100 180.560 ;
        RECT 4.400 179.160 419.100 179.200 ;
        RECT 4.400 177.800 419.500 179.160 ;
        RECT 4.000 171.720 419.500 177.800 ;
        RECT 4.400 170.320 419.500 171.720 ;
        RECT 4.000 164.240 419.500 170.320 ;
        RECT 4.400 162.840 419.500 164.240 ;
        RECT 4.000 159.480 419.500 162.840 ;
        RECT 4.000 158.080 419.100 159.480 ;
        RECT 4.000 156.760 419.500 158.080 ;
        RECT 4.400 155.360 419.500 156.760 ;
        RECT 4.000 149.280 419.500 155.360 ;
        RECT 4.400 147.880 419.500 149.280 ;
        RECT 4.000 141.800 419.500 147.880 ;
        RECT 4.400 140.400 419.500 141.800 ;
        RECT 4.000 138.400 419.500 140.400 ;
        RECT 4.000 137.000 419.100 138.400 ;
        RECT 4.000 134.320 419.500 137.000 ;
        RECT 4.400 132.920 419.500 134.320 ;
        RECT 4.000 126.840 419.500 132.920 ;
        RECT 4.400 125.440 419.500 126.840 ;
        RECT 4.000 119.360 419.500 125.440 ;
        RECT 4.400 117.960 419.500 119.360 ;
        RECT 4.000 117.320 419.500 117.960 ;
        RECT 4.000 115.920 419.100 117.320 ;
        RECT 4.000 111.880 419.500 115.920 ;
        RECT 4.400 110.480 419.500 111.880 ;
        RECT 4.000 104.400 419.500 110.480 ;
        RECT 4.400 103.000 419.500 104.400 ;
        RECT 4.000 96.920 419.500 103.000 ;
        RECT 4.400 96.240 419.500 96.920 ;
        RECT 4.400 95.520 419.100 96.240 ;
        RECT 4.000 94.840 419.100 95.520 ;
        RECT 4.000 89.440 419.500 94.840 ;
        RECT 4.400 88.040 419.500 89.440 ;
        RECT 4.000 81.960 419.500 88.040 ;
        RECT 4.400 80.560 419.500 81.960 ;
        RECT 4.000 75.160 419.500 80.560 ;
        RECT 4.000 74.480 419.100 75.160 ;
        RECT 4.400 73.760 419.100 74.480 ;
        RECT 4.400 73.080 419.500 73.760 ;
        RECT 4.000 67.000 419.500 73.080 ;
        RECT 4.400 65.600 419.500 67.000 ;
        RECT 4.000 59.520 419.500 65.600 ;
        RECT 4.400 58.120 419.500 59.520 ;
        RECT 4.000 54.080 419.500 58.120 ;
        RECT 4.000 52.680 419.100 54.080 ;
        RECT 4.000 52.040 419.500 52.680 ;
        RECT 4.400 50.640 419.500 52.040 ;
        RECT 4.000 44.560 419.500 50.640 ;
        RECT 4.400 43.160 419.500 44.560 ;
        RECT 4.000 37.080 419.500 43.160 ;
        RECT 4.400 35.680 419.500 37.080 ;
        RECT 4.000 33.000 419.500 35.680 ;
        RECT 4.000 31.600 419.100 33.000 ;
        RECT 4.000 29.600 419.500 31.600 ;
        RECT 4.400 28.200 419.500 29.600 ;
        RECT 4.000 22.120 419.500 28.200 ;
        RECT 4.400 20.720 419.500 22.120 ;
        RECT 4.000 14.640 419.500 20.720 ;
        RECT 4.400 13.240 419.500 14.640 ;
        RECT 4.000 11.920 419.500 13.240 ;
        RECT 4.000 10.520 419.100 11.920 ;
        RECT 4.000 10.000 419.500 10.520 ;
        RECT 257.140 288.760 258.870 296.420 ;
        RECT 257.150 70.140 258.880 77.800 ;
      LAYER met4 ;
        RECT 31.575 10.000 40.320 390.840 ;
        RECT 42.720 10.000 43.620 390.840 ;
        RECT 46.020 10.000 64.320 390.840 ;
        RECT 66.720 225.445 67.620 390.840 ;
        RECT 70.020 266.930 398.850 390.840 ;
        RECT 70.020 225.445 88.320 266.930 ;
        RECT 90.720 225.445 91.620 266.930 ;
        RECT 94.020 225.445 112.320 266.930 ;
        RECT 114.720 225.445 115.620 266.930 ;
        RECT 118.020 225.445 136.320 266.930 ;
        RECT 66.720 176.515 136.320 225.445 ;
        RECT 66.720 10.000 67.620 176.515 ;
        RECT 70.020 133.910 88.320 176.515 ;
        RECT 90.720 133.910 91.620 176.515 ;
        RECT 94.020 133.910 112.320 176.515 ;
        RECT 114.720 133.910 115.620 176.515 ;
        RECT 118.020 133.910 136.320 176.515 ;
        RECT 138.720 133.910 139.620 266.930 ;
        RECT 142.020 133.910 160.320 266.930 ;
        RECT 162.720 133.910 163.620 266.930 ;
        RECT 166.020 133.910 184.320 266.930 ;
        RECT 186.720 229.260 187.620 266.930 ;
        RECT 190.020 229.260 208.320 266.930 ;
        RECT 186.720 166.580 208.320 229.260 ;
        RECT 186.720 133.910 187.620 166.580 ;
        RECT 190.020 133.910 208.320 166.580 ;
        RECT 210.720 229.260 211.620 266.930 ;
        RECT 214.020 229.260 232.320 266.930 ;
        RECT 210.720 166.580 232.320 229.260 ;
        RECT 210.720 133.910 211.620 166.580 ;
        RECT 214.020 133.910 232.320 166.580 ;
        RECT 234.720 133.910 235.620 266.930 ;
        RECT 238.020 215.790 256.320 266.930 ;
        RECT 258.720 215.790 259.620 266.930 ;
        RECT 262.020 215.790 280.320 266.930 ;
        RECT 238.020 182.140 280.320 215.790 ;
        RECT 238.020 133.910 256.320 182.140 ;
        RECT 258.720 133.910 259.620 182.140 ;
        RECT 262.020 133.910 280.320 182.140 ;
        RECT 282.720 133.910 283.620 266.930 ;
        RECT 286.020 226.100 398.850 266.930 ;
        RECT 286.020 196.560 304.320 226.100 ;
        RECT 306.720 196.560 307.620 226.100 ;
        RECT 310.020 196.560 328.320 226.100 ;
        RECT 330.720 196.560 331.620 226.100 ;
        RECT 334.020 196.560 352.320 226.100 ;
        RECT 354.720 196.560 355.620 226.100 ;
        RECT 358.020 204.870 398.850 226.100 ;
        RECT 358.020 196.560 376.320 204.870 ;
        RECT 286.020 173.900 376.320 196.560 ;
        RECT 378.720 173.900 398.850 204.870 ;
        RECT 286.020 133.910 398.850 173.900 ;
        RECT 70.020 10.000 398.850 133.910 ;
        RECT 257.140 288.760 258.870 296.420 ;
        RECT 257.150 70.140 258.880 77.800 ;
      LAYER met5 ;
        RECT 85.400 256.580 245.960 364.890 ;
        RECT 85.400 232.580 245.960 248.480 ;
        RECT 85.400 208.580 245.960 224.480 ;
        RECT 85.400 184.580 245.960 200.480 ;
        RECT 85.400 160.580 245.960 176.480 ;
        RECT 85.400 136.580 245.960 152.480 ;
        RECT 85.400 35.950 245.960 131.780 ;
        RECT 256.820 70.000 289.350 78.110 ;
        RECT 256.860 288.500 289.390 296.610 ;
  END
END adc_top
END LIBRARY

