* SPICE3 file created from Extract.ext - technology: sky130A

C0 cbot_4 ctop_4 30.99fF
C1 cbot_dummy cbot_8 14.65fF
C2 cbot_4 cbot_dummy 16.03fF
C3 cbot_2 ctop_2 29.86fF
C4 cbot_dummy cbot_1 15.99fF
C5 cbot_dummy cbot_2 16.01fF
C6 cbot_dummy ctop_dummy 247.72fF
C7 ctop_8 cbot_8 28.51fF
C8 ctop_1 cbot_1 29.29fF
C9 cbot_dummy VSUBS 43.58fF
