magic
tech sky130A
magscale 1 2
timestamp 1670857138
<< nwell >>
rect -38 414 2246 582
rect -38 247 822 414
rect 1556 247 2246 414
<< pwell >>
rect 822 214 1556 414
rect 1 -17 2207 214
<< scnmos >>
rect 113 80 851 164
rect 1021 71 1430 346
rect 1602 71 1632 155
rect 1698 71 1728 155
rect 1907 71 1937 155
rect 2003 71 2033 155
<< scpmoshvt >>
rect 285 283 569 443
rect 1661 329 1691 489
rect 1757 329 1787 489
rect 1995 329 2025 489
rect 2091 329 2121 489
<< ndiff >>
rect 963 334 1021 346
rect 55 127 113 164
rect 55 92 67 127
rect 101 92 113 127
rect 55 80 113 92
rect 851 144 909 164
rect 851 92 863 144
rect 897 92 909 144
rect 851 80 909 92
rect 963 79 975 334
rect 1009 79 1021 334
rect 963 71 1021 79
rect 1430 334 1488 346
rect 1430 79 1442 334
rect 1476 79 1488 334
rect 1430 71 1488 79
rect 1542 143 1602 155
rect 1542 83 1552 143
rect 1586 83 1602 143
rect 1542 71 1602 83
rect 1632 143 1698 155
rect 1632 85 1648 143
rect 1682 85 1698 143
rect 1632 71 1698 85
rect 1728 143 1786 155
rect 1728 85 1744 143
rect 1778 85 1786 143
rect 1728 71 1786 85
rect 1845 124 1907 155
rect 1845 85 1857 124
rect 1891 85 1907 124
rect 1845 71 1907 85
rect 1937 143 2003 155
rect 1937 85 1953 143
rect 1987 85 2003 143
rect 1937 71 2003 85
rect 2033 143 2095 155
rect 2033 85 2049 143
rect 2083 85 2095 143
rect 2033 71 2095 85
<< pdiff >>
rect 1601 477 1661 489
rect 227 431 285 443
rect 227 379 239 431
rect 273 379 285 431
rect 227 283 285 379
rect 569 431 627 443
rect 569 305 581 431
rect 615 305 627 431
rect 569 283 627 305
rect 1601 341 1611 477
rect 1645 341 1661 477
rect 1601 329 1661 341
rect 1691 475 1757 489
rect 1691 354 1707 475
rect 1741 354 1757 475
rect 1691 329 1757 354
rect 1787 475 1847 489
rect 1787 341 1803 475
rect 1837 341 1847 475
rect 1787 329 1847 341
rect 1933 475 1995 489
rect 1933 400 1945 475
rect 1979 400 1995 475
rect 1933 329 1995 400
rect 2025 475 2091 489
rect 2025 341 2041 475
rect 2075 341 2091 475
rect 2025 329 2091 341
rect 2121 475 2181 489
rect 2121 341 2137 475
rect 2171 341 2181 475
rect 2121 329 2181 341
<< ndiffc >>
rect 67 92 101 127
rect 863 92 897 144
rect 975 79 1009 334
rect 1442 79 1476 334
rect 1552 83 1586 143
rect 1648 85 1682 143
rect 1744 85 1778 143
rect 1857 85 1891 124
rect 1953 85 1987 143
rect 2049 85 2083 143
<< pdiffc >>
rect 239 379 273 431
rect 581 305 615 431
rect 1611 341 1645 477
rect 1707 354 1741 475
rect 1803 341 1837 475
rect 1945 400 1979 475
rect 2041 341 2075 475
rect 2137 341 2171 475
<< poly >>
rect 1661 489 1691 515
rect 1757 489 1787 515
rect 1995 489 2025 515
rect 2091 489 2121 515
rect 285 443 569 479
rect 650 428 1430 438
rect 649 418 1430 428
rect 649 384 1112 418
rect 1291 384 1430 418
rect 649 361 1430 384
rect 113 263 181 281
rect 113 225 126 263
rect 167 228 181 263
rect 285 228 569 283
rect 649 235 943 361
rect 1021 346 1430 361
rect 167 225 569 228
rect 113 190 569 225
rect 113 164 851 190
rect 113 54 851 80
rect 1661 314 1691 329
rect 1757 314 1787 329
rect 1661 284 1787 314
rect 1995 305 2025 329
rect 2091 305 2121 329
rect 1661 248 1691 284
rect 1602 236 1691 248
rect 1995 275 2121 305
rect 1995 265 2088 275
rect 1602 202 1641 236
rect 1675 214 1691 236
rect 1824 227 1890 238
rect 1675 202 1728 214
rect 1602 184 1728 202
rect 1602 155 1632 184
rect 1698 155 1728 184
rect 1824 193 1840 227
rect 1874 219 1890 227
rect 1995 231 2038 265
rect 2072 231 2088 265
rect 1995 219 2088 231
rect 1874 193 2033 219
rect 1824 189 2033 193
rect 1824 182 1937 189
rect 1907 155 1937 182
rect 2003 155 2033 189
rect 1021 32 1430 71
rect 1602 44 1632 71
rect 1698 44 1728 71
rect 1907 44 1937 71
rect 2003 44 2033 71
<< polycont >>
rect 1112 384 1291 418
rect 126 225 167 263
rect 1641 202 1675 236
rect 1840 193 1874 227
rect 2038 231 2072 265
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 1611 477 1645 527
rect 239 431 273 447
rect 238 379 239 400
rect 238 361 273 379
rect 581 431 615 447
rect 581 289 615 305
rect 650 336 1016 460
rect 1095 418 1407 425
rect 1095 384 1112 418
rect 1291 384 1407 418
rect 1095 374 1407 384
rect 1442 336 1476 351
rect 650 334 1476 336
rect 113 264 181 281
rect 21 263 181 264
rect 21 225 126 263
rect 167 225 181 263
rect 21 209 181 225
rect 21 198 75 209
rect 113 195 181 209
rect 650 196 975 334
rect 863 144 897 160
rect 67 127 101 143
rect 67 76 101 92
rect 863 58 897 92
rect 973 79 975 196
rect 1009 79 1442 334
rect 1611 325 1645 341
rect 1707 475 1741 491
rect 1707 325 1741 354
rect 1803 475 1837 491
rect 1542 268 1576 279
rect 1542 235 1586 268
rect 973 17 1476 79
rect 1552 143 1586 235
rect 1620 202 1631 236
rect 1675 202 1691 236
rect 1803 228 1837 341
rect 1871 296 1905 527
rect 1939 475 1979 491
rect 1939 400 1945 475
rect 1939 383 1979 400
rect 2041 475 2075 491
rect 2041 309 2075 341
rect 2137 475 2177 491
rect 2171 341 2177 475
rect 2137 325 2177 341
rect 1871 262 1987 296
rect 1803 227 1890 228
rect 1803 210 1840 227
rect 1744 193 1840 210
rect 1874 193 1890 227
rect 1744 176 1837 193
rect 1552 17 1586 83
rect 1648 143 1682 159
rect 1648 69 1682 85
rect 1744 143 1778 176
rect 1953 143 1987 262
rect 2022 231 2038 265
rect 2072 231 2089 265
rect 2043 193 2089 231
rect 1744 69 1778 85
rect 1857 133 1891 143
rect 1857 69 1891 85
rect 1953 69 1987 85
rect 2049 143 2083 159
rect 2049 69 2083 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 239 379 273 431
rect 581 305 615 417
rect 1136 384 1172 418
rect 1234 384 1270 418
rect 67 92 101 127
rect 863 92 897 128
rect 1707 354 1741 445
rect 1542 279 1576 313
rect 1631 202 1641 236
rect 1641 202 1675 236
rect 1945 412 1979 451
rect 2041 341 2075 389
rect 2137 361 2171 443
rect 1648 105 1682 143
rect 1857 124 1891 133
rect 1857 99 1891 124
rect 2049 105 2083 139
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 233 431 279 496
rect 233 379 239 431
rect 273 379 279 431
rect 233 362 279 379
rect 573 417 1016 460
rect 1701 451 2177 458
rect 1701 445 1945 451
rect 238 361 273 362
rect 573 305 581 417
rect 615 336 1016 417
rect 1124 418 1282 424
rect 1124 384 1136 418
rect 1172 384 1234 418
rect 1270 384 1282 418
rect 1124 378 1282 384
rect 1181 336 1226 378
rect 1701 354 1707 445
rect 1741 430 1945 445
rect 1741 354 1747 430
rect 1939 412 1945 430
rect 1979 443 2177 451
rect 1979 430 2137 443
rect 1979 412 1985 430
rect 1939 400 1985 412
rect 1701 342 1747 354
rect 2035 389 2081 402
rect 2035 341 2041 389
rect 2075 341 2081 389
rect 2131 361 2137 430
rect 2171 361 2177 443
rect 2131 349 2177 361
rect 615 305 1496 336
rect 573 223 1496 305
rect 1530 314 1582 320
rect 2035 314 2081 341
rect 1530 313 2081 314
rect 1530 279 1542 313
rect 1576 279 2081 313
rect 1530 275 2081 279
rect 1530 273 1582 275
rect 1601 236 1691 242
rect 1601 223 1631 236
rect 573 202 1631 223
rect 1675 202 1691 236
rect 573 196 1691 202
rect 955 184 1691 196
rect 955 142 1496 184
rect 61 127 107 140
rect 61 92 67 127
rect 101 92 107 127
rect 61 48 107 92
rect 856 128 1496 142
rect 856 92 863 128
rect 897 93 1496 128
rect 1642 143 1688 155
rect 1642 105 1648 143
rect 1682 121 1688 143
rect 2037 139 2095 147
rect 1845 133 1903 139
rect 1845 121 1857 133
rect 1682 105 1857 121
rect 1642 99 1857 105
rect 1891 121 1903 133
rect 2037 121 2049 139
rect 1891 105 2049 121
rect 2083 113 2095 139
rect 2083 105 2089 113
rect 1891 99 2089 105
rect 1642 93 2089 99
rect 897 92 940 93
rect 856 78 940 92
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel metal1 s 0 496 2208 592 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -48 2208 48 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 673 527 707 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel metal1 s 673 -17 707 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 673 527 707 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 673 -17 707 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 121 -17 155 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 121 527 155 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 121 527 155 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 121 -17 155 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 1225 -17 1259 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 1225 -17 1259 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel locali s 40 221 74 255 7 FreeSans 160 0 0 0 in
port 2 nsew signal input
rlabel metal1 982 285 982 285 1 mid
flabel pwell s 1777 -17 1811 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 1777 -17 1811 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 1409 527 1443 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 1409 527 1443 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 1869 527 1903 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 1869 527 1903 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 2053 527 2087 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 2053 527 2087 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel locali s 2049 207 2083 241 0 FreeSans 160 0 0 0 out
port 3 nsew signal output
flabel metal1 s 1317 -17 1351 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 1317 -17 1351 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 949 -17 983 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 949 -17 983 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
string LEFsource USER
<< end >>
