* SPICE3 file created from adc_array_cap_16.ext - technology: sky130A

.subckt adc_array_circuit SAMPLE_N SAMPLE COLON_N COL_N ROW_N VCOM CBOT VINT VINT2
+ VDRV VDD VSS
X0 VINT2 COLON_N VDRV VSS sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.86e+06u as=2.52e+11p ps=2.88e+06u w=420000u l=180000u
X1 VINT2 ROW_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.26e+11p ps=1.44e+06u w=420000u l=180000u
X2 VSS COL_N VINT2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X3 CBOT SAMPLE_N VCOM VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=4.5e+11p ps=2.8e+06u w=900000u l=180000u
X4 VDRV SAMPLE CBOT VDD sky130_fd_pr__pfet_01v8 ad=1.305e+12p pd=8.3e+06u as=0p ps=0u w=900000u l=180000u
X5 VINT COL_N VDRV VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=0p ps=0u w=900000u l=180000u
X6 CBOT SAMPLE_N VDRV VSS sky130_fd_pr__nfet_01v8 ad=1.26e+11p pd=1.44e+06u as=0p ps=0u w=420000u l=180000u
X7 VCOM SAMPLE CBOT VSS sky130_fd_pr__nfet_01v8 ad=1.26e+11p pd=1.44e+06u as=0p ps=0u w=420000u l=180000u
X8 VDD ROW_N VINT VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=0p ps=0u w=900000u l=180000u
X9 VDRV COLON_N VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=180000u
C0 COLON_N COL_N 1.23fF
C1 VDRV COL_N 0.98fF
C2 SAMPLE_N VDD 1.16fF
C3 COLON_N SAMPLE 0.69fF
C4 VCOM VSS 1.65fF
C5 ROW_N VSS 1.02fF
C6 VDD VSS 2.65fF
.ends

.subckt adc_array_cap_16 COL_N COLON_N CTOP ROW_N SAMPLE SAMPLE_N VCOM VDD CBOT VSS
Xadc_array_circuit_0 SAMPLE_N SAMPLE COLON_N COL_N ROW_N VCOM CBOT adc_array_circuit_0/VINT
+ adc_array_circuit_0/VINT2 adc_array_circuit_0/VDRV VDD VSS adc_array_circuit
C0 CBOT adc_array_circuit_0/VDRV 0.42fF
C1 VCOM CBOT 0.47fF
C2 VDD CBOT 0.91fF
C3 CTOP CBOT 7.87fF
C4 CTOP VSS 0.91fF
C5 CBOT VSS 2.82fF
C6 VCOM VSS 1.65fF
C7 ROW_N VSS 1.02fF
C8 VDD VSS 2.65fF
.ends

