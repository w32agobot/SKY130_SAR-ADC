magic
tech sky130A
magscale 1 2
timestamp 1663078155
<< nwell >>
rect -53 -53 3939 3873
<< pmos >>
rect 143 95 3743 3683
<< pdiff >>
rect 85 3647 143 3683
rect 85 107 97 3647
rect 131 107 143 3647
rect 85 95 143 107
rect 3743 3647 3801 3683
rect 3743 107 3755 3647
rect 3789 107 3801 3647
rect 3743 95 3801 107
<< pdiffc >>
rect 97 107 131 3647
rect 3755 107 3789 3647
<< nsubdiff >>
rect -17 3803 79 3837
rect 3807 3803 3903 3837
rect -17 3741 17 3803
rect 3869 3741 3903 3803
rect -17 17 17 79
rect 3869 17 3903 79
rect -17 -17 79 17
rect 3807 -17 3903 17
<< nsubdiffcont >>
rect 79 3803 3807 3837
rect -17 79 17 3741
rect 3869 79 3903 3741
rect 79 -17 3807 17
<< poly >>
rect 143 3764 3743 3777
rect 143 3730 182 3764
rect 220 3730 262 3764
rect 300 3730 342 3764
rect 380 3730 422 3764
rect 460 3730 502 3764
rect 540 3730 582 3764
rect 620 3730 662 3764
rect 700 3730 742 3764
rect 780 3730 822 3764
rect 860 3730 902 3764
rect 940 3730 982 3764
rect 1020 3730 1062 3764
rect 1100 3730 1142 3764
rect 1180 3730 1222 3764
rect 1260 3730 1302 3764
rect 1340 3730 1382 3764
rect 1420 3730 1462 3764
rect 1500 3730 1542 3764
rect 1580 3730 1622 3764
rect 1660 3730 1702 3764
rect 1740 3730 1782 3764
rect 1820 3730 1862 3764
rect 1900 3730 1942 3764
rect 1980 3730 2022 3764
rect 2060 3730 2102 3764
rect 2140 3730 2182 3764
rect 2220 3730 2262 3764
rect 2300 3730 2342 3764
rect 2380 3730 2422 3764
rect 2460 3730 2502 3764
rect 2540 3730 2582 3764
rect 2620 3730 2662 3764
rect 2700 3730 2742 3764
rect 2780 3730 2822 3764
rect 2860 3730 2902 3764
rect 2940 3730 2982 3764
rect 3020 3730 3062 3764
rect 3100 3730 3142 3764
rect 3180 3730 3222 3764
rect 3260 3730 3302 3764
rect 3340 3730 3382 3764
rect 3420 3730 3462 3764
rect 3500 3730 3542 3764
rect 3580 3730 3622 3764
rect 3660 3730 3743 3764
rect 143 3683 3743 3730
rect 143 69 3743 95
<< polycont >>
rect 182 3730 220 3764
rect 262 3730 300 3764
rect 342 3730 380 3764
rect 422 3730 460 3764
rect 502 3730 540 3764
rect 582 3730 620 3764
rect 662 3730 700 3764
rect 742 3730 780 3764
rect 822 3730 860 3764
rect 902 3730 940 3764
rect 982 3730 1020 3764
rect 1062 3730 1100 3764
rect 1142 3730 1180 3764
rect 1222 3730 1260 3764
rect 1302 3730 1340 3764
rect 1382 3730 1420 3764
rect 1462 3730 1500 3764
rect 1542 3730 1580 3764
rect 1622 3730 1660 3764
rect 1702 3730 1740 3764
rect 1782 3730 1820 3764
rect 1862 3730 1900 3764
rect 1942 3730 1980 3764
rect 2022 3730 2060 3764
rect 2102 3730 2140 3764
rect 2182 3730 2220 3764
rect 2262 3730 2300 3764
rect 2342 3730 2380 3764
rect 2422 3730 2460 3764
rect 2502 3730 2540 3764
rect 2582 3730 2620 3764
rect 2662 3730 2700 3764
rect 2742 3730 2780 3764
rect 2822 3730 2860 3764
rect 2902 3730 2940 3764
rect 2982 3730 3020 3764
rect 3062 3730 3100 3764
rect 3142 3730 3180 3764
rect 3222 3730 3260 3764
rect 3302 3730 3340 3764
rect 3382 3730 3420 3764
rect 3462 3730 3500 3764
rect 3542 3730 3580 3764
rect 3622 3730 3660 3764
<< locali >>
rect 63 3803 79 3837
rect 3807 3803 3823 3837
rect -17 3741 17 3757
rect 166 3730 182 3764
rect 220 3730 262 3764
rect 300 3730 342 3764
rect 380 3730 422 3764
rect 460 3730 502 3764
rect 540 3730 582 3764
rect 620 3730 662 3764
rect 700 3730 742 3764
rect 780 3730 822 3764
rect 860 3730 902 3764
rect 940 3730 982 3764
rect 1020 3730 1062 3764
rect 1100 3730 1142 3764
rect 1180 3730 1222 3764
rect 1260 3730 1302 3764
rect 1340 3730 1382 3764
rect 1420 3730 1462 3764
rect 1500 3730 1542 3764
rect 1580 3730 1622 3764
rect 1660 3730 1702 3764
rect 1740 3730 1782 3764
rect 1820 3730 1862 3764
rect 1900 3730 1942 3764
rect 1980 3730 2022 3764
rect 2060 3730 2102 3764
rect 2140 3730 2182 3764
rect 2220 3730 2262 3764
rect 2300 3730 2342 3764
rect 2380 3730 2422 3764
rect 2460 3730 2502 3764
rect 2540 3730 2582 3764
rect 2620 3730 2662 3764
rect 2700 3730 2742 3764
rect 2780 3730 2822 3764
rect 2860 3730 2902 3764
rect 2940 3730 2982 3764
rect 3020 3730 3062 3764
rect 3100 3730 3142 3764
rect 3180 3730 3222 3764
rect 3260 3730 3302 3764
rect 3340 3730 3382 3764
rect 3420 3730 3462 3764
rect 3500 3730 3542 3764
rect 3580 3730 3622 3764
rect 3660 3730 3694 3764
rect 3869 3741 3903 3757
rect 97 3647 131 3687
rect 97 91 131 107
rect 3755 3647 3789 3687
rect 3755 91 3789 107
rect -17 63 17 79
rect 3869 63 3903 79
rect 63 -17 79 17
rect 3807 -17 3823 17
<< viali >>
rect 182 3730 220 3764
rect 262 3730 300 3764
rect 342 3730 380 3764
rect 422 3730 460 3764
rect 502 3730 540 3764
rect 582 3730 620 3764
rect 662 3730 700 3764
rect 742 3730 780 3764
rect 822 3730 860 3764
rect 902 3730 940 3764
rect 982 3730 1020 3764
rect 1062 3730 1100 3764
rect 1142 3730 1180 3764
rect 1222 3730 1260 3764
rect 1302 3730 1340 3764
rect 1382 3730 1420 3764
rect 1462 3730 1500 3764
rect 1542 3730 1580 3764
rect 1622 3730 1660 3764
rect 1702 3730 1740 3764
rect 1782 3730 1820 3764
rect 1862 3730 1900 3764
rect 1942 3730 1980 3764
rect 2022 3730 2060 3764
rect 2102 3730 2140 3764
rect 2182 3730 2220 3764
rect 2262 3730 2300 3764
rect 2342 3730 2380 3764
rect 2422 3730 2460 3764
rect 2502 3730 2540 3764
rect 2582 3730 2620 3764
rect 2662 3730 2700 3764
rect 2742 3730 2780 3764
rect 2822 3730 2860 3764
rect 2902 3730 2940 3764
rect 2982 3730 3020 3764
rect 3062 3730 3100 3764
rect 3142 3730 3180 3764
rect 3222 3730 3260 3764
rect 3302 3730 3340 3764
rect 3382 3730 3420 3764
rect 3462 3730 3500 3764
rect 3542 3730 3580 3764
rect 3622 3730 3660 3764
rect 97 107 131 3647
rect 3755 107 3789 3647
<< metal1 >>
rect 168 3722 174 3774
rect 226 3722 254 3774
rect 306 3722 334 3774
rect 386 3722 414 3774
rect 466 3722 494 3774
rect 546 3722 574 3774
rect 626 3722 654 3774
rect 706 3722 734 3774
rect 786 3722 814 3774
rect 866 3722 894 3774
rect 946 3722 974 3774
rect 1026 3722 1054 3774
rect 1106 3722 1134 3774
rect 1186 3722 1214 3774
rect 1266 3722 1294 3774
rect 1346 3722 1374 3774
rect 1426 3722 1454 3774
rect 1506 3722 1534 3774
rect 1586 3722 1614 3774
rect 1666 3722 1694 3774
rect 1746 3722 1774 3774
rect 1826 3722 1854 3774
rect 1906 3722 1934 3774
rect 1986 3722 2014 3774
rect 2066 3722 2094 3774
rect 2146 3722 2174 3774
rect 2226 3722 2254 3774
rect 2306 3722 2334 3774
rect 2386 3722 2414 3774
rect 2466 3722 2494 3774
rect 2546 3722 2574 3774
rect 2626 3722 2654 3774
rect 2706 3722 2734 3774
rect 2786 3722 2814 3774
rect 2866 3722 2894 3774
rect 2946 3722 2974 3774
rect 3026 3722 3054 3774
rect 3106 3722 3134 3774
rect 3186 3722 3214 3774
rect 3266 3722 3294 3774
rect 3346 3722 3374 3774
rect 3426 3722 3454 3774
rect 3506 3722 3534 3774
rect 3586 3722 3614 3774
rect 3666 3722 3694 3774
rect 90 3647 3796 3662
rect 90 107 97 3647
rect 131 107 3755 3647
rect 3789 107 3796 3647
rect 90 94 3796 107
<< via1 >>
rect 174 3764 226 3774
rect 174 3730 182 3764
rect 182 3730 220 3764
rect 220 3730 226 3764
rect 174 3722 226 3730
rect 254 3764 306 3774
rect 254 3730 262 3764
rect 262 3730 300 3764
rect 300 3730 306 3764
rect 254 3722 306 3730
rect 334 3764 386 3774
rect 334 3730 342 3764
rect 342 3730 380 3764
rect 380 3730 386 3764
rect 334 3722 386 3730
rect 414 3764 466 3774
rect 414 3730 422 3764
rect 422 3730 460 3764
rect 460 3730 466 3764
rect 414 3722 466 3730
rect 494 3764 546 3774
rect 494 3730 502 3764
rect 502 3730 540 3764
rect 540 3730 546 3764
rect 494 3722 546 3730
rect 574 3764 626 3774
rect 574 3730 582 3764
rect 582 3730 620 3764
rect 620 3730 626 3764
rect 574 3722 626 3730
rect 654 3764 706 3774
rect 654 3730 662 3764
rect 662 3730 700 3764
rect 700 3730 706 3764
rect 654 3722 706 3730
rect 734 3764 786 3774
rect 734 3730 742 3764
rect 742 3730 780 3764
rect 780 3730 786 3764
rect 734 3722 786 3730
rect 814 3764 866 3774
rect 814 3730 822 3764
rect 822 3730 860 3764
rect 860 3730 866 3764
rect 814 3722 866 3730
rect 894 3764 946 3774
rect 894 3730 902 3764
rect 902 3730 940 3764
rect 940 3730 946 3764
rect 894 3722 946 3730
rect 974 3764 1026 3774
rect 974 3730 982 3764
rect 982 3730 1020 3764
rect 1020 3730 1026 3764
rect 974 3722 1026 3730
rect 1054 3764 1106 3774
rect 1054 3730 1062 3764
rect 1062 3730 1100 3764
rect 1100 3730 1106 3764
rect 1054 3722 1106 3730
rect 1134 3764 1186 3774
rect 1134 3730 1142 3764
rect 1142 3730 1180 3764
rect 1180 3730 1186 3764
rect 1134 3722 1186 3730
rect 1214 3764 1266 3774
rect 1214 3730 1222 3764
rect 1222 3730 1260 3764
rect 1260 3730 1266 3764
rect 1214 3722 1266 3730
rect 1294 3764 1346 3774
rect 1294 3730 1302 3764
rect 1302 3730 1340 3764
rect 1340 3730 1346 3764
rect 1294 3722 1346 3730
rect 1374 3764 1426 3774
rect 1374 3730 1382 3764
rect 1382 3730 1420 3764
rect 1420 3730 1426 3764
rect 1374 3722 1426 3730
rect 1454 3764 1506 3774
rect 1454 3730 1462 3764
rect 1462 3730 1500 3764
rect 1500 3730 1506 3764
rect 1454 3722 1506 3730
rect 1534 3764 1586 3774
rect 1534 3730 1542 3764
rect 1542 3730 1580 3764
rect 1580 3730 1586 3764
rect 1534 3722 1586 3730
rect 1614 3764 1666 3774
rect 1614 3730 1622 3764
rect 1622 3730 1660 3764
rect 1660 3730 1666 3764
rect 1614 3722 1666 3730
rect 1694 3764 1746 3774
rect 1694 3730 1702 3764
rect 1702 3730 1740 3764
rect 1740 3730 1746 3764
rect 1694 3722 1746 3730
rect 1774 3764 1826 3774
rect 1774 3730 1782 3764
rect 1782 3730 1820 3764
rect 1820 3730 1826 3764
rect 1774 3722 1826 3730
rect 1854 3764 1906 3774
rect 1854 3730 1862 3764
rect 1862 3730 1900 3764
rect 1900 3730 1906 3764
rect 1854 3722 1906 3730
rect 1934 3764 1986 3774
rect 1934 3730 1942 3764
rect 1942 3730 1980 3764
rect 1980 3730 1986 3764
rect 1934 3722 1986 3730
rect 2014 3764 2066 3774
rect 2014 3730 2022 3764
rect 2022 3730 2060 3764
rect 2060 3730 2066 3764
rect 2014 3722 2066 3730
rect 2094 3764 2146 3774
rect 2094 3730 2102 3764
rect 2102 3730 2140 3764
rect 2140 3730 2146 3764
rect 2094 3722 2146 3730
rect 2174 3764 2226 3774
rect 2174 3730 2182 3764
rect 2182 3730 2220 3764
rect 2220 3730 2226 3764
rect 2174 3722 2226 3730
rect 2254 3764 2306 3774
rect 2254 3730 2262 3764
rect 2262 3730 2300 3764
rect 2300 3730 2306 3764
rect 2254 3722 2306 3730
rect 2334 3764 2386 3774
rect 2334 3730 2342 3764
rect 2342 3730 2380 3764
rect 2380 3730 2386 3764
rect 2334 3722 2386 3730
rect 2414 3764 2466 3774
rect 2414 3730 2422 3764
rect 2422 3730 2460 3764
rect 2460 3730 2466 3764
rect 2414 3722 2466 3730
rect 2494 3764 2546 3774
rect 2494 3730 2502 3764
rect 2502 3730 2540 3764
rect 2540 3730 2546 3764
rect 2494 3722 2546 3730
rect 2574 3764 2626 3774
rect 2574 3730 2582 3764
rect 2582 3730 2620 3764
rect 2620 3730 2626 3764
rect 2574 3722 2626 3730
rect 2654 3764 2706 3774
rect 2654 3730 2662 3764
rect 2662 3730 2700 3764
rect 2700 3730 2706 3764
rect 2654 3722 2706 3730
rect 2734 3764 2786 3774
rect 2734 3730 2742 3764
rect 2742 3730 2780 3764
rect 2780 3730 2786 3764
rect 2734 3722 2786 3730
rect 2814 3764 2866 3774
rect 2814 3730 2822 3764
rect 2822 3730 2860 3764
rect 2860 3730 2866 3764
rect 2814 3722 2866 3730
rect 2894 3764 2946 3774
rect 2894 3730 2902 3764
rect 2902 3730 2940 3764
rect 2940 3730 2946 3764
rect 2894 3722 2946 3730
rect 2974 3764 3026 3774
rect 2974 3730 2982 3764
rect 2982 3730 3020 3764
rect 3020 3730 3026 3764
rect 2974 3722 3026 3730
rect 3054 3764 3106 3774
rect 3054 3730 3062 3764
rect 3062 3730 3100 3764
rect 3100 3730 3106 3764
rect 3054 3722 3106 3730
rect 3134 3764 3186 3774
rect 3134 3730 3142 3764
rect 3142 3730 3180 3764
rect 3180 3730 3186 3764
rect 3134 3722 3186 3730
rect 3214 3764 3266 3774
rect 3214 3730 3222 3764
rect 3222 3730 3260 3764
rect 3260 3730 3266 3764
rect 3214 3722 3266 3730
rect 3294 3764 3346 3774
rect 3294 3730 3302 3764
rect 3302 3730 3340 3764
rect 3340 3730 3346 3764
rect 3294 3722 3346 3730
rect 3374 3764 3426 3774
rect 3374 3730 3382 3764
rect 3382 3730 3420 3764
rect 3420 3730 3426 3764
rect 3374 3722 3426 3730
rect 3454 3764 3506 3774
rect 3454 3730 3462 3764
rect 3462 3730 3500 3764
rect 3500 3730 3506 3764
rect 3454 3722 3506 3730
rect 3534 3764 3586 3774
rect 3534 3730 3542 3764
rect 3542 3730 3580 3764
rect 3580 3730 3586 3764
rect 3534 3722 3586 3730
rect 3614 3764 3666 3774
rect 3614 3730 3622 3764
rect 3622 3730 3660 3764
rect 3660 3730 3666 3764
rect 3614 3722 3666 3730
<< metal2 >>
rect 168 3722 174 3774
rect 226 3722 254 3774
rect 306 3722 334 3774
rect 386 3722 414 3774
rect 466 3722 494 3774
rect 546 3722 574 3774
rect 626 3722 654 3774
rect 706 3722 734 3774
rect 786 3722 814 3774
rect 866 3722 894 3774
rect 946 3722 974 3774
rect 1026 3722 1054 3774
rect 1106 3722 1134 3774
rect 1186 3722 1214 3774
rect 1266 3722 1294 3774
rect 1346 3722 1374 3774
rect 1426 3722 1454 3774
rect 1506 3722 1534 3774
rect 1586 3722 1614 3774
rect 1666 3722 1694 3774
rect 1746 3722 1774 3774
rect 1826 3722 1854 3774
rect 1906 3722 1934 3774
rect 1986 3722 2014 3774
rect 2066 3722 2094 3774
rect 2146 3722 2174 3774
rect 2226 3722 2254 3774
rect 2306 3722 2334 3774
rect 2386 3722 2414 3774
rect 2466 3722 2494 3774
rect 2546 3722 2574 3774
rect 2626 3722 2654 3774
rect 2706 3722 2734 3774
rect 2786 3722 2814 3774
rect 2866 3722 2894 3774
rect 2946 3722 2974 3774
rect 3026 3722 3054 3774
rect 3106 3722 3134 3774
rect 3186 3722 3214 3774
rect 3266 3722 3294 3774
rect 3346 3722 3374 3774
rect 3426 3722 3454 3774
rect 3506 3722 3534 3774
rect 3586 3722 3614 3774
rect 3666 3722 3694 3774
rect 168 106 196 3722
rect 224 78 252 3688
rect 280 106 308 3722
rect 336 78 364 3688
rect 392 106 420 3722
rect 448 78 476 3688
rect 504 106 532 3722
rect 560 78 588 3688
rect 616 106 644 3722
rect 672 78 700 3688
rect 728 106 756 3722
rect 784 78 812 3688
rect 840 106 868 3722
rect 896 78 924 3688
rect 952 106 980 3722
rect 1008 78 1036 3688
rect 1064 106 1092 3722
rect 1120 78 1148 3688
rect 1176 106 1204 3722
rect 1232 78 1260 3688
rect 1288 106 1316 3722
rect 1344 78 1372 3688
rect 1400 106 1428 3722
rect 1456 78 1484 3688
rect 1512 106 1540 3722
rect 1568 78 1596 3688
rect 1624 106 1652 3722
rect 1680 78 1708 3688
rect 1736 106 1764 3722
rect 1792 78 1820 3688
rect 1848 106 1876 3722
rect 1904 78 1932 3688
rect 1960 106 1988 3722
rect 2016 78 2044 3688
rect 2072 106 2100 3722
rect 2128 78 2156 3688
rect 2184 106 2212 3722
rect 2240 78 2268 3688
rect 2296 106 2324 3722
rect 2352 78 2380 3688
rect 2408 106 2436 3722
rect 2464 78 2492 3688
rect 2520 106 2548 3722
rect 2576 78 2604 3688
rect 2632 106 2660 3722
rect 2688 78 2716 3688
rect 2744 106 2772 3722
rect 2800 78 2828 3688
rect 2856 106 2884 3722
rect 2912 78 2940 3688
rect 2968 106 2996 3722
rect 3024 78 3052 3688
rect 3080 106 3108 3722
rect 3136 78 3164 3688
rect 3192 106 3220 3722
rect 3248 78 3276 3688
rect 3304 106 3332 3722
rect 3360 78 3388 3688
rect 3416 106 3444 3722
rect 3472 78 3500 3688
rect 3528 106 3556 3722
rect 3584 78 3612 3688
rect 3640 106 3668 3722
rect 3696 78 3724 3688
rect 168 50 3724 78
<< metal3 >>
rect 86 3668 3785 3696
rect 86 124 3701 3668
rect 3765 124 3785 3668
rect 86 96 3785 124
<< via3 >>
rect 3701 124 3765 3668
<< mimcap >>
rect 186 3556 3586 3596
rect 186 236 226 3556
rect 3546 236 3586 3556
rect 186 196 3586 236
<< mimcapcontact >>
rect 226 236 3546 3556
<< metal4 >>
rect 86 3668 4188 3696
rect 86 3556 3701 3668
rect 86 236 226 3556
rect 3546 236 3701 3556
rect 86 124 3701 236
rect 3765 3655 4188 3668
rect 3765 137 3932 3655
rect 4168 137 4188 3655
rect 3765 124 4188 137
rect 86 96 4188 124
<< via4 >>
rect 3932 137 4168 3655
<< mimcap2 >>
rect 186 3556 3586 3596
rect 186 236 226 3556
rect 3546 236 3586 3556
rect 186 196 3586 236
<< mimcap2contact >>
rect 226 236 3546 3556
<< metal5 >>
rect 3890 3655 4210 3697
rect 202 3556 3570 3580
rect 202 236 226 3556
rect 3546 236 3570 3556
rect 202 212 3570 236
rect 3890 137 3932 3655
rect 4168 137 4210 3655
rect 3890 95 4210 137
<< end >>
