VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO emptybox_50_35
  CLASS BLOCK ;
  FOREIGN emptybox_50_35 ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 35.000 ;
  OBS
      LAYER met1 ;
        RECT 0.120 0.100 49.500 34.710 ;
  END
END emptybox_50_35
END LIBRARY

