magic
tech sky130A
magscale 1 2
timestamp 1666972778
<< nwell >>
rect 2877 34830 2941 34831
rect 1279 34265 3154 34830
rect 1279 34264 1569 34265
rect 1629 33421 3020 33437
rect 1463 33177 3020 33421
rect 1463 33176 1925 33177
<< psubdiff >>
rect 944 35679 5204 35727
rect 944 35519 1306 35679
rect 1466 35519 1706 35679
rect 1866 35519 2106 35679
rect 2266 35519 2506 35679
rect 2666 35519 2906 35679
rect 3066 35519 3306 35679
rect 3466 35519 3706 35679
rect 3866 35519 4106 35679
rect 4266 35519 4506 35679
rect 4666 35519 5204 35679
rect 944 35496 5204 35519
rect 944 35336 1008 35496
rect 1168 35476 4983 35496
rect 1168 35336 1237 35476
rect 944 35096 1237 35336
rect 944 34936 1008 35096
rect 1168 34936 1237 35096
rect 4915 35336 4983 35476
rect 5143 35476 5204 35496
rect 5143 35336 5203 35476
rect 4915 35096 5203 35336
rect 944 34696 1237 34936
rect 4915 34936 4983 35096
rect 5143 34936 5203 35096
rect 944 34536 1008 34696
rect 1168 34536 1237 34696
rect 944 34296 1237 34536
rect 944 34136 1008 34296
rect 1168 34136 1237 34296
rect 944 33896 1237 34136
rect 944 33736 1008 33896
rect 1168 33736 1237 33896
rect 944 33496 1237 33736
rect 944 33336 1008 33496
rect 1168 33336 1237 33496
rect 944 33096 1237 33336
rect 4915 34696 5203 34936
rect 4915 34536 4983 34696
rect 5143 34536 5203 34696
rect 4915 34296 5203 34536
rect 4915 34136 4983 34296
rect 5143 34136 5203 34296
rect 4915 33896 5203 34136
rect 4915 33736 4983 33896
rect 5143 33736 5203 33896
rect 4915 33496 5203 33736
rect 4915 33336 4983 33496
rect 5143 33336 5203 33496
rect 944 32936 1008 33096
rect 1168 32936 1237 33096
rect 4915 33096 5203 33336
rect 944 32650 1237 32936
rect 4915 32936 4983 33096
rect 5143 32936 5203 33096
rect 4915 32732 5203 32936
rect 4915 32650 5204 32732
rect 944 32649 2538 32650
rect 2685 32649 5204 32650
rect 944 32614 5204 32649
rect 944 32454 1008 32614
rect 1168 32454 1408 32614
rect 1568 32454 1808 32614
rect 1968 32454 2208 32614
rect 2368 32609 3408 32614
rect 2368 32454 2742 32609
rect 944 32449 2742 32454
rect 2902 32449 3069 32609
rect 3229 32454 3408 32609
rect 3568 32454 3808 32614
rect 3968 32454 4208 32614
rect 4368 32454 4608 32614
rect 4768 32454 4983 32614
rect 5143 32454 5204 32614
rect 3229 32449 5204 32454
rect 944 32411 5203 32449
<< psubdiffcont >>
rect 1306 35519 1466 35679
rect 1706 35519 1866 35679
rect 2106 35519 2266 35679
rect 2506 35519 2666 35679
rect 2906 35519 3066 35679
rect 3306 35519 3466 35679
rect 3706 35519 3866 35679
rect 4106 35519 4266 35679
rect 4506 35519 4666 35679
rect 1008 35336 1168 35496
rect 1008 34936 1168 35096
rect 4983 35336 5143 35496
rect 4983 34936 5143 35096
rect 1008 34536 1168 34696
rect 1008 34136 1168 34296
rect 1008 33736 1168 33896
rect 1008 33336 1168 33496
rect 4983 34536 5143 34696
rect 4983 34136 5143 34296
rect 4983 33736 5143 33896
rect 4983 33336 5143 33496
rect 1008 32936 1168 33096
rect 4983 32936 5143 33096
rect 1008 32454 1168 32614
rect 1408 32454 1568 32614
rect 1808 32454 1968 32614
rect 2208 32454 2368 32614
rect 2742 32449 2902 32609
rect 3069 32449 3229 32609
rect 3408 32454 3568 32614
rect 3808 32454 3968 32614
rect 4208 32454 4368 32614
rect 4608 32454 4768 32614
rect 4983 32454 5143 32614
<< poly >>
rect 2885 34981 2951 34994
rect 2885 34966 2901 34981
rect 2039 34964 2901 34966
rect 1650 34947 2901 34964
rect 2935 34947 2951 34981
rect 1650 34934 2951 34947
rect 1650 34870 2965 34892
rect 1650 34862 2921 34870
rect 1650 34819 1750 34862
rect 1808 34819 1908 34862
rect 2081 34816 2181 34862
rect 2239 34817 2339 34862
rect 2526 34817 2626 34862
rect 2684 34817 2784 34862
rect 2911 34836 2921 34862
rect 2955 34836 2965 34870
rect 2911 34820 2965 34836
rect 2526 34816 2538 34817
rect 2003 33144 2103 33197
rect 2161 33144 2261 33198
rect 2483 33144 2583 33198
rect 2641 33144 2741 33197
rect 2944 33172 3012 33182
rect 2944 33144 2962 33172
rect 2003 33138 2962 33144
rect 2996 33138 3012 33172
rect 2003 33114 3012 33138
rect 2003 33040 2969 33070
rect 2900 33038 2969 33040
rect 2900 33003 2916 33038
rect 2953 33003 2969 33038
rect 2900 32992 2969 33003
<< polycont >>
rect 2901 34947 2935 34981
rect 2921 34836 2955 34870
rect 2962 33138 2996 33172
rect 2916 33003 2953 33038
<< locali >>
rect 463 67060 946 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 946 67060
rect 463 66913 946 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 946 66913
rect 463 66776 946 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 946 66776
rect 463 66650 946 66700
rect 463 65300 946 65349
rect 463 65224 504 65300
rect 576 65224 626 65300
rect 698 65224 752 65300
rect 824 65224 946 65300
rect 463 65153 946 65224
rect 463 65077 504 65153
rect 576 65077 626 65153
rect 698 65077 752 65153
rect 824 65077 946 65153
rect 463 65016 946 65077
rect 463 64940 504 65016
rect 576 64940 626 65016
rect 698 64940 752 65016
rect 824 64940 946 65016
rect 463 64890 946 64940
rect 463 63060 946 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 946 63060
rect 463 62913 946 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 946 62913
rect 463 62776 946 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 946 62776
rect 463 62650 946 62700
rect 463 61301 946 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 946 61301
rect 463 61154 946 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 946 61154
rect 463 61017 946 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 946 61017
rect 463 60891 946 60941
rect 464 59068 947 59109
rect 463 59060 947 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 947 59060
rect 463 58913 947 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 947 58913
rect 463 58776 947 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 947 58776
rect 463 58650 947 58700
rect 463 57301 946 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 946 57301
rect 463 57154 946 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 946 57154
rect 463 57017 946 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 946 57017
rect 463 56891 946 56941
rect 464 55068 947 55109
rect 463 55060 947 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 947 55060
rect 463 54913 947 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 947 54913
rect 463 54776 947 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 947 54776
rect 463 54650 947 54700
rect 463 53299 946 53348
rect 463 53223 504 53299
rect 576 53223 626 53299
rect 698 53223 752 53299
rect 824 53223 946 53299
rect 463 53152 946 53223
rect 463 53076 504 53152
rect 576 53076 626 53152
rect 698 53076 752 53152
rect 824 53076 946 53152
rect 463 53015 946 53076
rect 463 52939 504 53015
rect 576 52939 626 53015
rect 698 52939 752 53015
rect 824 52939 946 53015
rect 463 52889 946 52939
rect 463 51060 946 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 946 51060
rect 463 50913 946 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 946 50913
rect 463 50776 946 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 946 50776
rect 463 50650 946 50700
rect 463 49301 946 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 946 49301
rect 463 49154 946 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 946 49154
rect 463 49017 946 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 946 49017
rect 463 48891 946 48941
rect 463 47060 946 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 946 47060
rect 463 46913 946 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 946 46913
rect 463 46776 946 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 946 46776
rect 463 46650 946 46700
rect 463 45301 946 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 946 45301
rect 463 45154 946 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 946 45154
rect 463 45017 946 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 946 45017
rect 463 44891 946 44941
rect 463 43060 946 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 946 43060
rect 463 42913 946 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 946 42913
rect 463 42776 946 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 946 42776
rect 463 42650 946 42700
rect 463 41300 946 41350
rect 463 41224 504 41300
rect 576 41224 626 41300
rect 698 41224 752 41300
rect 824 41224 946 41300
rect 463 41153 946 41224
rect 463 41077 504 41153
rect 576 41077 626 41153
rect 698 41077 752 41153
rect 824 41077 946 41153
rect 463 41016 946 41077
rect 463 40940 504 41016
rect 576 40940 626 41016
rect 698 40940 752 41016
rect 824 40940 946 41016
rect 463 40891 946 40940
rect 463 40890 836 40891
rect 944 35679 5204 35727
rect 944 35519 1306 35679
rect 1466 35519 1706 35679
rect 1866 35519 2106 35679
rect 2266 35519 2506 35679
rect 2666 35519 2906 35679
rect 3066 35519 3306 35679
rect 3466 35519 3706 35679
rect 3866 35519 4106 35679
rect 4266 35519 4506 35679
rect 4666 35519 5204 35679
rect 944 35496 5204 35519
rect 944 35336 1008 35496
rect 1168 35476 4983 35496
rect 1168 35336 1238 35476
rect 944 35138 1238 35336
rect 1868 35395 2503 35410
rect 1650 35321 1796 35329
rect 1650 35279 1662 35321
rect 1704 35279 1742 35321
rect 1784 35279 1796 35321
rect 1650 35241 1796 35279
rect 1868 35281 1885 35395
rect 2003 35281 2041 35395
rect 2159 35281 2197 35395
rect 2315 35281 2503 35395
rect 4914 35336 4983 35476
rect 5143 35336 5204 35496
rect 1868 35271 2503 35281
rect 1868 35270 2009 35271
rect 1650 35199 1662 35241
rect 1704 35199 1742 35241
rect 1784 35223 1796 35241
rect 2192 35230 2227 35237
rect 1784 35199 2192 35223
rect 1650 35191 2192 35199
rect 1650 35189 2227 35191
rect 944 35137 1126 35138
rect 944 35062 969 35137
rect 1041 35096 1126 35137
rect 1166 35096 1238 35138
rect 944 35021 1008 35062
rect 1168 35024 1238 35096
rect 1604 35125 1638 35139
rect 1919 35124 1954 35139
rect 1604 35052 1638 35059
rect 944 34946 972 35021
rect 1198 34949 1238 35024
rect 1762 34999 1796 35090
rect 1919 35069 1920 35124
rect 2192 35078 2227 35189
rect 2351 35085 2503 35271
rect 2539 35328 2685 35336
rect 2539 35286 2551 35328
rect 2593 35286 2631 35328
rect 2673 35286 2685 35328
rect 2539 35248 2685 35286
rect 2539 35206 2551 35248
rect 2593 35206 2631 35248
rect 2673 35206 2685 35248
rect 2539 35196 2685 35206
rect 2638 35085 2672 35196
rect 4914 35108 5204 35336
rect 4721 35096 5204 35108
rect 1919 35058 1953 35069
rect 944 34936 1008 34946
rect 1168 34936 1238 34949
rect 944 34696 1238 34936
rect 1604 34944 1638 34989
rect 1604 34797 1638 34889
rect 1762 34798 1796 34977
rect 1920 34944 1954 34989
rect 1920 34797 1954 34889
rect 2035 34944 2069 34997
rect 2035 34796 2069 34889
rect 2193 34795 2227 34988
rect 2351 34977 2514 35085
rect 2793 34977 2831 35085
rect 4721 35074 4983 35096
rect 2351 34944 2385 34977
rect 2351 34796 2385 34889
rect 2479 34949 2514 34977
rect 2479 34851 2514 34889
rect 2480 34797 2514 34851
rect 2638 34797 2672 34977
rect 2796 34949 2831 34977
rect 2796 34890 2797 34949
rect 2885 34981 2951 34982
rect 2885 34947 2901 34981
rect 2935 34947 2951 34981
rect 2885 34946 2951 34947
rect 4914 34936 4983 35074
rect 5143 34936 5204 35096
rect 2796 34851 2831 34890
rect 4315 34870 4557 34876
rect 2796 34797 2830 34851
rect 2900 34836 2921 34870
rect 2955 34836 2973 34870
rect 4315 34836 4339 34870
rect 4373 34836 4557 34870
rect 4315 34828 4557 34836
rect 4591 34871 4663 34876
rect 4591 34836 4615 34871
rect 4650 34836 4663 34871
rect 4591 34829 4663 34836
rect 4591 34828 4638 34829
rect 944 34536 1008 34696
rect 1168 34536 1238 34696
rect 944 34296 1238 34536
rect 4914 34696 5204 34936
rect 4914 34536 4983 34696
rect 5143 34536 5204 34696
rect 944 34136 1008 34296
rect 1168 34136 1238 34296
rect 1339 34260 1523 34269
rect 1339 34225 1479 34260
rect 1515 34225 1523 34260
rect 1339 34217 1523 34225
rect 2818 34202 2942 34343
rect 3740 34202 3864 34343
rect 4914 34296 5204 34536
rect 4632 34258 4704 34262
rect 4632 34224 4662 34258
rect 4696 34224 4704 34258
rect 4632 34207 4704 34224
rect 944 33896 1238 34136
rect 4914 34136 4983 34296
rect 5143 34136 5204 34296
rect 4914 34020 5204 34136
rect 4812 33986 5204 34020
rect 944 33736 1008 33896
rect 1168 33736 1238 33896
rect 4914 33896 5204 33986
rect 24526 34392 25428 34442
rect 24526 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 24526 34245 25428 34316
rect 24526 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 24526 34108 25428 34169
rect 24526 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 24526 33983 25428 34032
rect 24526 33982 25401 33983
rect 1573 33745 1769 33788
rect 944 33496 1238 33736
rect 2818 33663 2942 33804
rect 3740 33663 3864 33804
rect 4696 33748 4704 33780
rect 4675 33745 4704 33748
rect 4914 33736 4983 33896
rect 5143 33736 5204 33896
rect 944 33336 1008 33496
rect 1168 33336 1238 33496
rect 4914 33496 5204 33736
rect 1963 33442 1997 33465
rect 944 33096 1238 33336
rect 1680 33358 1739 33375
rect 1680 33310 1686 33358
rect 1732 33310 1739 33358
rect 2114 33312 2149 33451
rect 4914 33336 4983 33496
rect 5143 33336 5204 33496
rect 1680 33245 1739 33310
rect 1680 33200 1686 33245
rect 1732 33200 1739 33245
rect 1680 33187 1739 33200
rect 944 33079 1008 33096
rect 1168 33079 1238 33096
rect 944 32991 975 33079
rect 1203 32991 1238 33079
rect 1957 33144 1991 33257
rect 1957 33029 1991 33090
rect 2115 33029 2149 33256
rect 2273 33143 2307 33257
rect 2273 33029 2307 33089
rect 2436 33146 2471 33255
rect 2436 33029 2471 33095
rect 2595 33029 2629 33258
rect 2753 33143 2787 33267
rect 2944 33138 2962 33172
rect 2996 33138 3012 33172
rect 4315 33170 4557 33178
rect 4315 33136 4523 33170
rect 4315 33130 4557 33136
rect 4591 33170 4661 33178
rect 4591 33136 4615 33170
rect 4649 33136 4661 33170
rect 4591 33131 4661 33136
rect 4591 33130 4657 33131
rect 2753 33029 2787 33092
rect 4914 33096 5204 33336
rect 2913 33038 2956 33058
rect 944 32949 1008 32991
rect 1168 32949 1238 32991
rect 944 32861 975 32949
rect 1070 32861 1109 32936
rect 1204 32861 1238 32949
rect 1946 32921 1991 33029
rect 2273 32921 2318 33029
rect 2423 32921 2471 33029
rect 2753 32928 2800 33029
rect 2913 33003 2916 33038
rect 2953 33003 2956 33038
rect 2913 32987 2956 33003
rect 4914 32936 4983 33096
rect 5143 32936 5204 33096
rect 4914 32932 5204 32936
rect 944 32650 1238 32861
rect 2595 32838 2629 32921
rect 2753 32838 2879 32928
rect 4721 32898 5204 32932
rect 2538 32830 2685 32838
rect 2538 32788 2551 32830
rect 2593 32788 2631 32830
rect 2673 32788 2685 32830
rect 2538 32750 2685 32788
rect 2538 32711 2551 32750
rect 2593 32711 2631 32750
rect 2673 32711 2685 32750
rect 2538 32703 2685 32711
rect 2752 32830 2899 32838
rect 2752 32788 2765 32830
rect 2807 32788 2845 32830
rect 2887 32788 2899 32830
rect 2752 32747 2899 32788
rect 2752 32713 2765 32747
rect 2807 32713 2845 32747
rect 2887 32713 2899 32747
rect 2752 32707 2899 32713
rect 4914 32650 5204 32898
rect 944 32614 5204 32650
rect 944 32454 1008 32614
rect 1168 32454 1408 32614
rect 1568 32454 1808 32614
rect 1968 32454 2208 32614
rect 2368 32609 3408 32614
rect 2368 32454 2742 32609
rect 944 32449 2742 32454
rect 2902 32449 3069 32609
rect 3229 32454 3408 32609
rect 3568 32454 3808 32614
rect 3968 32454 4208 32614
rect 4368 32454 4608 32614
rect 4768 32454 4983 32614
rect 5143 32454 5204 32614
rect 3229 32449 5204 32454
rect 24526 32632 25428 32682
rect 24526 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 24526 32485 25428 32556
rect 944 32411 5203 32449
rect 24526 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 24526 32348 25428 32409
rect 24526 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 24526 32223 25428 32272
rect 24526 32222 25401 32223
rect 485 27110 847 27111
rect 463 27061 1116 27110
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 1116 27061
rect 463 26914 1116 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 1116 26914
rect 463 26777 1116 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 1116 26777
rect 463 26652 1116 26701
rect 463 26651 946 26652
rect 463 25294 1026 25350
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 1026 25294
rect 463 25147 1026 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 1026 25147
rect 463 25010 1026 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 1026 25010
rect 463 24890 1026 24934
rect 463 24885 863 24890
rect 463 24884 862 24885
rect 463 23060 946 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 946 23060
rect 463 22913 946 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 946 22913
rect 463 22776 946 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 946 22776
rect 463 22650 946 22700
rect 463 21300 946 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 946 21300
rect 463 21153 946 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 946 21153
rect 463 21016 946 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 946 21016
rect 463 20890 946 20940
rect 463 19060 946 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 946 19060
rect 463 18913 946 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 946 18913
rect 463 18776 946 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 946 18776
rect 463 18650 946 18700
rect 463 17301 946 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 946 17301
rect 463 17154 946 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 946 17154
rect 463 17017 946 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 946 17017
rect 463 16891 946 16941
rect 463 15060 946 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 946 15060
rect 463 14913 946 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 946 14913
rect 463 14776 946 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 946 14776
rect 463 14650 946 14700
rect 463 13300 946 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 946 13300
rect 463 13153 946 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 946 13153
rect 463 13016 946 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 946 13016
rect 463 12890 946 12940
rect 463 11060 946 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 946 11060
rect 463 10913 946 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 946 10913
rect 463 10776 946 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 946 10776
rect 463 10650 946 10700
rect 463 9300 946 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 946 9300
rect 463 9153 946 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 946 9153
rect 463 9016 946 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 946 9016
rect 463 8890 946 8940
rect 463 7061 946 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 946 7061
rect 463 6914 946 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 946 6914
rect 463 6777 946 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 946 6777
rect 463 6651 946 6701
rect 463 5299 946 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 946 5299
rect 463 5152 946 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 946 5152
rect 463 5015 946 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 946 5015
rect 463 4889 946 4939
rect 463 3061 946 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 946 3061
rect 463 2914 946 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 946 2914
rect 463 2777 946 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 946 2777
rect 463 2651 946 2701
rect 463 1300 946 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 946 1300
rect 463 1153 946 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 946 1153
rect 463 1016 946 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 946 1016
rect 463 890 946 940
<< viali >>
rect 503 67376 575 67452
rect 629 67376 701 67452
rect 749 67376 821 67452
rect 25068 67416 25140 67492
rect 25194 67416 25266 67492
rect 25314 67416 25386 67492
rect 503 67258 575 67334
rect 629 67258 701 67334
rect 749 67258 821 67334
rect 25068 67298 25140 67374
rect 25194 67298 25266 67374
rect 25314 67298 25386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 26010 65995 26082 66071
rect 26136 65995 26208 66071
rect 26256 65995 26328 66071
rect 26010 65877 26082 65953
rect 26136 65877 26208 65953
rect 26256 65877 26328 65953
rect 504 65224 576 65300
rect 626 65224 698 65300
rect 752 65224 824 65300
rect 504 65077 576 65153
rect 626 65077 698 65153
rect 752 65077 824 65153
rect 504 64940 576 65016
rect 626 64940 698 65016
rect 752 64940 824 65016
rect 503 64703 575 64779
rect 629 64703 701 64779
rect 749 64703 821 64779
rect 503 64585 575 64661
rect 629 64585 701 64661
rect 749 64585 821 64661
rect 25068 64619 25140 64695
rect 25194 64619 25266 64695
rect 25314 64619 25386 64695
rect 25068 64501 25140 64577
rect 25194 64501 25266 64577
rect 25314 64501 25386 64577
rect 503 63374 575 63450
rect 629 63374 701 63450
rect 749 63374 821 63450
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 503 63256 575 63332
rect 629 63256 701 63332
rect 749 63256 821 63332
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61982 26082 62058
rect 26136 61982 26208 62058
rect 26256 61982 26328 62058
rect 26010 61864 26082 61940
rect 26136 61864 26208 61940
rect 26256 61864 26328 61940
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60634 575 60710
rect 629 60634 701 60710
rect 749 60634 821 60710
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 503 60516 575 60592
rect 629 60516 701 60592
rect 749 60516 821 60592
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59456 575 59532
rect 629 59456 701 59532
rect 749 59456 821 59532
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 503 59338 575 59414
rect 629 59338 701 59414
rect 749 59338 821 59414
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57981 26082 58057
rect 26136 57981 26208 58057
rect 26256 57981 26328 58057
rect 26010 57863 26082 57939
rect 26136 57863 26208 57939
rect 26256 57863 26328 57939
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56608 575 56684
rect 629 56608 701 56684
rect 749 56608 821 56684
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 503 56490 575 56566
rect 629 56490 701 56566
rect 749 56490 821 56566
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55405 575 55481
rect 629 55405 701 55481
rect 749 55405 821 55481
rect 25068 55470 25140 55546
rect 25194 55470 25266 55546
rect 25314 55470 25386 55546
rect 503 55287 575 55363
rect 629 55287 701 55363
rect 749 55287 821 55363
rect 25068 55352 25140 55428
rect 25194 55352 25266 55428
rect 25314 55352 25386 55428
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 54020 26082 54096
rect 26136 54020 26208 54096
rect 26256 54020 26328 54096
rect 26010 53902 26082 53978
rect 26136 53902 26208 53978
rect 26256 53902 26328 53978
rect 504 53223 576 53299
rect 626 53223 698 53299
rect 752 53223 824 53299
rect 504 53076 576 53152
rect 626 53076 698 53152
rect 752 53076 824 53152
rect 504 52939 576 53015
rect 626 52939 698 53015
rect 752 52939 824 53015
rect 503 52628 575 52704
rect 629 52628 701 52704
rect 749 52628 821 52704
rect 503 52510 575 52586
rect 629 52510 701 52586
rect 749 52510 821 52586
rect 25068 52554 25140 52630
rect 25194 52554 25266 52630
rect 25314 52554 25386 52630
rect 25068 52436 25140 52512
rect 25194 52436 25266 52512
rect 25314 52436 25386 52512
rect 503 51421 575 51497
rect 629 51421 701 51497
rect 749 51421 821 51497
rect 503 51303 575 51379
rect 629 51303 701 51379
rect 749 51303 821 51379
rect 25068 51371 25140 51447
rect 25194 51371 25266 51447
rect 25314 51371 25386 51447
rect 25068 51253 25140 51329
rect 25194 51253 25266 51329
rect 25314 51253 25386 51329
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50003 26082 50079
rect 26136 50003 26208 50079
rect 26256 50003 26328 50079
rect 26010 49885 26082 49961
rect 26136 49885 26208 49961
rect 26256 49885 26328 49961
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48655 575 48731
rect 629 48655 701 48731
rect 749 48655 821 48731
rect 503 48537 575 48613
rect 629 48537 701 48613
rect 749 48537 821 48613
rect 25068 48499 25140 48575
rect 25194 48499 25266 48575
rect 25314 48499 25386 48575
rect 25068 48381 25140 48457
rect 25194 48381 25266 48457
rect 25314 48381 25386 48457
rect 503 47468 575 47544
rect 629 47468 701 47544
rect 749 47468 821 47544
rect 503 47350 575 47426
rect 629 47350 701 47426
rect 749 47350 821 47426
rect 25068 47364 25140 47440
rect 25194 47364 25266 47440
rect 25314 47364 25386 47440
rect 25068 47246 25140 47322
rect 25194 47246 25266 47322
rect 25314 47246 25386 47322
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46082 26082 46158
rect 26136 46082 26208 46158
rect 26256 46082 26328 46158
rect 26010 45964 26082 46040
rect 26136 45964 26208 46040
rect 26256 45964 26328 46040
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44646 575 44722
rect 629 44646 701 44722
rect 749 44646 821 44722
rect 25068 44605 25140 44681
rect 25194 44605 25266 44681
rect 25314 44605 25386 44681
rect 503 44528 575 44604
rect 629 44528 701 44604
rect 749 44528 821 44604
rect 25068 44487 25140 44563
rect 25194 44487 25266 44563
rect 25314 44487 25386 44563
rect 503 43493 575 43569
rect 629 43493 701 43569
rect 749 43493 821 43569
rect 25068 43452 25140 43528
rect 25194 43452 25266 43528
rect 25314 43452 25386 43528
rect 503 43375 575 43451
rect 629 43375 701 43451
rect 749 43375 821 43451
rect 25068 43334 25140 43410
rect 25194 43334 25266 43410
rect 25314 43334 25386 43410
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 41824 26082 41900
rect 26136 41824 26208 41900
rect 26256 41824 26328 41900
rect 26010 41706 26082 41782
rect 26136 41706 26208 41782
rect 26256 41706 26328 41782
rect 504 41224 576 41300
rect 626 41224 698 41300
rect 752 41224 824 41300
rect 504 41077 576 41153
rect 626 41077 698 41153
rect 752 41077 824 41153
rect 504 40940 576 41016
rect 626 40940 698 41016
rect 752 40940 824 41016
rect 503 40433 575 40509
rect 629 40433 701 40509
rect 749 40433 821 40509
rect 503 40315 575 40391
rect 629 40315 701 40391
rect 749 40315 821 40391
rect 25068 40336 25140 40412
rect 25194 40336 25266 40412
rect 25314 40336 25386 40412
rect 25068 40218 25140 40294
rect 25194 40218 25266 40294
rect 25314 40218 25386 40294
rect 1662 35279 1704 35321
rect 1742 35279 1784 35321
rect 1885 35281 2003 35395
rect 2041 35281 2159 35395
rect 2197 35281 2315 35395
rect 1662 35199 1704 35241
rect 1742 35199 1784 35241
rect 2192 35191 2227 35230
rect 969 35096 1041 35137
rect 1126 35096 1166 35138
rect 969 35062 1008 35096
rect 1008 35062 1041 35096
rect 1126 35063 1166 35096
rect 1604 35059 1638 35125
rect 972 34946 1008 35021
rect 1008 34946 1044 35021
rect 1126 34949 1168 35024
rect 1168 34949 1198 35024
rect 1920 35069 1954 35124
rect 2551 35286 2593 35328
rect 2631 35286 2673 35328
rect 2551 35206 2593 35248
rect 2631 35206 2673 35248
rect 1604 34889 1638 34944
rect 1920 34889 1954 34944
rect 2035 34889 2069 34944
rect 2351 34889 2385 34944
rect 2479 34889 2514 34949
rect 2797 34890 2831 34949
rect 2901 34947 2935 34981
rect 4251 34926 4285 34960
rect 2921 34836 2955 34870
rect 3253 34836 3288 34870
rect 3553 34836 3587 34870
rect 4105 34836 4139 34870
rect 4339 34836 4373 34870
rect 4615 34836 4650 34871
rect 1762 34706 1796 34782
rect 3800 34779 3835 34813
rect 1479 34225 1515 34260
rect 1715 34224 1749 34258
rect 1807 34227 1841 34261
rect 1899 34224 1933 34258
rect 2029 34218 2063 34252
rect 4662 34224 4696 34258
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 1481 33748 1515 33782
rect 1805 33753 1839 33787
rect 1889 33754 1923 33788
rect 1986 33748 2020 33782
rect 4662 33748 4696 33782
rect 1686 33310 1732 33358
rect 1686 33200 1732 33245
rect 975 32991 1008 33079
rect 1008 32991 1070 33079
rect 1108 32991 1168 33079
rect 1168 32991 1203 33079
rect 1957 33090 1991 33144
rect 2273 33089 2307 33143
rect 2436 33095 2471 33146
rect 3807 33193 3841 33227
rect 2753 33092 2787 33143
rect 2962 33138 2996 33172
rect 3237 33137 3271 33171
rect 3553 33136 3587 33170
rect 4105 33136 4139 33170
rect 4523 33136 4557 33170
rect 4615 33136 4649 33170
rect 4251 33046 4285 33080
rect 975 32936 1008 32949
rect 1008 32936 1070 32949
rect 1109 32936 1168 32949
rect 1168 32936 1204 32949
rect 975 32861 1070 32936
rect 1109 32861 1204 32936
rect 2916 33003 2953 33038
rect 2551 32788 2593 32830
rect 2631 32788 2673 32830
rect 2551 32711 2593 32750
rect 2631 32711 2673 32750
rect 2765 32788 2807 32830
rect 2845 32788 2887 32830
rect 2765 32713 2807 32747
rect 2845 32713 2887 32747
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal1 >>
rect 24946 67492 25426 67517
rect 463 67452 947 67477
rect 463 67376 503 67452
rect 575 67376 629 67452
rect 701 67376 749 67452
rect 821 67376 947 67452
rect 463 67334 947 67376
rect 463 67258 503 67334
rect 575 67258 629 67334
rect 701 67258 749 67334
rect 821 67258 947 67334
rect 24946 67416 25068 67492
rect 25140 67416 25194 67492
rect 25266 67416 25314 67492
rect 25386 67416 25426 67492
rect 24946 67374 25426 67416
rect 24946 67298 25068 67374
rect 25140 67298 25194 67374
rect 25266 67298 25314 67374
rect 25386 67298 25426 67374
rect 24946 67262 25426 67298
rect 463 67222 947 67258
rect 463 67060 863 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 66650 863 66700
rect 24946 66071 26370 66096
rect 24946 65995 26010 66071
rect 26082 65995 26136 66071
rect 26208 65995 26256 66071
rect 26328 65995 26370 66071
rect 24946 65953 26370 65995
rect 24946 65877 26010 65953
rect 26082 65877 26136 65953
rect 26208 65877 26256 65953
rect 26328 65877 26370 65953
rect 24946 65841 26370 65877
rect 463 65300 863 65349
rect 463 65224 504 65300
rect 576 65224 626 65300
rect 698 65224 752 65300
rect 824 65224 863 65300
rect 463 65153 863 65224
rect 463 65077 504 65153
rect 576 65077 626 65153
rect 698 65077 752 65153
rect 824 65077 863 65153
rect 463 65016 863 65077
rect 463 64940 504 65016
rect 576 64940 626 65016
rect 698 64940 752 65016
rect 824 64940 863 65016
rect 463 64890 863 64940
rect 463 64779 947 64804
rect 463 64703 503 64779
rect 575 64703 629 64779
rect 701 64703 749 64779
rect 821 64703 947 64779
rect 463 64661 947 64703
rect 463 64585 503 64661
rect 575 64585 629 64661
rect 701 64585 749 64661
rect 821 64585 947 64661
rect 463 64549 947 64585
rect 24946 64695 25428 64720
rect 24946 64619 25068 64695
rect 25140 64619 25194 64695
rect 25266 64619 25314 64695
rect 25386 64619 25428 64695
rect 24946 64577 25428 64619
rect 24946 64501 25068 64577
rect 25140 64501 25194 64577
rect 25266 64501 25314 64577
rect 25386 64501 25428 64577
rect 24946 64465 25428 64501
rect 24945 63517 24946 63530
rect 24945 63492 25426 63517
rect 463 63450 947 63475
rect 463 63374 503 63450
rect 575 63374 629 63450
rect 701 63374 749 63450
rect 821 63374 947 63450
rect 463 63332 947 63374
rect 463 63256 503 63332
rect 575 63256 629 63332
rect 701 63256 749 63332
rect 821 63256 947 63332
rect 24945 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25426 63492
rect 24945 63374 25426 63416
rect 24945 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25426 63374
rect 24945 63275 25426 63298
rect 24946 63262 25426 63275
rect 463 63220 947 63256
rect 463 63060 863 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 62650 863 62700
rect 24946 62058 26370 62083
rect 24946 61982 26010 62058
rect 26082 61982 26136 62058
rect 26208 61982 26256 62058
rect 26328 61982 26370 62058
rect 24946 61940 26370 61982
rect 24946 61864 26010 61940
rect 26082 61864 26136 61940
rect 26208 61864 26256 61940
rect 26328 61864 26370 61940
rect 24946 61828 26370 61864
rect 463 61301 863 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60891 863 60941
rect 463 60710 947 60735
rect 463 60634 503 60710
rect 575 60634 629 60710
rect 701 60634 749 60710
rect 821 60634 947 60710
rect 463 60592 947 60634
rect 463 60516 503 60592
rect 575 60516 629 60592
rect 701 60516 749 60592
rect 821 60516 947 60592
rect 463 60480 947 60516
rect 24945 60720 24946 60760
rect 24945 60695 25428 60720
rect 24945 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 24945 60577 25428 60619
rect 24945 60505 25068 60577
rect 24946 60501 25068 60505
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 24946 60465 25428 60501
rect 463 59532 947 59557
rect 463 59456 503 59532
rect 575 59456 629 59532
rect 701 59456 749 59532
rect 821 59456 947 59532
rect 463 59414 947 59456
rect 463 59338 503 59414
rect 575 59338 629 59414
rect 701 59338 749 59414
rect 821 59338 947 59414
rect 463 59302 947 59338
rect 24944 59492 25426 59517
rect 24944 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25426 59492
rect 24944 59374 25426 59416
rect 24944 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25426 59374
rect 24944 59262 25426 59298
rect 464 59068 864 59109
rect 463 59060 864 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 24946 58057 26370 58082
rect 24946 57981 26010 58057
rect 26082 57981 26136 58057
rect 26208 57981 26256 58057
rect 26328 57981 26370 58057
rect 24946 57939 26370 57981
rect 24946 57863 26010 57939
rect 26082 57863 26136 57939
rect 26208 57863 26256 57939
rect 26328 57863 26370 57939
rect 24946 57827 26370 57863
rect 463 57301 863 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56891 863 56941
rect 463 56684 949 56709
rect 463 56608 503 56684
rect 575 56608 629 56684
rect 701 56608 749 56684
rect 821 56608 949 56684
rect 463 56566 949 56608
rect 463 56490 503 56566
rect 575 56490 629 56566
rect 701 56490 749 56566
rect 821 56490 949 56566
rect 463 56454 949 56490
rect 24946 56695 25428 56720
rect 24946 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 24946 56577 25428 56619
rect 24946 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 24946 56465 25428 56501
rect 24945 55546 25427 55571
rect 463 55481 947 55506
rect 463 55405 503 55481
rect 575 55405 629 55481
rect 701 55405 749 55481
rect 821 55405 947 55481
rect 463 55363 947 55405
rect 463 55287 503 55363
rect 575 55287 629 55363
rect 701 55287 749 55363
rect 821 55287 947 55363
rect 24945 55470 25068 55546
rect 25140 55470 25194 55546
rect 25266 55470 25314 55546
rect 25386 55470 25427 55546
rect 24945 55428 25427 55470
rect 24945 55352 25068 55428
rect 25140 55352 25194 55428
rect 25266 55352 25314 55428
rect 25386 55352 25427 55428
rect 24945 55316 25427 55352
rect 463 55251 947 55287
rect 464 55068 864 55109
rect 463 55060 864 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 24946 54096 26370 54121
rect 24946 54020 26010 54096
rect 26082 54020 26136 54096
rect 26208 54020 26256 54096
rect 26328 54020 26370 54096
rect 24946 53978 26370 54020
rect 24946 53902 26010 53978
rect 26082 53902 26136 53978
rect 26208 53902 26256 53978
rect 26328 53902 26370 53978
rect 24946 53866 26370 53902
rect 463 53299 863 53348
rect 463 53223 504 53299
rect 576 53223 626 53299
rect 698 53223 752 53299
rect 824 53223 863 53299
rect 463 53152 863 53223
rect 463 53076 504 53152
rect 576 53076 626 53152
rect 698 53076 752 53152
rect 824 53076 863 53152
rect 463 53015 863 53076
rect 463 52939 504 53015
rect 576 52939 626 53015
rect 698 52939 752 53015
rect 824 52939 863 53015
rect 463 52889 863 52939
rect 463 52704 947 52729
rect 463 52628 503 52704
rect 575 52628 629 52704
rect 701 52628 749 52704
rect 821 52628 947 52704
rect 463 52586 947 52628
rect 463 52510 503 52586
rect 575 52510 629 52586
rect 701 52510 749 52586
rect 821 52510 947 52586
rect 463 52474 947 52510
rect 24946 52630 25428 52655
rect 24946 52554 25068 52630
rect 25140 52554 25194 52630
rect 25266 52554 25314 52630
rect 25386 52554 25428 52630
rect 24946 52512 25428 52554
rect 24946 52436 25068 52512
rect 25140 52436 25194 52512
rect 25266 52436 25314 52512
rect 25386 52436 25428 52512
rect 24946 52400 25428 52436
rect 463 51497 949 51522
rect 463 51421 503 51497
rect 575 51421 629 51497
rect 701 51421 749 51497
rect 821 51421 949 51497
rect 463 51379 949 51421
rect 463 51303 503 51379
rect 575 51303 629 51379
rect 701 51303 749 51379
rect 821 51303 949 51379
rect 463 51267 949 51303
rect 24945 51447 25427 51472
rect 24945 51371 25068 51447
rect 25140 51371 25194 51447
rect 25266 51371 25314 51447
rect 25386 51371 25427 51447
rect 24945 51329 25427 51371
rect 24945 51253 25068 51329
rect 25140 51253 25194 51329
rect 25266 51253 25314 51329
rect 25386 51253 25427 51329
rect 24945 51217 25427 51253
rect 463 51060 863 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 50650 863 50700
rect 24946 50079 26370 50104
rect 24946 50003 26010 50079
rect 26082 50003 26136 50079
rect 26208 50003 26256 50079
rect 26328 50003 26370 50079
rect 24946 49961 26370 50003
rect 24946 49885 26010 49961
rect 26082 49885 26136 49961
rect 26208 49885 26256 49961
rect 26328 49885 26370 49961
rect 24946 49849 26370 49885
rect 463 49301 863 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48891 863 48941
rect 463 48731 947 48756
rect 463 48655 503 48731
rect 575 48655 629 48731
rect 701 48655 749 48731
rect 821 48655 947 48731
rect 463 48613 947 48655
rect 463 48537 503 48613
rect 575 48537 629 48613
rect 701 48537 749 48613
rect 821 48537 947 48613
rect 463 48501 947 48537
rect 24946 48575 25428 48600
rect 24946 48499 25068 48575
rect 25140 48499 25194 48575
rect 25266 48499 25314 48575
rect 25386 48499 25428 48575
rect 24946 48457 25428 48499
rect 24946 48381 25068 48457
rect 25140 48381 25194 48457
rect 25266 48381 25314 48457
rect 25386 48381 25428 48457
rect 24946 48345 25428 48381
rect 463 47544 947 47569
rect 463 47468 503 47544
rect 575 47468 629 47544
rect 701 47468 749 47544
rect 821 47468 947 47544
rect 463 47426 947 47468
rect 463 47350 503 47426
rect 575 47350 629 47426
rect 701 47350 749 47426
rect 821 47350 947 47426
rect 463 47314 947 47350
rect 24946 47440 25428 47465
rect 24946 47364 25068 47440
rect 25140 47364 25194 47440
rect 25266 47364 25314 47440
rect 25386 47364 25428 47440
rect 24946 47322 25428 47364
rect 24946 47246 25068 47322
rect 25140 47246 25194 47322
rect 25266 47246 25314 47322
rect 25386 47246 25428 47322
rect 24946 47210 25428 47246
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 24946 46158 26370 46183
rect 24946 46082 26010 46158
rect 26082 46082 26136 46158
rect 26208 46082 26256 46158
rect 26328 46082 26370 46158
rect 24946 46040 26370 46082
rect 24946 45964 26010 46040
rect 26082 45964 26136 46040
rect 26208 45964 26256 46040
rect 26328 45964 26370 46040
rect 24946 45928 26370 45964
rect 463 45301 863 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44891 863 44941
rect 463 44722 947 44747
rect 463 44646 503 44722
rect 575 44646 629 44722
rect 701 44646 749 44722
rect 821 44646 947 44722
rect 463 44604 947 44646
rect 463 44528 503 44604
rect 575 44528 629 44604
rect 701 44528 749 44604
rect 821 44528 947 44604
rect 463 44492 947 44528
rect 24946 44681 25428 44706
rect 24946 44605 25068 44681
rect 25140 44605 25194 44681
rect 25266 44605 25314 44681
rect 25386 44605 25428 44681
rect 24946 44563 25428 44605
rect 24946 44487 25068 44563
rect 25140 44487 25194 44563
rect 25266 44487 25314 44563
rect 25386 44487 25428 44563
rect 24946 44451 25428 44487
rect 463 43569 947 43594
rect 463 43493 503 43569
rect 575 43493 629 43569
rect 701 43493 749 43569
rect 821 43493 947 43569
rect 463 43451 947 43493
rect 463 43375 503 43451
rect 575 43375 629 43451
rect 701 43375 749 43451
rect 821 43375 947 43451
rect 463 43339 947 43375
rect 24946 43528 25428 43553
rect 24946 43452 25068 43528
rect 25140 43452 25194 43528
rect 25266 43452 25314 43528
rect 25386 43452 25428 43528
rect 24946 43410 25428 43452
rect 24946 43334 25068 43410
rect 25140 43334 25194 43410
rect 25266 43334 25314 43410
rect 25386 43334 25428 43410
rect 24946 43298 25428 43334
rect 463 43060 863 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 42650 863 42700
rect 24946 41900 26370 41925
rect 24946 41824 26010 41900
rect 26082 41824 26136 41900
rect 26208 41824 26256 41900
rect 26328 41824 26370 41900
rect 24946 41782 26370 41824
rect 24946 41706 26010 41782
rect 26082 41706 26136 41782
rect 26208 41706 26256 41782
rect 26328 41706 26370 41782
rect 24946 41670 26370 41706
rect 463 41300 863 41350
rect 463 41224 504 41300
rect 576 41224 626 41300
rect 698 41224 752 41300
rect 824 41224 863 41300
rect 463 41153 863 41224
rect 463 41077 504 41153
rect 576 41077 626 41153
rect 698 41077 752 41153
rect 824 41077 863 41153
rect 463 41016 863 41077
rect 463 40940 504 41016
rect 576 40940 626 41016
rect 698 40940 752 41016
rect 824 40940 863 41016
rect 463 40891 863 40940
rect 463 40890 836 40891
rect 463 40509 946 40534
rect 463 40433 503 40509
rect 575 40433 629 40509
rect 701 40433 749 40509
rect 821 40433 946 40509
rect 463 40391 946 40433
rect 463 40315 503 40391
rect 575 40315 629 40391
rect 701 40315 749 40391
rect 821 40315 946 40391
rect 463 40279 946 40315
rect 24946 40412 25428 40437
rect 24946 40336 25068 40412
rect 25140 40336 25194 40412
rect 25266 40336 25314 40412
rect 25386 40336 25428 40412
rect 24946 40294 25428 40336
rect 24946 40218 25068 40294
rect 25140 40218 25194 40294
rect 25266 40218 25314 40294
rect 25386 40218 25428 40294
rect 24946 40182 25428 40218
rect 3287 35752 4421 35753
rect 0 35741 25902 35752
rect 0 35661 32 35741
rect 112 35661 157 35741
rect 237 35661 282 35741
rect 362 35726 25902 35741
rect 362 35661 25535 35726
rect 0 35646 25535 35661
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 0 35635 25902 35646
rect 0 35555 32 35635
rect 112 35555 157 35635
rect 237 35555 282 35635
rect 362 35606 25902 35635
rect 362 35555 25534 35606
rect 0 35526 25534 35555
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 0 35497 25902 35526
rect 1868 35395 2335 35410
rect 1650 35321 1796 35329
rect 1650 35269 1662 35321
rect 1714 35269 1732 35321
rect 1784 35269 1796 35321
rect 1868 35281 1885 35395
rect 2003 35281 2041 35395
rect 2159 35281 2197 35395
rect 2315 35281 2335 35395
rect 1868 35270 2335 35281
rect 2539 35328 2685 35336
rect 2539 35276 2551 35328
rect 2603 35276 2621 35328
rect 2673 35276 2685 35328
rect 1650 35251 1796 35269
rect 1650 35199 1662 35251
rect 1714 35199 1732 35251
rect 1784 35233 1796 35251
rect 2539 35258 2685 35276
rect 2167 35233 2239 35236
rect 1784 35230 2239 35233
rect 1784 35199 2192 35230
rect 1650 35191 2192 35199
rect 2227 35191 2239 35230
rect 2539 35206 2551 35258
rect 2603 35206 2621 35258
rect 2673 35206 2685 35258
rect 2539 35196 2685 35206
rect 1650 35189 2239 35191
rect 2167 35185 2239 35189
rect 944 35139 1238 35173
rect 463 35138 2973 35139
rect 463 35137 1126 35138
rect 463 35130 969 35137
rect 463 35052 479 35130
rect 561 35052 593 35130
rect 675 35052 707 35130
rect 789 35062 969 35130
rect 1041 35063 1126 35137
rect 1166 35125 2973 35138
rect 1166 35063 1604 35125
rect 1041 35062 1604 35063
rect 789 35059 1604 35062
rect 1638 35124 2973 35125
rect 1638 35069 1920 35124
rect 1954 35069 2973 35124
rect 1638 35059 2973 35069
rect 789 35052 2973 35059
rect 463 35043 2973 35052
rect 944 35024 1238 35043
rect 944 35021 1126 35024
rect 944 34946 972 35021
rect 1044 34949 1126 35021
rect 1198 34949 1238 35024
rect 2889 34982 2950 34987
rect 2889 34981 3370 34982
rect 1044 34946 1238 34949
rect 944 34923 1238 34946
rect 1592 34944 1966 34954
rect 1592 34889 1604 34944
rect 1638 34889 1920 34944
rect 1954 34889 1966 34944
rect 1592 34882 1966 34889
rect 2022 34944 2397 34954
rect 2022 34889 2035 34944
rect 2069 34889 2351 34944
rect 2385 34889 2397 34944
rect 2022 34882 2397 34889
rect 2467 34949 2843 34955
rect 2467 34889 2479 34949
rect 2514 34890 2797 34949
rect 2831 34890 2843 34949
rect 2889 34947 2901 34981
rect 2935 34947 3370 34981
rect 24527 34972 25428 34998
rect 2889 34946 3370 34947
rect 2889 34941 2950 34946
rect 2514 34889 2843 34890
rect 2467 34883 2843 34889
rect 2900 34870 3301 34876
rect 2900 34836 2921 34870
rect 2955 34836 3253 34870
rect 3288 34836 3301 34870
rect 2900 34829 3301 34836
rect 1755 34782 1802 34794
rect 1495 34774 1569 34781
rect 1495 34722 1503 34774
rect 1563 34770 1569 34774
rect 1755 34770 1762 34782
rect 1563 34722 1762 34770
rect 1495 34717 1762 34722
rect 1755 34706 1762 34717
rect 1796 34706 1802 34782
rect 3342 34772 3370 34946
rect 3615 34960 4297 34966
rect 3615 34926 4251 34960
rect 4285 34926 4297 34960
rect 3615 34920 4297 34926
rect 3523 34828 3529 34880
rect 3581 34876 3587 34880
rect 3615 34876 3650 34920
rect 24527 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 4610 34879 4662 34885
rect 4092 34876 4156 34878
rect 3581 34870 3650 34876
rect 3587 34836 3650 34870
rect 3581 34830 3650 34836
rect 4075 34870 4385 34876
rect 4075 34836 4105 34870
rect 4139 34836 4339 34870
rect 4373 34836 4385 34870
rect 4075 34830 4385 34836
rect 3581 34828 3587 34830
rect 4092 34826 4156 34830
rect 4608 34829 4610 34877
rect 3792 34813 3841 34825
rect 4610 34821 4662 34827
rect 24527 34852 25428 34892
rect 3792 34779 3800 34813
rect 3835 34779 3841 34813
rect 3792 34772 3841 34779
rect 3341 34737 3841 34772
rect 24527 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 24527 34743 25428 34772
rect 1755 34694 1802 34706
rect 0 34586 1593 34595
rect 0 34508 16 34586
rect 98 34508 130 34586
rect 212 34508 244 34586
rect 326 34508 1593 34586
rect 0 34499 1593 34508
rect 25028 34392 25428 34442
rect 3608 34348 3660 34354
rect 1893 34305 3608 34334
rect 1465 34217 1471 34269
rect 1523 34268 1529 34269
rect 1523 34258 1773 34268
rect 1523 34224 1715 34258
rect 1749 34224 1773 34258
rect 1523 34218 1773 34224
rect 1801 34261 1847 34275
rect 1801 34227 1807 34261
rect 1841 34227 1847 34261
rect 1523 34217 1529 34218
rect 1801 34210 1847 34227
rect 1893 34258 1941 34305
rect 3608 34290 3660 34296
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 1893 34224 1899 34258
rect 1933 34224 1941 34258
rect 1893 34212 1941 34224
rect 2019 34252 2076 34275
rect 2019 34218 2029 34252
rect 2063 34218 2076 34252
rect 1805 34184 1847 34210
rect 2019 34202 2076 34218
rect 4652 34267 4704 34273
rect 4652 34209 4704 34215
rect 25028 34245 25428 34316
rect 2019 34184 2063 34202
rect 1805 34155 2063 34184
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 463 34042 2056 34051
rect 463 33964 479 34042
rect 561 33964 593 34042
rect 675 33964 707 34042
rect 789 33964 2056 34042
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 25028 33983 25428 34032
rect 25028 33982 25401 33983
rect 463 33955 2056 33964
rect 3517 33889 3523 33897
rect 1874 33854 3523 33889
rect 1457 33738 1463 33790
rect 1515 33738 1539 33790
rect 1799 33787 1845 33851
rect 1799 33753 1805 33787
rect 1839 33753 1845 33787
rect 1799 33708 1845 33753
rect 1874 33788 1940 33854
rect 3517 33845 3523 33854
rect 3575 33845 3581 33897
rect 1874 33754 1889 33788
rect 1923 33754 1940 33788
rect 1874 33738 1940 33754
rect 1980 33782 2032 33795
rect 1980 33748 1986 33782
rect 2020 33748 2032 33782
rect 1980 33708 2032 33748
rect 4652 33791 4704 33797
rect 4652 33733 4704 33739
rect 1799 33680 2032 33708
rect 0 33498 1317 33507
rect 0 33420 16 33498
rect 98 33420 130 33498
rect 212 33420 244 33498
rect 326 33420 1317 33498
rect 0 33411 1317 33420
rect 24526 33476 25902 33502
rect 24526 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 1680 33358 1739 33375
rect 1680 33306 1683 33358
rect 1735 33306 1739 33358
rect 1680 33252 1739 33306
rect 24526 33356 25902 33396
rect 1680 33200 1683 33252
rect 1735 33200 1739 33252
rect 1680 33150 1739 33200
rect 3332 33265 3841 33300
rect 2927 33172 3295 33178
rect 1680 33144 2320 33150
rect 944 33079 1238 33111
rect 1680 33090 1957 33144
rect 1991 33143 2320 33144
rect 1991 33090 2273 33143
rect 1680 33089 2273 33090
rect 2307 33089 2320 33143
rect 1680 33084 2320 33089
rect 2416 33146 2804 33152
rect 2416 33095 2436 33146
rect 2471 33143 2804 33146
rect 2471 33095 2753 33143
rect 2416 33092 2753 33095
rect 2787 33092 2804 33143
rect 2927 33138 2962 33172
rect 2996 33171 3295 33172
rect 2996 33138 3237 33171
rect 2927 33137 3237 33138
rect 3271 33137 3295 33171
rect 2927 33131 3295 33137
rect 2416 33085 2804 33092
rect 1680 33083 1739 33084
rect 1945 33083 2320 33084
rect 944 32991 975 33079
rect 1070 32991 1108 33079
rect 1203 32991 1238 33079
rect 3332 33069 3375 33265
rect 3806 33233 3841 33265
rect 24526 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 24526 33247 25902 33276
rect 3801 33227 3848 33233
rect 3801 33193 3807 33227
rect 3841 33193 3848 33227
rect 3547 33176 3553 33182
rect 3523 33130 3553 33176
rect 3605 33130 3646 33182
rect 3801 33181 3848 33193
rect 4609 33181 4661 33187
rect 2969 33058 3375 33069
rect 2910 33038 3375 33058
rect 3610 33086 3646 33130
rect 4075 33178 4156 33180
rect 4075 33170 4569 33178
rect 4075 33136 4105 33170
rect 4139 33136 4523 33170
rect 4557 33136 4569 33170
rect 4075 33130 4569 33136
rect 4075 33128 4156 33130
rect 4609 33123 4661 33129
rect 3610 33080 4297 33086
rect 3610 33046 4251 33080
rect 4285 33046 4297 33080
rect 3610 33038 4297 33046
rect 2910 33003 2916 33038
rect 2953 33034 3375 33038
rect 2953 33023 2987 33034
rect 2953 33003 2959 33023
rect 2910 32991 2959 33003
rect 944 32963 1238 32991
rect 463 32954 2973 32963
rect 463 32876 479 32954
rect 561 32876 593 32954
rect 675 32876 707 32954
rect 789 32949 2973 32954
rect 789 32876 975 32949
rect 463 32867 975 32876
rect 944 32861 975 32867
rect 1070 32861 1109 32949
rect 1204 32867 2973 32949
rect 1204 32861 1238 32867
rect 944 32835 1238 32861
rect 2538 32830 2685 32838
rect 2538 32778 2551 32830
rect 2603 32778 2621 32830
rect 2673 32778 2685 32830
rect 2538 32763 2685 32778
rect 2538 32711 2551 32763
rect 2603 32711 2621 32763
rect 2673 32711 2685 32763
rect 2538 32649 2685 32711
rect 2752 32830 2899 32838
rect 2752 32778 2765 32830
rect 2817 32778 2835 32830
rect 2887 32778 2899 32830
rect 2752 32765 2899 32778
rect 2752 32713 2765 32765
rect 2817 32713 2835 32765
rect 2887 32713 2899 32765
rect 2752 32707 2899 32713
rect 25028 32632 25428 32682
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 32223 25428 32272
rect 25028 32222 25401 32223
rect 24514 31917 25427 31943
rect 24514 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25427 31917
rect 24514 31797 25427 31837
rect 24514 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25427 31797
rect 24514 31688 25427 31717
rect 463 28302 25428 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 463 28184 25428 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 463 28073 25428 28108
rect 463 28072 1825 28073
rect 2313 28072 25428 28073
rect 463 27520 946 27545
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 946 27520
rect 463 27402 946 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 946 27402
rect 463 27290 946 27326
rect 24946 27520 25428 27545
rect 24946 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 24946 27402 25428 27444
rect 24946 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 24946 27290 25428 27326
rect 463 27061 863 27111
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 26651 863 26701
rect 24946 26130 26370 26155
rect 24946 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 24946 26012 26370 26054
rect 24946 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 24946 25900 26370 25936
rect 463 25294 863 25350
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24884 862 24885
rect 944 24681 946 24880
rect 463 24608 946 24633
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 946 24608
rect 463 24490 946 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 946 24490
rect 463 24378 946 24414
rect 24946 24559 25428 24584
rect 24946 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 24946 24441 25428 24483
rect 24946 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 24946 24329 25428 24365
rect 463 23604 946 23629
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 946 23604
rect 463 23486 946 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 946 23486
rect 463 23374 946 23410
rect 24945 23442 25427 23467
rect 24945 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25427 23442
rect 24945 23324 25427 23366
rect 24945 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25427 23324
rect 24945 23212 25427 23248
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 24946 21971 26370 21996
rect 24946 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 24946 21853 26370 21895
rect 24946 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 24946 21741 26370 21777
rect 463 21300 863 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20890 863 20940
rect 463 20626 947 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 947 20626
rect 463 20508 947 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 947 20508
rect 463 20396 947 20432
rect 24946 20599 25428 20624
rect 24946 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 24946 20481 25428 20523
rect 24946 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 24946 20369 25428 20405
rect 463 19544 947 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 947 19544
rect 463 19426 947 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 947 19426
rect 463 19314 947 19350
rect 24946 19424 25428 19449
rect 24946 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 24946 19306 25428 19348
rect 24946 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 24946 19194 25428 19230
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 24946 18181 26370 18206
rect 24946 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 24946 18063 26370 18105
rect 24946 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 24946 17951 26370 17987
rect 463 17301 863 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16891 863 16941
rect 463 16669 947 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 947 16669
rect 463 16551 947 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 947 16551
rect 463 16439 947 16475
rect 24945 16583 25427 16608
rect 24945 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25427 16583
rect 24945 16465 25427 16507
rect 24945 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25427 16465
rect 24945 16353 25427 16389
rect 463 15568 947 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 947 15568
rect 463 15450 947 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 947 15450
rect 463 15338 947 15374
rect 24945 15412 25427 15437
rect 24945 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25427 15412
rect 24945 15294 25427 15336
rect 24945 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25427 15294
rect 24945 15182 25427 15218
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 24946 14074 26370 14099
rect 24946 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 24946 13956 26370 13998
rect 24946 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 24946 13844 26370 13880
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12702 948 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 948 12702
rect 463 12584 948 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 948 12584
rect 463 12472 948 12508
rect 24945 12651 25427 12676
rect 24945 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25427 12651
rect 24945 12533 25427 12575
rect 24945 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25427 12533
rect 24945 12421 25427 12457
rect 463 11486 949 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 949 11486
rect 463 11368 949 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 949 11368
rect 463 11256 949 11292
rect 24945 11437 25427 11462
rect 24945 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25427 11437
rect 24945 11319 25427 11361
rect 24945 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25427 11319
rect 24945 11207 25427 11243
rect 463 11060 863 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 10650 863 10700
rect 24946 10256 26370 10281
rect 24946 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 24946 10138 26370 10180
rect 24946 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 24946 10026 26370 10062
rect 463 9300 863 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8890 863 8940
rect 463 8621 947 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 947 8621
rect 463 8503 947 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 947 8503
rect 463 8391 947 8427
rect 24946 8594 25428 8619
rect 24946 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 24946 8476 25428 8518
rect 24946 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 24946 8364 25428 8400
rect 463 7499 947 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 947 7499
rect 463 7381 947 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 947 7381
rect 463 7269 947 7305
rect 24946 7437 25427 7462
rect 24946 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25427 7437
rect 24946 7319 25427 7361
rect 24946 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25427 7319
rect 24946 7207 25427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 24946 6292 26370 6317
rect 24946 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 24946 6174 26370 6216
rect 24946 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 24946 6062 26370 6098
rect 463 5299 863 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4889 863 4939
rect 463 4639 946 4664
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 946 4639
rect 463 4521 946 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 946 4521
rect 463 4409 946 4445
rect 24946 4594 25428 4619
rect 24946 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 24946 4476 25428 4518
rect 24946 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 24946 4364 25428 4400
rect 463 3528 946 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 946 3528
rect 463 3410 946 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 946 3410
rect 463 3298 946 3334
rect 24946 3437 25427 3462
rect 24946 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25427 3437
rect 24946 3319 25427 3361
rect 24946 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25427 3319
rect 24946 3207 25427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 24946 2280 26370 2305
rect 24946 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 24946 2162 26370 2204
rect 24946 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 24946 2050 26370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 948 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 948 705
rect 463 587 948 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 948 587
rect 463 475 948 511
rect 24946 594 25428 619
rect 24946 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 24946 476 25428 518
rect 24946 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 24946 364 25428 400
<< via1 >>
rect 503 67376 575 67452
rect 629 67376 701 67452
rect 749 67376 821 67452
rect 503 67258 575 67334
rect 629 67258 701 67334
rect 749 67258 821 67334
rect 25068 67416 25140 67492
rect 25194 67416 25266 67492
rect 25314 67416 25386 67492
rect 25068 67298 25140 67374
rect 25194 67298 25266 67374
rect 25314 67298 25386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 26010 65995 26082 66071
rect 26136 65995 26208 66071
rect 26256 65995 26328 66071
rect 26010 65877 26082 65953
rect 26136 65877 26208 65953
rect 26256 65877 26328 65953
rect 504 65224 576 65300
rect 626 65224 698 65300
rect 752 65224 824 65300
rect 504 65077 576 65153
rect 626 65077 698 65153
rect 752 65077 824 65153
rect 504 64940 576 65016
rect 626 64940 698 65016
rect 752 64940 824 65016
rect 503 64703 575 64779
rect 629 64703 701 64779
rect 749 64703 821 64779
rect 503 64585 575 64661
rect 629 64585 701 64661
rect 749 64585 821 64661
rect 25068 64619 25140 64695
rect 25194 64619 25266 64695
rect 25314 64619 25386 64695
rect 25068 64501 25140 64577
rect 25194 64501 25266 64577
rect 25314 64501 25386 64577
rect 503 63374 575 63450
rect 629 63374 701 63450
rect 749 63374 821 63450
rect 503 63256 575 63332
rect 629 63256 701 63332
rect 749 63256 821 63332
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61982 26082 62058
rect 26136 61982 26208 62058
rect 26256 61982 26328 62058
rect 26010 61864 26082 61940
rect 26136 61864 26208 61940
rect 26256 61864 26328 61940
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60634 575 60710
rect 629 60634 701 60710
rect 749 60634 821 60710
rect 503 60516 575 60592
rect 629 60516 701 60592
rect 749 60516 821 60592
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59456 575 59532
rect 629 59456 701 59532
rect 749 59456 821 59532
rect 503 59338 575 59414
rect 629 59338 701 59414
rect 749 59338 821 59414
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57981 26082 58057
rect 26136 57981 26208 58057
rect 26256 57981 26328 58057
rect 26010 57863 26082 57939
rect 26136 57863 26208 57939
rect 26256 57863 26328 57939
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56608 575 56684
rect 629 56608 701 56684
rect 749 56608 821 56684
rect 503 56490 575 56566
rect 629 56490 701 56566
rect 749 56490 821 56566
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55405 575 55481
rect 629 55405 701 55481
rect 749 55405 821 55481
rect 503 55287 575 55363
rect 629 55287 701 55363
rect 749 55287 821 55363
rect 25068 55470 25140 55546
rect 25194 55470 25266 55546
rect 25314 55470 25386 55546
rect 25068 55352 25140 55428
rect 25194 55352 25266 55428
rect 25314 55352 25386 55428
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 54020 26082 54096
rect 26136 54020 26208 54096
rect 26256 54020 26328 54096
rect 26010 53902 26082 53978
rect 26136 53902 26208 53978
rect 26256 53902 26328 53978
rect 504 53223 576 53299
rect 626 53223 698 53299
rect 752 53223 824 53299
rect 504 53076 576 53152
rect 626 53076 698 53152
rect 752 53076 824 53152
rect 504 52939 576 53015
rect 626 52939 698 53015
rect 752 52939 824 53015
rect 503 52628 575 52704
rect 629 52628 701 52704
rect 749 52628 821 52704
rect 503 52510 575 52586
rect 629 52510 701 52586
rect 749 52510 821 52586
rect 25068 52554 25140 52630
rect 25194 52554 25266 52630
rect 25314 52554 25386 52630
rect 25068 52436 25140 52512
rect 25194 52436 25266 52512
rect 25314 52436 25386 52512
rect 503 51421 575 51497
rect 629 51421 701 51497
rect 749 51421 821 51497
rect 503 51303 575 51379
rect 629 51303 701 51379
rect 749 51303 821 51379
rect 25068 51371 25140 51447
rect 25194 51371 25266 51447
rect 25314 51371 25386 51447
rect 25068 51253 25140 51329
rect 25194 51253 25266 51329
rect 25314 51253 25386 51329
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50003 26082 50079
rect 26136 50003 26208 50079
rect 26256 50003 26328 50079
rect 26010 49885 26082 49961
rect 26136 49885 26208 49961
rect 26256 49885 26328 49961
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48655 575 48731
rect 629 48655 701 48731
rect 749 48655 821 48731
rect 503 48537 575 48613
rect 629 48537 701 48613
rect 749 48537 821 48613
rect 25068 48499 25140 48575
rect 25194 48499 25266 48575
rect 25314 48499 25386 48575
rect 25068 48381 25140 48457
rect 25194 48381 25266 48457
rect 25314 48381 25386 48457
rect 503 47468 575 47544
rect 629 47468 701 47544
rect 749 47468 821 47544
rect 503 47350 575 47426
rect 629 47350 701 47426
rect 749 47350 821 47426
rect 25068 47364 25140 47440
rect 25194 47364 25266 47440
rect 25314 47364 25386 47440
rect 25068 47246 25140 47322
rect 25194 47246 25266 47322
rect 25314 47246 25386 47322
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46082 26082 46158
rect 26136 46082 26208 46158
rect 26256 46082 26328 46158
rect 26010 45964 26082 46040
rect 26136 45964 26208 46040
rect 26256 45964 26328 46040
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44646 575 44722
rect 629 44646 701 44722
rect 749 44646 821 44722
rect 503 44528 575 44604
rect 629 44528 701 44604
rect 749 44528 821 44604
rect 25068 44605 25140 44681
rect 25194 44605 25266 44681
rect 25314 44605 25386 44681
rect 25068 44487 25140 44563
rect 25194 44487 25266 44563
rect 25314 44487 25386 44563
rect 503 43493 575 43569
rect 629 43493 701 43569
rect 749 43493 821 43569
rect 503 43375 575 43451
rect 629 43375 701 43451
rect 749 43375 821 43451
rect 25068 43452 25140 43528
rect 25194 43452 25266 43528
rect 25314 43452 25386 43528
rect 25068 43334 25140 43410
rect 25194 43334 25266 43410
rect 25314 43334 25386 43410
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 41824 26082 41900
rect 26136 41824 26208 41900
rect 26256 41824 26328 41900
rect 26010 41706 26082 41782
rect 26136 41706 26208 41782
rect 26256 41706 26328 41782
rect 504 41224 576 41300
rect 626 41224 698 41300
rect 752 41224 824 41300
rect 504 41077 576 41153
rect 626 41077 698 41153
rect 752 41077 824 41153
rect 504 40940 576 41016
rect 626 40940 698 41016
rect 752 40940 824 41016
rect 503 40433 575 40509
rect 629 40433 701 40509
rect 749 40433 821 40509
rect 503 40315 575 40391
rect 629 40315 701 40391
rect 749 40315 821 40391
rect 25068 40336 25140 40412
rect 25194 40336 25266 40412
rect 25314 40336 25386 40412
rect 25068 40218 25140 40294
rect 25194 40218 25266 40294
rect 25314 40218 25386 40294
rect 32 35661 112 35741
rect 157 35661 237 35741
rect 282 35661 362 35741
rect 25535 35646 25615 35726
rect 25660 35646 25740 35726
rect 25785 35646 25865 35726
rect 32 35555 112 35635
rect 157 35555 237 35635
rect 282 35555 362 35635
rect 25534 35526 25614 35606
rect 25659 35526 25739 35606
rect 25784 35526 25864 35606
rect 1662 35279 1704 35321
rect 1704 35279 1714 35321
rect 1662 35269 1714 35279
rect 1732 35279 1742 35321
rect 1742 35279 1784 35321
rect 1732 35269 1784 35279
rect 1885 35281 2003 35395
rect 2041 35281 2159 35395
rect 2197 35281 2315 35395
rect 2551 35286 2593 35328
rect 2593 35286 2603 35328
rect 2551 35276 2603 35286
rect 2621 35286 2631 35328
rect 2631 35286 2673 35328
rect 2621 35276 2673 35286
rect 1662 35241 1714 35251
rect 1662 35199 1704 35241
rect 1704 35199 1714 35241
rect 1732 35241 1784 35251
rect 1732 35199 1742 35241
rect 1742 35199 1784 35241
rect 2551 35248 2603 35258
rect 2551 35206 2593 35248
rect 2593 35206 2603 35248
rect 2621 35248 2673 35258
rect 2621 35206 2631 35248
rect 2631 35206 2673 35248
rect 479 35052 561 35130
rect 593 35052 675 35130
rect 707 35052 789 35130
rect 1503 34722 1563 34774
rect 3529 34870 3581 34880
rect 25061 34892 25141 34972
rect 25186 34892 25266 34972
rect 25311 34892 25391 34972
rect 3529 34836 3553 34870
rect 3553 34836 3581 34870
rect 3529 34828 3581 34836
rect 4610 34871 4662 34879
rect 4610 34836 4615 34871
rect 4615 34836 4650 34871
rect 4650 34836 4662 34871
rect 4610 34827 4662 34836
rect 25060 34772 25140 34852
rect 25185 34772 25265 34852
rect 25310 34772 25390 34852
rect 16 34508 98 34586
rect 130 34508 212 34586
rect 244 34508 326 34586
rect 1471 34260 1523 34269
rect 1471 34225 1479 34260
rect 1479 34225 1515 34260
rect 1515 34225 1523 34260
rect 1471 34217 1523 34225
rect 3608 34296 3660 34348
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 4652 34258 4704 34267
rect 4652 34224 4662 34258
rect 4662 34224 4696 34258
rect 4696 34224 4704 34258
rect 4652 34215 4704 34224
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 479 33964 561 34042
rect 593 33964 675 34042
rect 707 33964 789 34042
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 1463 33782 1515 33790
rect 1463 33748 1481 33782
rect 1481 33748 1515 33782
rect 1463 33738 1515 33748
rect 3523 33845 3575 33897
rect 4652 33782 4704 33791
rect 4652 33748 4662 33782
rect 4662 33748 4696 33782
rect 4696 33748 4704 33782
rect 4652 33739 4704 33748
rect 16 33420 98 33498
rect 130 33420 212 33498
rect 244 33420 326 33498
rect 24560 33396 24640 33476
rect 24685 33396 24765 33476
rect 24810 33396 24890 33476
rect 25535 33396 25615 33476
rect 25660 33396 25740 33476
rect 25785 33396 25865 33476
rect 1683 33310 1686 33358
rect 1686 33310 1732 33358
rect 1732 33310 1735 33358
rect 1683 33306 1735 33310
rect 1683 33245 1735 33252
rect 1683 33200 1686 33245
rect 1686 33200 1732 33245
rect 1732 33200 1735 33245
rect 24559 33276 24639 33356
rect 24684 33276 24764 33356
rect 24809 33276 24889 33356
rect 25534 33276 25614 33356
rect 25659 33276 25739 33356
rect 25784 33276 25864 33356
rect 3553 33170 3605 33182
rect 3553 33136 3587 33170
rect 3587 33136 3605 33170
rect 3553 33130 3605 33136
rect 4609 33170 4661 33181
rect 4609 33136 4615 33170
rect 4615 33136 4649 33170
rect 4649 33136 4661 33170
rect 4609 33129 4661 33136
rect 479 32876 561 32954
rect 593 32876 675 32954
rect 707 32876 789 32954
rect 2551 32788 2593 32830
rect 2593 32788 2603 32830
rect 2551 32778 2603 32788
rect 2621 32788 2631 32830
rect 2631 32788 2673 32830
rect 2621 32778 2673 32788
rect 2551 32750 2603 32763
rect 2551 32711 2593 32750
rect 2593 32711 2603 32750
rect 2621 32750 2673 32763
rect 2621 32711 2631 32750
rect 2631 32711 2673 32750
rect 2765 32788 2807 32830
rect 2807 32788 2817 32830
rect 2765 32778 2817 32788
rect 2835 32788 2845 32830
rect 2845 32788 2887 32830
rect 2835 32778 2887 32788
rect 2765 32747 2817 32765
rect 2765 32713 2807 32747
rect 2807 32713 2817 32747
rect 2835 32747 2887 32765
rect 2835 32713 2845 32747
rect 2845 32713 2887 32747
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 25060 31837 25140 31917
rect 25185 31837 25265 31917
rect 25310 31837 25390 31917
rect 25059 31717 25139 31797
rect 25184 31717 25264 31797
rect 25309 31717 25389 31797
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal2 >>
rect 25026 67492 25426 67517
rect 463 67452 864 67477
rect 463 67376 503 67452
rect 575 67376 629 67452
rect 701 67376 749 67452
rect 821 67376 864 67452
rect 463 67334 864 67376
rect 463 67258 503 67334
rect 575 67258 629 67334
rect 701 67258 749 67334
rect 821 67258 864 67334
rect 25026 67416 25068 67492
rect 25140 67416 25194 67492
rect 25266 67416 25314 67492
rect 25386 67416 25426 67492
rect 25026 67374 25426 67416
rect 25026 67298 25068 67374
rect 25140 67298 25194 67374
rect 25266 67298 25314 67374
rect 25386 67298 25426 67374
rect 25026 67262 25426 67298
rect 463 67222 864 67258
rect 463 67060 863 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 66650 863 66700
rect 25970 66071 26370 66096
rect 25970 65995 26010 66071
rect 26082 65995 26136 66071
rect 26208 65995 26256 66071
rect 26328 65995 26370 66071
rect 25970 65953 26370 65995
rect 25970 65877 26010 65953
rect 26082 65877 26136 65953
rect 26208 65877 26256 65953
rect 26328 65877 26370 65953
rect 25970 65841 26370 65877
rect 463 65300 863 65349
rect 463 65224 504 65300
rect 576 65224 626 65300
rect 698 65224 752 65300
rect 824 65224 863 65300
rect 463 65153 863 65224
rect 463 65077 504 65153
rect 576 65077 626 65153
rect 698 65077 752 65153
rect 824 65077 863 65153
rect 463 65016 863 65077
rect 463 64940 504 65016
rect 576 64940 626 65016
rect 698 64940 752 65016
rect 824 64940 863 65016
rect 463 64890 863 64940
rect 463 64779 864 64804
rect 463 64703 503 64779
rect 575 64703 629 64779
rect 701 64703 749 64779
rect 821 64703 864 64779
rect 463 64661 864 64703
rect 463 64585 503 64661
rect 575 64585 629 64661
rect 701 64585 749 64661
rect 821 64585 864 64661
rect 463 64549 864 64585
rect 25028 64695 25428 64720
rect 25028 64619 25068 64695
rect 25140 64619 25194 64695
rect 25266 64619 25314 64695
rect 25386 64619 25428 64695
rect 25028 64577 25428 64619
rect 25028 64501 25068 64577
rect 25140 64501 25194 64577
rect 25266 64501 25314 64577
rect 25386 64501 25428 64577
rect 25028 64465 25428 64501
rect 25026 63492 25426 63517
rect 463 63450 864 63475
rect 463 63374 503 63450
rect 575 63374 629 63450
rect 701 63374 749 63450
rect 821 63374 864 63450
rect 463 63332 864 63374
rect 463 63256 503 63332
rect 575 63256 629 63332
rect 701 63256 749 63332
rect 821 63256 864 63332
rect 25026 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25426 63492
rect 25026 63374 25426 63416
rect 25026 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25426 63374
rect 25026 63262 25426 63298
rect 463 63220 864 63256
rect 463 63060 863 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 62650 863 62700
rect 25970 62058 26370 62083
rect 25970 61982 26010 62058
rect 26082 61982 26136 62058
rect 26208 61982 26256 62058
rect 26328 61982 26370 62058
rect 25970 61940 26370 61982
rect 25970 61864 26010 61940
rect 26082 61864 26136 61940
rect 26208 61864 26256 61940
rect 26328 61864 26370 61940
rect 25970 61828 26370 61864
rect 463 61301 863 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60891 863 60941
rect 463 60710 864 60735
rect 463 60634 503 60710
rect 575 60634 629 60710
rect 701 60634 749 60710
rect 821 60634 864 60710
rect 463 60592 864 60634
rect 463 60516 503 60592
rect 575 60516 629 60592
rect 701 60516 749 60592
rect 821 60516 864 60592
rect 463 60480 864 60516
rect 25028 60695 25428 60720
rect 25028 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 25028 60577 25428 60619
rect 25028 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 25028 60465 25428 60501
rect 463 59532 864 59557
rect 463 59456 503 59532
rect 575 59456 629 59532
rect 701 59456 749 59532
rect 821 59456 864 59532
rect 463 59414 864 59456
rect 463 59338 503 59414
rect 575 59338 629 59414
rect 701 59338 749 59414
rect 821 59338 864 59414
rect 463 59302 864 59338
rect 25026 59492 25426 59517
rect 25026 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25426 59492
rect 25026 59374 25426 59416
rect 25026 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25426 59374
rect 25026 59262 25426 59298
rect 464 59068 864 59109
rect 463 59060 864 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 25970 58057 26370 58082
rect 25970 57981 26010 58057
rect 26082 57981 26136 58057
rect 26208 57981 26256 58057
rect 26328 57981 26370 58057
rect 25970 57939 26370 57981
rect 25970 57863 26010 57939
rect 26082 57863 26136 57939
rect 26208 57863 26256 57939
rect 26328 57863 26370 57939
rect 25970 57827 26370 57863
rect 463 57301 863 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56891 863 56941
rect 463 56684 866 56709
rect 463 56608 503 56684
rect 575 56608 629 56684
rect 701 56608 749 56684
rect 821 56608 866 56684
rect 463 56566 866 56608
rect 463 56490 503 56566
rect 575 56490 629 56566
rect 701 56490 749 56566
rect 821 56490 866 56566
rect 463 56454 866 56490
rect 25028 56695 25428 56720
rect 25028 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 25028 56577 25428 56619
rect 25028 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 25028 56465 25428 56501
rect 25027 55546 25427 55571
rect 463 55481 864 55506
rect 463 55405 503 55481
rect 575 55405 629 55481
rect 701 55405 749 55481
rect 821 55405 864 55481
rect 463 55363 864 55405
rect 463 55287 503 55363
rect 575 55287 629 55363
rect 701 55287 749 55363
rect 821 55287 864 55363
rect 25027 55470 25068 55546
rect 25140 55470 25194 55546
rect 25266 55470 25314 55546
rect 25386 55470 25427 55546
rect 25027 55428 25427 55470
rect 25027 55352 25068 55428
rect 25140 55352 25194 55428
rect 25266 55352 25314 55428
rect 25386 55352 25427 55428
rect 25027 55316 25427 55352
rect 463 55251 864 55287
rect 464 55068 864 55109
rect 463 55060 864 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 25970 54096 26370 54121
rect 25970 54020 26010 54096
rect 26082 54020 26136 54096
rect 26208 54020 26256 54096
rect 26328 54020 26370 54096
rect 25970 53978 26370 54020
rect 25970 53902 26010 53978
rect 26082 53902 26136 53978
rect 26208 53902 26256 53978
rect 26328 53902 26370 53978
rect 25970 53866 26370 53902
rect 463 53299 863 53348
rect 463 53223 504 53299
rect 576 53223 626 53299
rect 698 53223 752 53299
rect 824 53223 863 53299
rect 463 53152 863 53223
rect 463 53076 504 53152
rect 576 53076 626 53152
rect 698 53076 752 53152
rect 824 53076 863 53152
rect 463 53015 863 53076
rect 463 52939 504 53015
rect 576 52939 626 53015
rect 698 52939 752 53015
rect 824 52939 863 53015
rect 463 52889 863 52939
rect 463 52704 864 52729
rect 463 52628 503 52704
rect 575 52628 629 52704
rect 701 52628 749 52704
rect 821 52628 864 52704
rect 463 52586 864 52628
rect 463 52510 503 52586
rect 575 52510 629 52586
rect 701 52510 749 52586
rect 821 52510 864 52586
rect 463 52474 864 52510
rect 25028 52630 25428 52655
rect 25028 52554 25068 52630
rect 25140 52554 25194 52630
rect 25266 52554 25314 52630
rect 25386 52554 25428 52630
rect 25028 52512 25428 52554
rect 25028 52436 25068 52512
rect 25140 52436 25194 52512
rect 25266 52436 25314 52512
rect 25386 52436 25428 52512
rect 25028 52400 25428 52436
rect 463 51497 866 51522
rect 463 51421 503 51497
rect 575 51421 629 51497
rect 701 51421 749 51497
rect 821 51421 866 51497
rect 463 51379 866 51421
rect 463 51303 503 51379
rect 575 51303 629 51379
rect 701 51303 749 51379
rect 821 51303 866 51379
rect 463 51267 866 51303
rect 25027 51447 25427 51472
rect 25027 51371 25068 51447
rect 25140 51371 25194 51447
rect 25266 51371 25314 51447
rect 25386 51371 25427 51447
rect 25027 51329 25427 51371
rect 25027 51253 25068 51329
rect 25140 51253 25194 51329
rect 25266 51253 25314 51329
rect 25386 51253 25427 51329
rect 25027 51217 25427 51253
rect 463 51060 863 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 50650 863 50700
rect 25970 50079 26370 50104
rect 25970 50003 26010 50079
rect 26082 50003 26136 50079
rect 26208 50003 26256 50079
rect 26328 50003 26370 50079
rect 25970 49961 26370 50003
rect 25970 49885 26010 49961
rect 26082 49885 26136 49961
rect 26208 49885 26256 49961
rect 26328 49885 26370 49961
rect 25970 49849 26370 49885
rect 463 49301 863 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48891 863 48941
rect 463 48731 864 48756
rect 463 48655 503 48731
rect 575 48655 629 48731
rect 701 48655 749 48731
rect 821 48655 864 48731
rect 463 48613 864 48655
rect 463 48537 503 48613
rect 575 48537 629 48613
rect 701 48537 749 48613
rect 821 48537 864 48613
rect 463 48501 864 48537
rect 25028 48575 25428 48600
rect 25028 48499 25068 48575
rect 25140 48499 25194 48575
rect 25266 48499 25314 48575
rect 25386 48499 25428 48575
rect 25028 48457 25428 48499
rect 25028 48381 25068 48457
rect 25140 48381 25194 48457
rect 25266 48381 25314 48457
rect 25386 48381 25428 48457
rect 25028 48345 25428 48381
rect 463 47544 864 47569
rect 463 47468 503 47544
rect 575 47468 629 47544
rect 701 47468 749 47544
rect 821 47468 864 47544
rect 463 47426 864 47468
rect 463 47350 503 47426
rect 575 47350 629 47426
rect 701 47350 749 47426
rect 821 47350 864 47426
rect 463 47314 864 47350
rect 25028 47440 25428 47465
rect 25028 47364 25068 47440
rect 25140 47364 25194 47440
rect 25266 47364 25314 47440
rect 25386 47364 25428 47440
rect 25028 47322 25428 47364
rect 25028 47246 25068 47322
rect 25140 47246 25194 47322
rect 25266 47246 25314 47322
rect 25386 47246 25428 47322
rect 25028 47210 25428 47246
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 25970 46158 26370 46183
rect 25970 46082 26010 46158
rect 26082 46082 26136 46158
rect 26208 46082 26256 46158
rect 26328 46082 26370 46158
rect 25970 46040 26370 46082
rect 25970 45964 26010 46040
rect 26082 45964 26136 46040
rect 26208 45964 26256 46040
rect 26328 45964 26370 46040
rect 25970 45928 26370 45964
rect 463 45301 863 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44891 863 44941
rect 463 44722 864 44747
rect 463 44646 503 44722
rect 575 44646 629 44722
rect 701 44646 749 44722
rect 821 44646 864 44722
rect 463 44604 864 44646
rect 463 44528 503 44604
rect 575 44528 629 44604
rect 701 44528 749 44604
rect 821 44528 864 44604
rect 463 44492 864 44528
rect 25028 44681 25428 44706
rect 25028 44605 25068 44681
rect 25140 44605 25194 44681
rect 25266 44605 25314 44681
rect 25386 44605 25428 44681
rect 25028 44563 25428 44605
rect 25028 44487 25068 44563
rect 25140 44487 25194 44563
rect 25266 44487 25314 44563
rect 25386 44487 25428 44563
rect 25028 44451 25428 44487
rect 463 43569 864 43594
rect 463 43493 503 43569
rect 575 43493 629 43569
rect 701 43493 749 43569
rect 821 43493 864 43569
rect 463 43451 864 43493
rect 463 43375 503 43451
rect 575 43375 629 43451
rect 701 43375 749 43451
rect 821 43375 864 43451
rect 463 43339 864 43375
rect 25028 43528 25428 43553
rect 25028 43452 25068 43528
rect 25140 43452 25194 43528
rect 25266 43452 25314 43528
rect 25386 43452 25428 43528
rect 25028 43410 25428 43452
rect 25028 43334 25068 43410
rect 25140 43334 25194 43410
rect 25266 43334 25314 43410
rect 25386 43334 25428 43410
rect 25028 43298 25428 43334
rect 463 43060 863 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 42650 863 42700
rect 25970 41900 26370 41925
rect 25970 41824 26010 41900
rect 26082 41824 26136 41900
rect 26208 41824 26256 41900
rect 26328 41824 26370 41900
rect 25970 41782 26370 41824
rect 25970 41706 26010 41782
rect 26082 41706 26136 41782
rect 26208 41706 26256 41782
rect 26328 41706 26370 41782
rect 25970 41670 26370 41706
rect 463 41300 863 41350
rect 463 41224 504 41300
rect 576 41224 626 41300
rect 698 41224 752 41300
rect 824 41224 863 41300
rect 463 41153 863 41224
rect 463 41077 504 41153
rect 576 41077 626 41153
rect 698 41077 752 41153
rect 824 41077 863 41153
rect 463 41016 863 41077
rect 463 40940 504 41016
rect 576 40940 626 41016
rect 698 40940 752 41016
rect 824 40940 863 41016
rect 463 40891 863 40940
rect 463 40890 836 40891
rect 463 40509 863 40534
rect 463 40433 503 40509
rect 575 40433 629 40509
rect 701 40433 749 40509
rect 821 40433 863 40509
rect 463 40391 863 40433
rect 463 40315 503 40391
rect 575 40315 629 40391
rect 701 40315 749 40391
rect 821 40315 863 40391
rect 463 40279 863 40315
rect 25028 40412 25428 40437
rect 25028 40336 25068 40412
rect 25140 40336 25194 40412
rect 25266 40336 25314 40412
rect 25386 40336 25428 40412
rect 25028 40294 25428 40336
rect 25028 40218 25068 40294
rect 25140 40218 25194 40294
rect 25266 40218 25314 40294
rect 25386 40218 25428 40294
rect 25028 40182 25428 40218
rect 1650 35925 2398 35940
rect 1650 35869 2257 35925
rect 2313 35869 2337 35925
rect 2393 35869 2398 35925
rect 1650 35845 2398 35869
rect 1650 35789 2257 35845
rect 2313 35789 2337 35845
rect 2393 35789 2398 35845
rect 1650 35776 2398 35789
rect 1650 35774 2396 35776
rect 0 35741 400 35752
rect 0 35661 32 35741
rect 112 35661 157 35741
rect 237 35661 282 35741
rect 362 35661 400 35741
rect 0 35635 400 35661
rect 0 35555 32 35635
rect 112 35555 157 35635
rect 237 35555 282 35635
rect 362 35555 400 35635
rect 0 35528 400 35555
rect 1411 35320 1569 35333
rect 1411 35319 1498 35320
rect 1411 35263 1416 35319
rect 1472 35264 1498 35319
rect 1554 35264 1569 35320
rect 1472 35263 1569 35264
rect 1411 35240 1569 35263
rect 1411 35239 1499 35240
rect 1411 35183 1417 35239
rect 1473 35184 1499 35239
rect 1555 35184 1569 35240
rect 1650 35321 1796 35774
rect 2468 35711 2867 40000
rect 3352 35904 3502 35919
rect 3352 35848 3361 35904
rect 3417 35848 3441 35904
rect 3497 35848 3502 35904
rect 3352 35824 3502 35848
rect 3352 35768 3361 35824
rect 3417 35768 3441 35824
rect 3497 35768 3502 35824
rect 3352 35755 3502 35768
rect 3352 35754 3500 35755
rect 1867 35438 2868 35711
rect 1650 35269 1662 35321
rect 1714 35269 1732 35321
rect 1784 35269 1796 35321
rect 1650 35251 1796 35269
rect 1650 35199 1662 35251
rect 1714 35199 1732 35251
rect 1784 35199 1796 35251
rect 1650 35189 1796 35199
rect 1868 35410 2267 35438
rect 1868 35395 2335 35410
rect 1868 35281 1885 35395
rect 2003 35281 2041 35395
rect 2159 35281 2197 35395
rect 2315 35281 2335 35395
rect 1868 35270 2335 35281
rect 2538 35328 2685 35336
rect 2538 35276 2551 35328
rect 2603 35276 2621 35328
rect 2673 35276 2685 35328
rect 1473 35183 1569 35184
rect 1411 35169 1569 35183
rect 463 35130 805 35139
rect 463 35052 479 35130
rect 561 35052 593 35130
rect 675 35052 707 35130
rect 789 35052 805 35130
rect 463 35043 805 35052
rect 1495 34774 1569 35169
rect 1495 34722 1503 34774
rect 1563 34722 1569 34774
rect 1495 34717 1569 34722
rect 0 34586 342 34595
rect 0 34508 16 34586
rect 98 34508 130 34586
rect 212 34508 244 34586
rect 326 34508 342 34586
rect 0 34499 342 34508
rect 1471 34269 1523 34275
rect 1471 34211 1523 34217
rect 463 34042 805 34051
rect 463 33964 479 34042
rect 561 33964 593 34042
rect 675 33964 707 34042
rect 789 33964 805 34042
rect 463 33955 805 33964
rect 1471 33797 1504 34211
rect 1463 33790 1515 33797
rect 1463 33732 1515 33738
rect 0 33498 342 33507
rect 0 33420 16 33498
rect 98 33420 130 33498
rect 212 33420 244 33498
rect 326 33420 342 33498
rect 0 33411 342 33420
rect 1680 33358 1739 35189
rect 1680 33306 1683 33358
rect 1735 33306 1739 33358
rect 1680 33252 1739 33306
rect 1680 33200 1683 33252
rect 1735 33200 1739 33252
rect 1680 33187 1739 33200
rect 463 32954 805 32963
rect 463 32876 479 32954
rect 561 32876 593 32954
rect 675 32876 707 32954
rect 789 32876 805 32954
rect 463 32867 805 32876
rect 1868 28936 2267 35270
rect 2538 35258 2685 35276
rect 2538 35206 2551 35258
rect 2603 35206 2621 35258
rect 2673 35206 2685 35258
rect 2751 35318 2899 35332
rect 2751 35262 2760 35318
rect 2816 35317 2899 35318
rect 2816 35262 2840 35317
rect 2751 35261 2840 35262
rect 2896 35261 2899 35317
rect 2751 35253 2899 35261
rect 2538 32830 2685 35206
rect 2538 32778 2551 32830
rect 2603 32778 2621 32830
rect 2673 32778 2685 32830
rect 2538 32763 2685 32778
rect 2538 32711 2551 32763
rect 2603 32711 2621 32763
rect 2673 32711 2685 32763
rect 2538 32476 2685 32711
rect 2752 35237 2899 35253
rect 2752 35181 2761 35237
rect 2817 35181 2841 35237
rect 2897 35181 2899 35237
rect 2752 32830 2899 35181
rect 3352 35317 3499 35754
rect 25502 35726 25902 35752
rect 25502 35646 25535 35726
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 25502 35606 25902 35646
rect 25502 35526 25534 35606
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 25502 35497 25902 35526
rect 3352 35261 3360 35317
rect 3416 35316 3499 35317
rect 3416 35261 3440 35316
rect 3352 35260 3440 35261
rect 3496 35260 3499 35316
rect 3352 35236 3499 35260
rect 3352 35180 3361 35236
rect 3417 35180 3441 35236
rect 3497 35180 3499 35236
rect 3352 35169 3499 35180
rect 25028 34972 25428 34998
rect 25028 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 3523 34828 3529 34880
rect 3581 34828 3587 34880
rect 4610 34879 4704 34885
rect 3537 33897 3568 34828
rect 4662 34827 4704 34879
rect 4610 34821 4704 34827
rect 3608 34348 3660 34354
rect 3608 34290 3660 34296
rect 3517 33845 3523 33897
rect 3575 33845 3581 33897
rect 3620 33185 3649 34290
rect 4652 34267 4704 34821
rect 25028 34852 25428 34892
rect 25028 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 25028 34743 25428 34772
rect 4652 34209 4704 34215
rect 25028 34392 25428 34442
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 25028 34245 25428 34316
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 25028 33983 25428 34032
rect 25028 33982 25401 33983
rect 4652 33791 4704 33797
rect 4652 33187 4704 33739
rect 24527 33476 24927 33502
rect 24527 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 24927 33476
rect 24527 33356 24927 33396
rect 24527 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 24927 33356
rect 24527 33247 24927 33276
rect 25502 33476 25902 33502
rect 25502 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 25502 33356 25902 33396
rect 25502 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 25502 33247 25902 33276
rect 3536 33182 3649 33185
rect 3536 33130 3553 33182
rect 3605 33130 3649 33182
rect 3536 33126 3649 33130
rect 4609 33181 4704 33187
rect 4661 33129 4704 33181
rect 4609 33123 4704 33129
rect 2752 32778 2765 32830
rect 2817 32778 2835 32830
rect 2887 32778 2899 32830
rect 2752 32765 2899 32778
rect 2752 32713 2765 32765
rect 2817 32713 2835 32765
rect 2887 32713 2899 32765
rect 2752 32707 2899 32713
rect 2535 32475 2685 32476
rect 25028 32632 25428 32682
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 2535 32463 2689 32475
rect 2535 32401 2544 32463
rect 2600 32401 2624 32463
rect 2680 32401 2689 32463
rect 2535 32391 2689 32401
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 32223 25428 32272
rect 25028 32222 25401 32223
rect 25027 31917 25427 31943
rect 25027 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25427 31917
rect 25027 31797 25427 31837
rect 25027 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25427 31797
rect 25027 31688 25427 31717
rect 1868 28710 2742 28936
rect 1866 28485 2742 28710
rect 463 28302 866 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 866 28302
rect 463 28184 866 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 866 28184
rect 463 28072 866 28108
rect 2306 27967 2742 28485
rect 25025 28302 25428 28360
rect 25025 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 25025 28184 25428 28226
rect 25025 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 25025 28072 25428 28108
rect 463 27520 863 27545
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 863 27520
rect 463 27402 863 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 863 27402
rect 463 27290 863 27326
rect 25028 27520 25428 27545
rect 25028 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 25028 27402 25428 27444
rect 25028 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 25028 27290 25428 27326
rect 463 27061 863 27111
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 26651 863 26701
rect 25970 26130 26370 26155
rect 25970 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 25970 26012 26370 26054
rect 25970 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 25970 25900 26370 25936
rect 463 25294 863 25349
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24884 862 24885
rect 463 24608 863 24633
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 863 24608
rect 463 24490 863 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 863 24490
rect 463 24378 863 24414
rect 25028 24559 25428 24584
rect 25028 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 25028 24441 25428 24483
rect 25028 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 25028 24329 25428 24365
rect 463 23604 863 23629
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 863 23604
rect 463 23486 863 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 863 23486
rect 463 23374 863 23410
rect 25027 23442 25427 23467
rect 25027 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25427 23442
rect 25027 23324 25427 23366
rect 25027 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25427 23324
rect 25027 23212 25427 23248
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 25970 21971 26370 21996
rect 25970 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 25970 21853 26370 21895
rect 25970 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 25970 21741 26370 21777
rect 463 21300 863 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20890 863 20940
rect 463 20626 864 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 864 20626
rect 463 20508 864 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 864 20508
rect 463 20396 864 20432
rect 25028 20599 25428 20624
rect 25028 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 25028 20481 25428 20523
rect 25028 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 25028 20369 25428 20405
rect 463 19544 864 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 864 19544
rect 463 19426 864 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 864 19426
rect 463 19314 864 19350
rect 25028 19424 25428 19449
rect 25028 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 25028 19306 25428 19348
rect 25028 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 25028 19194 25428 19230
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 25970 18181 26370 18206
rect 25970 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 25970 18063 26370 18105
rect 25970 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 25970 17951 26370 17987
rect 463 17301 863 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16891 863 16941
rect 463 16669 864 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 864 16669
rect 463 16551 864 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 864 16551
rect 463 16439 864 16475
rect 25027 16583 25427 16608
rect 25027 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25427 16583
rect 25027 16465 25427 16507
rect 25027 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25427 16465
rect 25027 16353 25427 16389
rect 463 15568 864 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 864 15568
rect 463 15450 864 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 864 15450
rect 463 15338 864 15374
rect 25027 15412 25427 15437
rect 25027 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25427 15412
rect 25027 15294 25427 15336
rect 25027 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25427 15294
rect 25027 15182 25427 15218
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 25970 14074 26370 14099
rect 25970 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 25970 13956 26370 13998
rect 25970 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 25970 13844 26370 13880
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12702 865 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 865 12702
rect 463 12584 865 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 865 12584
rect 463 12472 865 12508
rect 25027 12651 25427 12676
rect 25027 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25427 12651
rect 25027 12533 25427 12575
rect 25027 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25427 12533
rect 25027 12421 25427 12457
rect 463 11486 866 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 866 11486
rect 463 11368 866 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 866 11368
rect 463 11256 866 11292
rect 25027 11437 25427 11462
rect 25027 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25427 11437
rect 25027 11319 25427 11361
rect 25027 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25427 11319
rect 25027 11207 25427 11243
rect 463 11060 863 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 10650 863 10700
rect 25970 10256 26370 10281
rect 25970 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 25970 10138 26370 10180
rect 25970 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 25970 10026 26370 10062
rect 463 9300 863 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8890 863 8940
rect 463 8621 864 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 864 8621
rect 463 8503 864 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 864 8503
rect 463 8391 864 8427
rect 25028 8594 25428 8619
rect 25028 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 25028 8476 25428 8518
rect 25028 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 25028 8364 25428 8400
rect 463 7499 864 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 864 7499
rect 463 7381 864 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 864 7381
rect 463 7269 864 7305
rect 25027 7437 25427 7462
rect 25027 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25427 7437
rect 25027 7319 25427 7361
rect 25027 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25427 7319
rect 25027 7207 25427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 25970 6292 26370 6317
rect 25970 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 25970 6174 26370 6216
rect 25970 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 25970 6062 26370 6098
rect 463 5299 863 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4889 863 4939
rect 463 4639 863 4664
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 863 4639
rect 463 4521 863 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 863 4521
rect 463 4409 863 4445
rect 25028 4594 25428 4619
rect 25028 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 25028 4476 25428 4518
rect 25028 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 25028 4364 25428 4400
rect 463 3528 863 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3298 863 3334
rect 25027 3437 25427 3462
rect 25027 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25427 3437
rect 25027 3319 25427 3361
rect 25027 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25427 3319
rect 25027 3207 25427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 25970 2280 26370 2305
rect 25970 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 25970 2162 26370 2204
rect 25970 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 25970 2050 26370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 25028 594 25428 619
rect 25028 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 25028 476 25428 518
rect 25028 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 25028 364 25428 400
<< via2 >>
rect 503 67376 575 67452
rect 629 67376 701 67452
rect 749 67376 821 67452
rect 503 67258 575 67334
rect 629 67258 701 67334
rect 749 67258 821 67334
rect 25068 67416 25140 67492
rect 25194 67416 25266 67492
rect 25314 67416 25386 67492
rect 25068 67298 25140 67374
rect 25194 67298 25266 67374
rect 25314 67298 25386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 26010 65995 26082 66071
rect 26136 65995 26208 66071
rect 26256 65995 26328 66071
rect 26010 65877 26082 65953
rect 26136 65877 26208 65953
rect 26256 65877 26328 65953
rect 504 65224 576 65300
rect 626 65224 698 65300
rect 752 65224 824 65300
rect 504 65077 576 65153
rect 626 65077 698 65153
rect 752 65077 824 65153
rect 504 64940 576 65016
rect 626 64940 698 65016
rect 752 64940 824 65016
rect 503 64703 575 64779
rect 629 64703 701 64779
rect 749 64703 821 64779
rect 503 64585 575 64661
rect 629 64585 701 64661
rect 749 64585 821 64661
rect 25068 64619 25140 64695
rect 25194 64619 25266 64695
rect 25314 64619 25386 64695
rect 25068 64501 25140 64577
rect 25194 64501 25266 64577
rect 25314 64501 25386 64577
rect 503 63374 575 63450
rect 629 63374 701 63450
rect 749 63374 821 63450
rect 503 63256 575 63332
rect 629 63256 701 63332
rect 749 63256 821 63332
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61982 26082 62058
rect 26136 61982 26208 62058
rect 26256 61982 26328 62058
rect 26010 61864 26082 61940
rect 26136 61864 26208 61940
rect 26256 61864 26328 61940
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60634 575 60710
rect 629 60634 701 60710
rect 749 60634 821 60710
rect 503 60516 575 60592
rect 629 60516 701 60592
rect 749 60516 821 60592
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59456 575 59532
rect 629 59456 701 59532
rect 749 59456 821 59532
rect 503 59338 575 59414
rect 629 59338 701 59414
rect 749 59338 821 59414
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57981 26082 58057
rect 26136 57981 26208 58057
rect 26256 57981 26328 58057
rect 26010 57863 26082 57939
rect 26136 57863 26208 57939
rect 26256 57863 26328 57939
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56608 575 56684
rect 629 56608 701 56684
rect 749 56608 821 56684
rect 503 56490 575 56566
rect 629 56490 701 56566
rect 749 56490 821 56566
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55405 575 55481
rect 629 55405 701 55481
rect 749 55405 821 55481
rect 503 55287 575 55363
rect 629 55287 701 55363
rect 749 55287 821 55363
rect 25068 55470 25140 55546
rect 25194 55470 25266 55546
rect 25314 55470 25386 55546
rect 25068 55352 25140 55428
rect 25194 55352 25266 55428
rect 25314 55352 25386 55428
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 54020 26082 54096
rect 26136 54020 26208 54096
rect 26256 54020 26328 54096
rect 26010 53902 26082 53978
rect 26136 53902 26208 53978
rect 26256 53902 26328 53978
rect 504 53223 576 53299
rect 626 53223 698 53299
rect 752 53223 824 53299
rect 504 53076 576 53152
rect 626 53076 698 53152
rect 752 53076 824 53152
rect 504 52939 576 53015
rect 626 52939 698 53015
rect 752 52939 824 53015
rect 503 52628 575 52704
rect 629 52628 701 52704
rect 749 52628 821 52704
rect 503 52510 575 52586
rect 629 52510 701 52586
rect 749 52510 821 52586
rect 25068 52554 25140 52630
rect 25194 52554 25266 52630
rect 25314 52554 25386 52630
rect 25068 52436 25140 52512
rect 25194 52436 25266 52512
rect 25314 52436 25386 52512
rect 503 51421 575 51497
rect 629 51421 701 51497
rect 749 51421 821 51497
rect 503 51303 575 51379
rect 629 51303 701 51379
rect 749 51303 821 51379
rect 25068 51371 25140 51447
rect 25194 51371 25266 51447
rect 25314 51371 25386 51447
rect 25068 51253 25140 51329
rect 25194 51253 25266 51329
rect 25314 51253 25386 51329
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50003 26082 50079
rect 26136 50003 26208 50079
rect 26256 50003 26328 50079
rect 26010 49885 26082 49961
rect 26136 49885 26208 49961
rect 26256 49885 26328 49961
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48655 575 48731
rect 629 48655 701 48731
rect 749 48655 821 48731
rect 503 48537 575 48613
rect 629 48537 701 48613
rect 749 48537 821 48613
rect 25068 48499 25140 48575
rect 25194 48499 25266 48575
rect 25314 48499 25386 48575
rect 25068 48381 25140 48457
rect 25194 48381 25266 48457
rect 25314 48381 25386 48457
rect 503 47468 575 47544
rect 629 47468 701 47544
rect 749 47468 821 47544
rect 503 47350 575 47426
rect 629 47350 701 47426
rect 749 47350 821 47426
rect 25068 47364 25140 47440
rect 25194 47364 25266 47440
rect 25314 47364 25386 47440
rect 25068 47246 25140 47322
rect 25194 47246 25266 47322
rect 25314 47246 25386 47322
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46082 26082 46158
rect 26136 46082 26208 46158
rect 26256 46082 26328 46158
rect 26010 45964 26082 46040
rect 26136 45964 26208 46040
rect 26256 45964 26328 46040
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44646 575 44722
rect 629 44646 701 44722
rect 749 44646 821 44722
rect 503 44528 575 44604
rect 629 44528 701 44604
rect 749 44528 821 44604
rect 25068 44605 25140 44681
rect 25194 44605 25266 44681
rect 25314 44605 25386 44681
rect 25068 44487 25140 44563
rect 25194 44487 25266 44563
rect 25314 44487 25386 44563
rect 503 43493 575 43569
rect 629 43493 701 43569
rect 749 43493 821 43569
rect 503 43375 575 43451
rect 629 43375 701 43451
rect 749 43375 821 43451
rect 25068 43452 25140 43528
rect 25194 43452 25266 43528
rect 25314 43452 25386 43528
rect 25068 43334 25140 43410
rect 25194 43334 25266 43410
rect 25314 43334 25386 43410
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 41824 26082 41900
rect 26136 41824 26208 41900
rect 26256 41824 26328 41900
rect 26010 41706 26082 41782
rect 26136 41706 26208 41782
rect 26256 41706 26328 41782
rect 504 41224 576 41300
rect 626 41224 698 41300
rect 752 41224 824 41300
rect 504 41077 576 41153
rect 626 41077 698 41153
rect 752 41077 824 41153
rect 504 40940 576 41016
rect 626 40940 698 41016
rect 752 40940 824 41016
rect 503 40433 575 40509
rect 629 40433 701 40509
rect 749 40433 821 40509
rect 503 40315 575 40391
rect 629 40315 701 40391
rect 749 40315 821 40391
rect 25068 40336 25140 40412
rect 25194 40336 25266 40412
rect 25314 40336 25386 40412
rect 25068 40218 25140 40294
rect 25194 40218 25266 40294
rect 25314 40218 25386 40294
rect 2257 35869 2313 35925
rect 2337 35869 2393 35925
rect 2257 35789 2313 35845
rect 2337 35789 2393 35845
rect 32 35661 112 35741
rect 157 35661 237 35741
rect 282 35661 362 35741
rect 32 35555 112 35635
rect 157 35555 237 35635
rect 282 35555 362 35635
rect 1416 35263 1472 35319
rect 1498 35264 1554 35320
rect 1417 35183 1473 35239
rect 1499 35184 1555 35240
rect 3361 35848 3417 35904
rect 3441 35848 3497 35904
rect 3361 35768 3417 35824
rect 3441 35768 3497 35824
rect 479 35052 561 35130
rect 593 35052 675 35130
rect 707 35052 789 35130
rect 16 34508 98 34586
rect 130 34508 212 34586
rect 244 34508 326 34586
rect 479 33964 561 34042
rect 593 33964 675 34042
rect 707 33964 789 34042
rect 16 33420 98 33498
rect 130 33420 212 33498
rect 244 33420 326 33498
rect 479 32876 561 32954
rect 593 32876 675 32954
rect 707 32876 789 32954
rect 2760 35262 2816 35318
rect 2840 35261 2896 35317
rect 2761 35181 2817 35237
rect 2841 35181 2897 35237
rect 25535 35646 25615 35726
rect 25660 35646 25740 35726
rect 25785 35646 25865 35726
rect 25534 35526 25614 35606
rect 25659 35526 25739 35606
rect 25784 35526 25864 35606
rect 3360 35261 3416 35317
rect 3440 35260 3496 35316
rect 3361 35180 3417 35236
rect 3441 35180 3497 35236
rect 25061 34892 25141 34972
rect 25186 34892 25266 34972
rect 25311 34892 25391 34972
rect 25060 34772 25140 34852
rect 25185 34772 25265 34852
rect 25310 34772 25390 34852
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 24560 33396 24640 33476
rect 24685 33396 24765 33476
rect 24810 33396 24890 33476
rect 24559 33276 24639 33356
rect 24684 33276 24764 33356
rect 24809 33276 24889 33356
rect 25535 33396 25615 33476
rect 25660 33396 25740 33476
rect 25785 33396 25865 33476
rect 25534 33276 25614 33356
rect 25659 33276 25739 33356
rect 25784 33276 25864 33356
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 2544 32401 2600 32463
rect 2624 32401 2680 32463
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 25060 31837 25140 31917
rect 25185 31837 25265 31917
rect 25310 31837 25390 31917
rect 25059 31717 25139 31797
rect 25184 31717 25264 31797
rect 25309 31717 25389 31797
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal3 >>
rect 25026 67492 25426 67517
rect 463 67452 864 67477
rect 463 67376 503 67452
rect 575 67376 629 67452
rect 701 67376 749 67452
rect 821 67376 864 67452
rect 463 67334 864 67376
rect 463 67258 503 67334
rect 575 67258 629 67334
rect 701 67258 749 67334
rect 821 67258 864 67334
rect 25026 67416 25068 67492
rect 25140 67416 25194 67492
rect 25266 67416 25314 67492
rect 25386 67416 25426 67492
rect 25026 67374 25426 67416
rect 25026 67298 25068 67374
rect 25140 67298 25194 67374
rect 25266 67298 25314 67374
rect 25386 67298 25426 67374
rect 25026 67262 25426 67298
rect 463 67222 864 67258
rect 463 67060 863 67109
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 66650 863 66700
rect 25970 66071 26370 66096
rect 25970 65995 26010 66071
rect 26082 65995 26136 66071
rect 26208 65995 26256 66071
rect 26328 65995 26370 66071
rect 25970 65953 26370 65995
rect 25970 65877 26010 65953
rect 26082 65877 26136 65953
rect 26208 65877 26256 65953
rect 26328 65877 26370 65953
rect 25970 65841 26370 65877
rect 463 65300 863 65349
rect 463 65224 504 65300
rect 576 65224 626 65300
rect 698 65224 752 65300
rect 824 65224 863 65300
rect 463 65153 863 65224
rect 463 65077 504 65153
rect 576 65077 626 65153
rect 698 65077 752 65153
rect 824 65077 863 65153
rect 463 65016 863 65077
rect 463 64940 504 65016
rect 576 64940 626 65016
rect 698 64940 752 65016
rect 824 64940 863 65016
rect 463 64890 863 64940
rect 463 64779 864 64804
rect 463 64703 503 64779
rect 575 64703 629 64779
rect 701 64703 749 64779
rect 821 64703 864 64779
rect 463 64661 864 64703
rect 463 64585 503 64661
rect 575 64585 629 64661
rect 701 64585 749 64661
rect 821 64585 864 64661
rect 463 64549 864 64585
rect 25028 64695 25428 64720
rect 25028 64619 25068 64695
rect 25140 64619 25194 64695
rect 25266 64619 25314 64695
rect 25386 64619 25428 64695
rect 25028 64577 25428 64619
rect 25028 64501 25068 64577
rect 25140 64501 25194 64577
rect 25266 64501 25314 64577
rect 25386 64501 25428 64577
rect 25028 64465 25428 64501
rect 25026 63492 25426 63517
rect 463 63450 864 63475
rect 463 63374 503 63450
rect 575 63374 629 63450
rect 701 63374 749 63450
rect 821 63374 864 63450
rect 463 63332 864 63374
rect 463 63256 503 63332
rect 575 63256 629 63332
rect 701 63256 749 63332
rect 821 63256 864 63332
rect 25026 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25426 63492
rect 25026 63374 25426 63416
rect 25026 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25426 63374
rect 25026 63262 25426 63298
rect 463 63220 864 63256
rect 463 63060 863 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 62650 863 62700
rect 25970 62058 26370 62083
rect 25970 61982 26010 62058
rect 26082 61982 26136 62058
rect 26208 61982 26256 62058
rect 26328 61982 26370 62058
rect 25970 61940 26370 61982
rect 25970 61864 26010 61940
rect 26082 61864 26136 61940
rect 26208 61864 26256 61940
rect 26328 61864 26370 61940
rect 25970 61828 26370 61864
rect 463 61301 863 61350
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60891 863 60941
rect 463 60710 864 60735
rect 463 60634 503 60710
rect 575 60634 629 60710
rect 701 60634 749 60710
rect 821 60634 864 60710
rect 463 60592 864 60634
rect 463 60516 503 60592
rect 575 60516 629 60592
rect 701 60516 749 60592
rect 821 60516 864 60592
rect 463 60480 864 60516
rect 25028 60695 25428 60720
rect 25028 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 25028 60577 25428 60619
rect 25028 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 25028 60465 25428 60501
rect 463 59532 864 59557
rect 463 59456 503 59532
rect 575 59456 629 59532
rect 701 59456 749 59532
rect 821 59456 864 59532
rect 463 59414 864 59456
rect 463 59338 503 59414
rect 575 59338 629 59414
rect 701 59338 749 59414
rect 821 59338 864 59414
rect 463 59302 864 59338
rect 25026 59492 25426 59517
rect 25026 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25426 59492
rect 25026 59374 25426 59416
rect 25026 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25426 59374
rect 25026 59262 25426 59298
rect 464 59068 864 59109
rect 463 59060 864 59068
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 25970 58057 26370 58082
rect 25970 57981 26010 58057
rect 26082 57981 26136 58057
rect 26208 57981 26256 58057
rect 26328 57981 26370 58057
rect 25970 57939 26370 57981
rect 25970 57863 26010 57939
rect 26082 57863 26136 57939
rect 26208 57863 26256 57939
rect 26328 57863 26370 57939
rect 25970 57827 26370 57863
rect 463 57301 863 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56891 863 56941
rect 463 56684 866 56709
rect 463 56608 503 56684
rect 575 56608 629 56684
rect 701 56608 749 56684
rect 821 56608 866 56684
rect 463 56566 866 56608
rect 463 56490 503 56566
rect 575 56490 629 56566
rect 701 56490 749 56566
rect 821 56490 866 56566
rect 463 56454 866 56490
rect 25028 56695 25428 56720
rect 25028 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 25028 56577 25428 56619
rect 25028 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 25028 56465 25428 56501
rect 25027 55546 25427 55571
rect 463 55481 864 55506
rect 463 55405 503 55481
rect 575 55405 629 55481
rect 701 55405 749 55481
rect 821 55405 864 55481
rect 463 55363 864 55405
rect 463 55287 503 55363
rect 575 55287 629 55363
rect 701 55287 749 55363
rect 821 55287 864 55363
rect 25027 55470 25068 55546
rect 25140 55470 25194 55546
rect 25266 55470 25314 55546
rect 25386 55470 25427 55546
rect 25027 55428 25427 55470
rect 25027 55352 25068 55428
rect 25140 55352 25194 55428
rect 25266 55352 25314 55428
rect 25386 55352 25427 55428
rect 25027 55316 25427 55352
rect 463 55251 864 55287
rect 464 55068 864 55109
rect 463 55060 864 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 25970 54096 26370 54121
rect 25970 54020 26010 54096
rect 26082 54020 26136 54096
rect 26208 54020 26256 54096
rect 26328 54020 26370 54096
rect 25970 53978 26370 54020
rect 25970 53902 26010 53978
rect 26082 53902 26136 53978
rect 26208 53902 26256 53978
rect 26328 53902 26370 53978
rect 25970 53866 26370 53902
rect 463 53299 863 53348
rect 463 53223 504 53299
rect 576 53223 626 53299
rect 698 53223 752 53299
rect 824 53223 863 53299
rect 463 53152 863 53223
rect 463 53076 504 53152
rect 576 53076 626 53152
rect 698 53076 752 53152
rect 824 53076 863 53152
rect 463 53015 863 53076
rect 463 52939 504 53015
rect 576 52939 626 53015
rect 698 52939 752 53015
rect 824 52939 863 53015
rect 463 52889 863 52939
rect 463 52704 864 52729
rect 463 52628 503 52704
rect 575 52628 629 52704
rect 701 52628 749 52704
rect 821 52628 864 52704
rect 463 52586 864 52628
rect 463 52510 503 52586
rect 575 52510 629 52586
rect 701 52510 749 52586
rect 821 52510 864 52586
rect 463 52474 864 52510
rect 25028 52630 25428 52655
rect 25028 52554 25068 52630
rect 25140 52554 25194 52630
rect 25266 52554 25314 52630
rect 25386 52554 25428 52630
rect 25028 52512 25428 52554
rect 25028 52436 25068 52512
rect 25140 52436 25194 52512
rect 25266 52436 25314 52512
rect 25386 52436 25428 52512
rect 25028 52400 25428 52436
rect 463 51497 866 51522
rect 463 51421 503 51497
rect 575 51421 629 51497
rect 701 51421 749 51497
rect 821 51421 866 51497
rect 463 51379 866 51421
rect 463 51303 503 51379
rect 575 51303 629 51379
rect 701 51303 749 51379
rect 821 51303 866 51379
rect 463 51267 866 51303
rect 25027 51447 25427 51472
rect 25027 51371 25068 51447
rect 25140 51371 25194 51447
rect 25266 51371 25314 51447
rect 25386 51371 25427 51447
rect 25027 51329 25427 51371
rect 25027 51253 25068 51329
rect 25140 51253 25194 51329
rect 25266 51253 25314 51329
rect 25386 51253 25427 51329
rect 25027 51217 25427 51253
rect 463 51060 863 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 50650 863 50700
rect 25970 50079 26370 50104
rect 25970 50003 26010 50079
rect 26082 50003 26136 50079
rect 26208 50003 26256 50079
rect 26328 50003 26370 50079
rect 25970 49961 26370 50003
rect 25970 49885 26010 49961
rect 26082 49885 26136 49961
rect 26208 49885 26256 49961
rect 26328 49885 26370 49961
rect 25970 49849 26370 49885
rect 463 49301 863 49350
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48891 863 48941
rect 463 48731 864 48756
rect 463 48655 503 48731
rect 575 48655 629 48731
rect 701 48655 749 48731
rect 821 48655 864 48731
rect 463 48613 864 48655
rect 463 48537 503 48613
rect 575 48537 629 48613
rect 701 48537 749 48613
rect 821 48537 864 48613
rect 463 48501 864 48537
rect 25028 48575 25428 48600
rect 25028 48499 25068 48575
rect 25140 48499 25194 48575
rect 25266 48499 25314 48575
rect 25386 48499 25428 48575
rect 25028 48457 25428 48499
rect 25028 48381 25068 48457
rect 25140 48381 25194 48457
rect 25266 48381 25314 48457
rect 25386 48381 25428 48457
rect 25028 48345 25428 48381
rect 463 47544 864 47569
rect 463 47468 503 47544
rect 575 47468 629 47544
rect 701 47468 749 47544
rect 821 47468 864 47544
rect 463 47426 864 47468
rect 463 47350 503 47426
rect 575 47350 629 47426
rect 701 47350 749 47426
rect 821 47350 864 47426
rect 463 47314 864 47350
rect 25028 47440 25428 47465
rect 25028 47364 25068 47440
rect 25140 47364 25194 47440
rect 25266 47364 25314 47440
rect 25386 47364 25428 47440
rect 25028 47322 25428 47364
rect 25028 47246 25068 47322
rect 25140 47246 25194 47322
rect 25266 47246 25314 47322
rect 25386 47246 25428 47322
rect 25028 47210 25428 47246
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 25970 46158 26370 46183
rect 25970 46082 26010 46158
rect 26082 46082 26136 46158
rect 26208 46082 26256 46158
rect 26328 46082 26370 46158
rect 25970 46040 26370 46082
rect 25970 45964 26010 46040
rect 26082 45964 26136 46040
rect 26208 45964 26256 46040
rect 26328 45964 26370 46040
rect 25970 45928 26370 45964
rect 463 45301 863 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44891 863 44941
rect 463 44722 864 44747
rect 463 44646 503 44722
rect 575 44646 629 44722
rect 701 44646 749 44722
rect 821 44646 864 44722
rect 463 44604 864 44646
rect 463 44528 503 44604
rect 575 44528 629 44604
rect 701 44528 749 44604
rect 821 44528 864 44604
rect 463 44492 864 44528
rect 25028 44681 25428 44706
rect 25028 44605 25068 44681
rect 25140 44605 25194 44681
rect 25266 44605 25314 44681
rect 25386 44605 25428 44681
rect 25028 44563 25428 44605
rect 25028 44487 25068 44563
rect 25140 44487 25194 44563
rect 25266 44487 25314 44563
rect 25386 44487 25428 44563
rect 25028 44451 25428 44487
rect 463 43569 864 43594
rect 463 43493 503 43569
rect 575 43493 629 43569
rect 701 43493 749 43569
rect 821 43493 864 43569
rect 463 43451 864 43493
rect 463 43375 503 43451
rect 575 43375 629 43451
rect 701 43375 749 43451
rect 821 43375 864 43451
rect 463 43339 864 43375
rect 25028 43528 25428 43553
rect 25028 43452 25068 43528
rect 25140 43452 25194 43528
rect 25266 43452 25314 43528
rect 25386 43452 25428 43528
rect 25028 43410 25428 43452
rect 25028 43334 25068 43410
rect 25140 43334 25194 43410
rect 25266 43334 25314 43410
rect 25386 43334 25428 43410
rect 25028 43298 25428 43334
rect 463 43060 863 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 42650 863 42700
rect 25970 41900 26370 41925
rect 25970 41824 26010 41900
rect 26082 41824 26136 41900
rect 26208 41824 26256 41900
rect 26328 41824 26370 41900
rect 25970 41782 26370 41824
rect 25970 41706 26010 41782
rect 26082 41706 26136 41782
rect 26208 41706 26256 41782
rect 26328 41706 26370 41782
rect 25970 41670 26370 41706
rect 463 41300 863 41350
rect 463 41224 504 41300
rect 576 41224 626 41300
rect 698 41224 752 41300
rect 824 41224 863 41300
rect 463 41153 863 41224
rect 463 41077 504 41153
rect 576 41077 626 41153
rect 698 41077 752 41153
rect 824 41077 863 41153
rect 463 41016 863 41077
rect 463 40940 504 41016
rect 576 40940 626 41016
rect 698 40940 752 41016
rect 824 40940 863 41016
rect 463 40891 863 40940
rect 463 40890 836 40891
rect 463 40509 863 40534
rect 463 40433 503 40509
rect 575 40433 629 40509
rect 701 40433 749 40509
rect 821 40433 863 40509
rect 463 40391 863 40433
rect 463 40315 503 40391
rect 575 40315 629 40391
rect 701 40315 749 40391
rect 821 40315 863 40391
rect 463 40279 863 40315
rect 25028 40412 25428 40437
rect 25028 40336 25068 40412
rect 25140 40336 25194 40412
rect 25266 40336 25314 40412
rect 25386 40336 25428 40412
rect 25028 40294 25428 40336
rect 25028 40218 25068 40294
rect 25140 40218 25194 40294
rect 25266 40218 25314 40294
rect 25386 40218 25428 40294
rect 25028 40182 25428 40218
rect 2248 35925 2401 35940
rect 2248 35861 2249 35925
rect 2313 35861 2337 35925
rect 2248 35845 2401 35861
rect 2248 35781 2249 35845
rect 2313 35781 2337 35845
rect 2248 35775 2401 35781
rect 3352 35905 4345 35920
rect 3352 35904 4192 35905
rect 3352 35848 3361 35904
rect 3417 35848 3441 35904
rect 3497 35848 4192 35904
rect 3352 35841 4192 35848
rect 4256 35841 4280 35905
rect 4344 35841 4345 35905
rect 3352 35825 4345 35841
rect 3352 35824 4192 35825
rect 3352 35768 3361 35824
rect 3417 35768 3441 35824
rect 3497 35768 4192 35824
rect 3352 35761 4192 35768
rect 4256 35761 4280 35825
rect 4344 35761 4345 35825
rect 3352 35754 4345 35761
rect 0 35741 400 35752
rect 0 35661 32 35741
rect 112 35661 156 35741
rect 237 35661 282 35741
rect 362 35661 400 35741
rect 0 35635 400 35661
rect 0 35555 32 35635
rect 112 35555 156 35635
rect 237 35555 282 35635
rect 362 35555 400 35635
rect 0 35528 400 35555
rect 25502 35726 25902 35752
rect 25502 35646 25535 35726
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 25502 35606 25902 35646
rect 25502 35526 25534 35606
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 25502 35497 25902 35526
rect 2689 35333 3502 35334
rect 1411 35320 3502 35333
rect 1411 35319 1498 35320
rect 1411 35263 1416 35319
rect 1472 35264 1498 35319
rect 1554 35318 3502 35320
rect 1554 35264 2760 35318
rect 1472 35263 2760 35264
rect 1411 35262 2760 35263
rect 2816 35317 3502 35318
rect 2816 35262 2840 35317
rect 1411 35261 2840 35262
rect 2896 35261 3360 35317
rect 3416 35316 3502 35317
rect 3416 35261 3440 35316
rect 1411 35260 3440 35261
rect 3496 35260 3502 35316
rect 1411 35240 3502 35260
rect 1411 35239 1499 35240
rect 1411 35183 1417 35239
rect 1473 35184 1499 35239
rect 1555 35237 3502 35240
rect 1555 35184 2761 35237
rect 1473 35183 2761 35184
rect 1411 35181 2761 35183
rect 2817 35181 2841 35237
rect 2897 35236 3502 35237
rect 2897 35181 3361 35236
rect 1411 35180 3361 35181
rect 3417 35180 3441 35236
rect 3497 35180 3502 35236
rect 1411 35169 3502 35180
rect 463 35131 805 35139
rect 463 35051 478 35131
rect 562 35051 592 35131
rect 676 35051 706 35131
rect 790 35051 805 35131
rect 463 35043 805 35051
rect 25028 34972 25428 34998
rect 25028 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 25028 34852 25428 34892
rect 25028 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 25028 34743 25428 34772
rect 0 34587 342 34595
rect 0 34507 15 34587
rect 99 34507 129 34587
rect 213 34507 243 34587
rect 327 34507 342 34587
rect 0 34499 342 34507
rect 25028 34392 25428 34442
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 25028 34245 25428 34316
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 463 34043 805 34051
rect 463 33963 478 34043
rect 562 33963 592 34043
rect 676 33963 706 34043
rect 790 33963 805 34043
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 25028 33983 25428 34032
rect 25028 33982 25401 33983
rect 463 33955 805 33963
rect 0 33499 342 33507
rect 0 33419 15 33499
rect 99 33419 129 33499
rect 213 33419 243 33499
rect 327 33419 342 33499
rect 0 33411 342 33419
rect 24527 33476 24927 33502
rect 24527 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 24927 33476
rect 24527 33356 24927 33396
rect 24527 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 24927 33356
rect 24527 33247 24927 33276
rect 25502 33476 25902 33502
rect 25502 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 25502 33356 25902 33396
rect 25502 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 25502 33247 25902 33276
rect 463 32955 805 32963
rect 463 32875 478 32955
rect 562 32875 592 32955
rect 676 32875 706 32955
rect 790 32875 805 32955
rect 463 32867 805 32875
rect 25028 32632 25428 32682
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 2535 32475 2688 32476
rect 2535 32463 2689 32475
rect 2535 32399 2536 32463
rect 2600 32399 2624 32463
rect 2688 32399 2689 32463
rect 2535 32391 2689 32399
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 32223 25428 32272
rect 25028 32222 25401 32223
rect 25027 31917 25427 31943
rect 25027 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25427 31917
rect 25027 31797 25427 31837
rect 25027 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25427 31797
rect 25027 31688 25427 31717
rect 463 28302 866 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 866 28302
rect 463 28184 866 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 866 28184
rect 463 28072 866 28108
rect 25025 28302 25428 28360
rect 25025 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 25025 28184 25428 28226
rect 25025 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 25025 28072 25428 28108
rect 463 27520 863 27545
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 863 27520
rect 463 27402 863 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 863 27402
rect 463 27290 863 27326
rect 25028 27520 25428 27545
rect 25028 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 25028 27402 25428 27444
rect 25028 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 25028 27290 25428 27326
rect 463 27061 863 27111
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 26651 863 26701
rect 25970 26130 26370 26155
rect 25970 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 25970 26012 26370 26054
rect 25970 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 25970 25900 26370 25936
rect 463 25294 863 25349
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24884 862 24885
rect 463 24608 863 24633
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 863 24608
rect 463 24490 863 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 863 24490
rect 463 24378 863 24414
rect 25028 24559 25428 24584
rect 25028 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 25028 24441 25428 24483
rect 25028 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 25028 24329 25428 24365
rect 463 23604 863 23629
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 863 23604
rect 463 23486 863 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 863 23486
rect 463 23374 863 23410
rect 25027 23442 25427 23467
rect 25027 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25427 23442
rect 25027 23324 25427 23366
rect 25027 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25427 23324
rect 25027 23212 25427 23248
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 25970 21971 26370 21996
rect 25970 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 25970 21853 26370 21895
rect 25970 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 25970 21741 26370 21777
rect 463 21300 863 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20890 863 20940
rect 463 20626 864 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 864 20626
rect 463 20508 864 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 864 20508
rect 463 20396 864 20432
rect 25028 20599 25428 20624
rect 25028 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 25028 20481 25428 20523
rect 25028 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 25028 20369 25428 20405
rect 463 19544 864 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 864 19544
rect 463 19426 864 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 864 19426
rect 463 19314 864 19350
rect 25028 19424 25428 19449
rect 25028 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 25028 19306 25428 19348
rect 25028 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 25028 19194 25428 19230
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 25970 18181 26370 18206
rect 25970 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 25970 18063 26370 18105
rect 25970 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 25970 17951 26370 17987
rect 463 17301 863 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16891 863 16941
rect 463 16669 864 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 864 16669
rect 463 16551 864 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 864 16551
rect 463 16439 864 16475
rect 25027 16583 25427 16608
rect 25027 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25427 16583
rect 25027 16465 25427 16507
rect 25027 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25427 16465
rect 25027 16353 25427 16389
rect 463 15568 864 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 864 15568
rect 463 15450 864 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 864 15450
rect 463 15338 864 15374
rect 25027 15412 25427 15437
rect 25027 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25427 15412
rect 25027 15294 25427 15336
rect 25027 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25427 15294
rect 25027 15182 25427 15218
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 25970 14074 26370 14099
rect 25970 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 25970 13956 26370 13998
rect 25970 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 25970 13844 26370 13880
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12702 865 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 865 12702
rect 463 12584 865 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 865 12584
rect 463 12472 865 12508
rect 25027 12651 25427 12676
rect 25027 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25427 12651
rect 25027 12533 25427 12575
rect 25027 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25427 12533
rect 25027 12421 25427 12457
rect 463 11486 866 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 866 11486
rect 463 11368 866 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 866 11368
rect 463 11256 866 11292
rect 25027 11437 25427 11462
rect 25027 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25427 11437
rect 25027 11319 25427 11361
rect 25027 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25427 11319
rect 25027 11207 25427 11243
rect 463 11060 863 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 10650 863 10700
rect 25970 10256 26370 10281
rect 25970 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 25970 10138 26370 10180
rect 25970 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 25970 10026 26370 10062
rect 463 9300 863 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8890 863 8940
rect 463 8621 864 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 864 8621
rect 463 8503 864 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 864 8503
rect 463 8391 864 8427
rect 25028 8594 25428 8619
rect 25028 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 25028 8476 25428 8518
rect 25028 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 25028 8364 25428 8400
rect 463 7499 864 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 864 7499
rect 463 7381 864 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 864 7381
rect 463 7269 864 7305
rect 25027 7437 25427 7462
rect 25027 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25427 7437
rect 25027 7319 25427 7361
rect 25027 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25427 7319
rect 25027 7207 25427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 25970 6292 26370 6317
rect 25970 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 25970 6174 26370 6216
rect 25970 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 25970 6062 26370 6098
rect 463 5299 863 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4889 863 4939
rect 463 4639 863 4664
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 863 4639
rect 463 4521 863 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 863 4521
rect 463 4409 863 4445
rect 25028 4594 25428 4619
rect 25028 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 25028 4476 25428 4518
rect 25028 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 25028 4364 25428 4400
rect 463 3528 863 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3298 863 3334
rect 25027 3437 25427 3462
rect 25027 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25427 3437
rect 25027 3319 25427 3361
rect 25027 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25427 3319
rect 25027 3207 25427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 25970 2280 26370 2305
rect 25970 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 25970 2162 26370 2204
rect 25970 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 25970 2050 26370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 25028 594 25428 619
rect 25028 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 25028 476 25428 518
rect 25028 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 25028 364 25428 400
<< via3 >>
rect 503 67376 575 67452
rect 629 67376 701 67452
rect 749 67376 821 67452
rect 503 67258 575 67334
rect 629 67258 701 67334
rect 749 67258 821 67334
rect 25068 67416 25140 67492
rect 25194 67416 25266 67492
rect 25314 67416 25386 67492
rect 25068 67298 25140 67374
rect 25194 67298 25266 67374
rect 25314 67298 25386 67374
rect 504 66984 576 67060
rect 626 66984 698 67060
rect 752 66984 824 67060
rect 504 66837 576 66913
rect 626 66837 698 66913
rect 752 66837 824 66913
rect 504 66700 576 66776
rect 626 66700 698 66776
rect 752 66700 824 66776
rect 26010 65995 26082 66071
rect 26136 65995 26208 66071
rect 26256 65995 26328 66071
rect 26010 65877 26082 65953
rect 26136 65877 26208 65953
rect 26256 65877 26328 65953
rect 504 65224 576 65300
rect 626 65224 698 65300
rect 752 65224 824 65300
rect 504 65077 576 65153
rect 626 65077 698 65153
rect 752 65077 824 65153
rect 504 64940 576 65016
rect 626 64940 698 65016
rect 752 64940 824 65016
rect 503 64703 575 64779
rect 629 64703 701 64779
rect 749 64703 821 64779
rect 503 64585 575 64661
rect 629 64585 701 64661
rect 749 64585 821 64661
rect 25068 64619 25140 64695
rect 25194 64619 25266 64695
rect 25314 64619 25386 64695
rect 25068 64501 25140 64577
rect 25194 64501 25266 64577
rect 25314 64501 25386 64577
rect 503 63374 575 63450
rect 629 63374 701 63450
rect 749 63374 821 63450
rect 503 63256 575 63332
rect 629 63256 701 63332
rect 749 63256 821 63332
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61982 26082 62058
rect 26136 61982 26208 62058
rect 26256 61982 26328 62058
rect 26010 61864 26082 61940
rect 26136 61864 26208 61940
rect 26256 61864 26328 61940
rect 504 61225 576 61301
rect 626 61225 698 61301
rect 752 61225 824 61301
rect 504 61078 576 61154
rect 626 61078 698 61154
rect 752 61078 824 61154
rect 504 60941 576 61017
rect 626 60941 698 61017
rect 752 60941 824 61017
rect 503 60634 575 60710
rect 629 60634 701 60710
rect 749 60634 821 60710
rect 503 60516 575 60592
rect 629 60516 701 60592
rect 749 60516 821 60592
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59456 575 59532
rect 629 59456 701 59532
rect 749 59456 821 59532
rect 503 59338 575 59414
rect 629 59338 701 59414
rect 749 59338 821 59414
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57981 26082 58057
rect 26136 57981 26208 58057
rect 26256 57981 26328 58057
rect 26010 57863 26082 57939
rect 26136 57863 26208 57939
rect 26256 57863 26328 57939
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56608 575 56684
rect 629 56608 701 56684
rect 749 56608 821 56684
rect 503 56490 575 56566
rect 629 56490 701 56566
rect 749 56490 821 56566
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55405 575 55481
rect 629 55405 701 55481
rect 749 55405 821 55481
rect 503 55287 575 55363
rect 629 55287 701 55363
rect 749 55287 821 55363
rect 25068 55470 25140 55546
rect 25194 55470 25266 55546
rect 25314 55470 25386 55546
rect 25068 55352 25140 55428
rect 25194 55352 25266 55428
rect 25314 55352 25386 55428
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 54020 26082 54096
rect 26136 54020 26208 54096
rect 26256 54020 26328 54096
rect 26010 53902 26082 53978
rect 26136 53902 26208 53978
rect 26256 53902 26328 53978
rect 504 53223 576 53299
rect 626 53223 698 53299
rect 752 53223 824 53299
rect 504 53076 576 53152
rect 626 53076 698 53152
rect 752 53076 824 53152
rect 504 52939 576 53015
rect 626 52939 698 53015
rect 752 52939 824 53015
rect 503 52628 575 52704
rect 629 52628 701 52704
rect 749 52628 821 52704
rect 503 52510 575 52586
rect 629 52510 701 52586
rect 749 52510 821 52586
rect 25068 52554 25140 52630
rect 25194 52554 25266 52630
rect 25314 52554 25386 52630
rect 25068 52436 25140 52512
rect 25194 52436 25266 52512
rect 25314 52436 25386 52512
rect 503 51421 575 51497
rect 629 51421 701 51497
rect 749 51421 821 51497
rect 503 51303 575 51379
rect 629 51303 701 51379
rect 749 51303 821 51379
rect 25068 51371 25140 51447
rect 25194 51371 25266 51447
rect 25314 51371 25386 51447
rect 25068 51253 25140 51329
rect 25194 51253 25266 51329
rect 25314 51253 25386 51329
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50003 26082 50079
rect 26136 50003 26208 50079
rect 26256 50003 26328 50079
rect 26010 49885 26082 49961
rect 26136 49885 26208 49961
rect 26256 49885 26328 49961
rect 504 49225 576 49301
rect 626 49225 698 49301
rect 752 49225 824 49301
rect 504 49078 576 49154
rect 626 49078 698 49154
rect 752 49078 824 49154
rect 504 48941 576 49017
rect 626 48941 698 49017
rect 752 48941 824 49017
rect 503 48655 575 48731
rect 629 48655 701 48731
rect 749 48655 821 48731
rect 503 48537 575 48613
rect 629 48537 701 48613
rect 749 48537 821 48613
rect 25068 48499 25140 48575
rect 25194 48499 25266 48575
rect 25314 48499 25386 48575
rect 25068 48381 25140 48457
rect 25194 48381 25266 48457
rect 25314 48381 25386 48457
rect 503 47468 575 47544
rect 629 47468 701 47544
rect 749 47468 821 47544
rect 503 47350 575 47426
rect 629 47350 701 47426
rect 749 47350 821 47426
rect 25068 47364 25140 47440
rect 25194 47364 25266 47440
rect 25314 47364 25386 47440
rect 25068 47246 25140 47322
rect 25194 47246 25266 47322
rect 25314 47246 25386 47322
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46082 26082 46158
rect 26136 46082 26208 46158
rect 26256 46082 26328 46158
rect 26010 45964 26082 46040
rect 26136 45964 26208 46040
rect 26256 45964 26328 46040
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44646 575 44722
rect 629 44646 701 44722
rect 749 44646 821 44722
rect 503 44528 575 44604
rect 629 44528 701 44604
rect 749 44528 821 44604
rect 25068 44605 25140 44681
rect 25194 44605 25266 44681
rect 25314 44605 25386 44681
rect 25068 44487 25140 44563
rect 25194 44487 25266 44563
rect 25314 44487 25386 44563
rect 503 43493 575 43569
rect 629 43493 701 43569
rect 749 43493 821 43569
rect 503 43375 575 43451
rect 629 43375 701 43451
rect 749 43375 821 43451
rect 25068 43452 25140 43528
rect 25194 43452 25266 43528
rect 25314 43452 25386 43528
rect 25068 43334 25140 43410
rect 25194 43334 25266 43410
rect 25314 43334 25386 43410
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 41824 26082 41900
rect 26136 41824 26208 41900
rect 26256 41824 26328 41900
rect 26010 41706 26082 41782
rect 26136 41706 26208 41782
rect 26256 41706 26328 41782
rect 504 41224 576 41300
rect 626 41224 698 41300
rect 752 41224 824 41300
rect 504 41077 576 41153
rect 626 41077 698 41153
rect 752 41077 824 41153
rect 504 40940 576 41016
rect 626 40940 698 41016
rect 752 40940 824 41016
rect 503 40433 575 40509
rect 629 40433 701 40509
rect 749 40433 821 40509
rect 503 40315 575 40391
rect 629 40315 701 40391
rect 749 40315 821 40391
rect 25068 40336 25140 40412
rect 25194 40336 25266 40412
rect 25314 40336 25386 40412
rect 25068 40218 25140 40294
rect 25194 40218 25266 40294
rect 25314 40218 25386 40294
rect 2249 35869 2257 35925
rect 2257 35869 2313 35925
rect 2249 35861 2313 35869
rect 2337 35869 2393 35925
rect 2393 35869 2401 35925
rect 2337 35861 2401 35869
rect 2249 35789 2257 35845
rect 2257 35789 2313 35845
rect 2249 35781 2313 35789
rect 2337 35789 2393 35845
rect 2393 35789 2401 35845
rect 2337 35781 2401 35789
rect 4192 35841 4256 35905
rect 4280 35841 4344 35905
rect 4192 35761 4256 35825
rect 4280 35761 4344 35825
rect 32 35661 111 35741
rect 156 35661 157 35741
rect 157 35661 236 35741
rect 282 35661 362 35741
rect 32 35555 111 35635
rect 156 35555 157 35635
rect 157 35555 236 35635
rect 282 35555 362 35635
rect 25535 35646 25615 35726
rect 25660 35646 25740 35726
rect 25785 35646 25865 35726
rect 25534 35526 25614 35606
rect 25659 35526 25739 35606
rect 25784 35526 25864 35606
rect 478 35130 562 35131
rect 478 35052 479 35130
rect 479 35052 561 35130
rect 561 35052 562 35130
rect 478 35051 562 35052
rect 592 35130 676 35131
rect 592 35052 593 35130
rect 593 35052 675 35130
rect 675 35052 676 35130
rect 592 35051 676 35052
rect 706 35130 790 35131
rect 706 35052 707 35130
rect 707 35052 789 35130
rect 789 35052 790 35130
rect 706 35051 790 35052
rect 25061 34892 25141 34972
rect 25186 34892 25266 34972
rect 25311 34892 25391 34972
rect 25060 34772 25140 34852
rect 25185 34772 25265 34852
rect 25310 34772 25390 34852
rect 15 34586 99 34587
rect 15 34508 16 34586
rect 16 34508 98 34586
rect 98 34508 99 34586
rect 15 34507 99 34508
rect 129 34586 213 34587
rect 129 34508 130 34586
rect 130 34508 212 34586
rect 212 34508 213 34586
rect 129 34507 213 34508
rect 243 34586 327 34587
rect 243 34508 244 34586
rect 244 34508 326 34586
rect 326 34508 327 34586
rect 243 34507 327 34508
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 478 34042 562 34043
rect 478 33964 479 34042
rect 479 33964 561 34042
rect 561 33964 562 34042
rect 478 33963 562 33964
rect 592 34042 676 34043
rect 592 33964 593 34042
rect 593 33964 675 34042
rect 675 33964 676 34042
rect 592 33963 676 33964
rect 706 34042 790 34043
rect 706 33964 707 34042
rect 707 33964 789 34042
rect 789 33964 790 34042
rect 706 33963 790 33964
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 15 33498 99 33499
rect 15 33420 16 33498
rect 16 33420 98 33498
rect 98 33420 99 33498
rect 15 33419 99 33420
rect 129 33498 213 33499
rect 129 33420 130 33498
rect 130 33420 212 33498
rect 212 33420 213 33498
rect 129 33419 213 33420
rect 243 33498 327 33499
rect 243 33420 244 33498
rect 244 33420 326 33498
rect 326 33420 327 33498
rect 243 33419 327 33420
rect 24560 33396 24640 33476
rect 24685 33396 24765 33476
rect 24810 33396 24890 33476
rect 24559 33276 24639 33356
rect 24684 33276 24764 33356
rect 24809 33276 24889 33356
rect 25535 33396 25615 33476
rect 25660 33396 25740 33476
rect 25785 33396 25865 33476
rect 25534 33276 25614 33356
rect 25659 33276 25739 33356
rect 25784 33276 25864 33356
rect 478 32954 562 32955
rect 478 32876 479 32954
rect 479 32876 561 32954
rect 561 32876 562 32954
rect 478 32875 562 32876
rect 592 32954 676 32955
rect 592 32876 593 32954
rect 593 32876 675 32954
rect 675 32876 676 32954
rect 592 32875 676 32876
rect 706 32954 790 32955
rect 706 32876 707 32954
rect 707 32876 789 32954
rect 789 32876 790 32954
rect 706 32875 790 32876
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 2536 32401 2544 32463
rect 2544 32401 2600 32463
rect 2536 32399 2600 32401
rect 2624 32401 2680 32463
rect 2680 32401 2688 32463
rect 2624 32399 2688 32401
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 25060 31837 25140 31917
rect 25185 31837 25265 31917
rect 25310 31837 25390 31917
rect 25059 31717 25139 31797
rect 25184 31717 25264 31797
rect 25309 31717 25389 31797
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal4 >>
rect 0 35741 400 68000
rect 0 35661 32 35741
rect 111 35661 156 35741
rect 236 35661 282 35741
rect 362 35661 400 35741
rect 0 35635 400 35661
rect 0 35555 32 35635
rect 111 35555 156 35635
rect 236 35555 282 35635
rect 362 35555 400 35635
rect 0 34587 400 35555
rect 0 34507 15 34587
rect 99 34507 129 34587
rect 213 34507 243 34587
rect 327 34507 400 34587
rect 0 33499 400 34507
rect 0 33419 15 33499
rect 99 33419 129 33499
rect 213 33419 243 33499
rect 327 33419 400 33499
rect 0 0 400 33419
rect 463 67477 863 68000
rect 25028 67517 25428 68000
rect 25026 67492 25428 67517
rect 463 67452 864 67477
rect 463 67376 503 67452
rect 575 67376 629 67452
rect 701 67376 749 67452
rect 821 67376 864 67452
rect 463 67334 864 67376
rect 463 67258 503 67334
rect 575 67258 629 67334
rect 701 67258 749 67334
rect 821 67258 864 67334
rect 25026 67416 25068 67492
rect 25140 67416 25194 67492
rect 25266 67416 25314 67492
rect 25386 67416 25428 67492
rect 25026 67374 25428 67416
rect 25026 67298 25068 67374
rect 25140 67298 25194 67374
rect 25266 67298 25314 67374
rect 25386 67298 25428 67374
rect 25026 67262 25428 67298
rect 463 67222 864 67258
rect 463 67060 863 67222
rect 463 66984 504 67060
rect 576 66984 626 67060
rect 698 66984 752 67060
rect 824 66984 863 67060
rect 463 66913 863 66984
rect 463 66837 504 66913
rect 576 66837 626 66913
rect 698 66837 752 66913
rect 824 66837 863 66913
rect 463 66776 863 66837
rect 463 66700 504 66776
rect 576 66700 626 66776
rect 698 66700 752 66776
rect 824 66700 863 66776
rect 463 65300 863 66700
rect 463 65224 504 65300
rect 576 65224 626 65300
rect 698 65224 752 65300
rect 824 65224 863 65300
rect 463 65153 863 65224
rect 463 65077 504 65153
rect 576 65077 626 65153
rect 698 65077 752 65153
rect 824 65077 863 65153
rect 463 65016 863 65077
rect 463 64940 504 65016
rect 576 64940 626 65016
rect 698 64940 752 65016
rect 824 64940 863 65016
rect 463 64804 863 64940
rect 463 64779 864 64804
rect 463 64703 503 64779
rect 575 64703 629 64779
rect 701 64703 749 64779
rect 821 64703 864 64779
rect 463 64661 864 64703
rect 463 64585 503 64661
rect 575 64585 629 64661
rect 701 64585 749 64661
rect 821 64585 864 64661
rect 463 64549 864 64585
rect 25028 64695 25428 67262
rect 25028 64619 25068 64695
rect 25140 64619 25194 64695
rect 25266 64619 25314 64695
rect 25386 64619 25428 64695
rect 25028 64577 25428 64619
rect 463 63475 863 64549
rect 25028 64501 25068 64577
rect 25140 64501 25194 64577
rect 25266 64501 25314 64577
rect 25386 64501 25428 64577
rect 25028 63517 25428 64501
rect 25026 63492 25428 63517
rect 463 63450 864 63475
rect 463 63374 503 63450
rect 575 63374 629 63450
rect 701 63374 749 63450
rect 821 63374 864 63450
rect 463 63332 864 63374
rect 463 63256 503 63332
rect 575 63256 629 63332
rect 701 63256 749 63332
rect 821 63256 864 63332
rect 25026 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25428 63492
rect 25026 63374 25428 63416
rect 25026 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25428 63374
rect 25026 63262 25428 63298
rect 463 63220 864 63256
rect 463 63060 863 63220
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 61301 863 62700
rect 463 61225 504 61301
rect 576 61225 626 61301
rect 698 61225 752 61301
rect 824 61225 863 61301
rect 463 61154 863 61225
rect 463 61078 504 61154
rect 576 61078 626 61154
rect 698 61078 752 61154
rect 824 61078 863 61154
rect 463 61017 863 61078
rect 463 60941 504 61017
rect 576 60941 626 61017
rect 698 60941 752 61017
rect 824 60941 863 61017
rect 463 60735 863 60941
rect 463 60710 864 60735
rect 463 60634 503 60710
rect 575 60634 629 60710
rect 701 60634 749 60710
rect 821 60634 864 60710
rect 463 60592 864 60634
rect 463 60516 503 60592
rect 575 60516 629 60592
rect 701 60516 749 60592
rect 821 60516 864 60592
rect 463 60480 864 60516
rect 25028 60695 25428 63262
rect 25028 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 25028 60577 25428 60619
rect 25028 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 463 59557 863 60480
rect 463 59532 864 59557
rect 463 59456 503 59532
rect 575 59456 629 59532
rect 701 59456 749 59532
rect 821 59456 864 59532
rect 25028 59517 25428 60501
rect 463 59414 864 59456
rect 463 59338 503 59414
rect 575 59338 629 59414
rect 701 59338 749 59414
rect 821 59338 864 59414
rect 463 59302 864 59338
rect 25026 59492 25428 59517
rect 25026 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25428 59492
rect 25026 59374 25428 59416
rect 463 59109 863 59302
rect 25026 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25428 59374
rect 25026 59262 25428 59298
rect 463 59060 864 59109
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 864 59060
rect 463 58913 864 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 864 58913
rect 463 58776 864 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 864 58776
rect 463 58650 864 58700
rect 463 57301 863 58650
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56709 863 56941
rect 463 56684 866 56709
rect 463 56608 503 56684
rect 575 56608 629 56684
rect 701 56608 749 56684
rect 821 56608 866 56684
rect 463 56566 866 56608
rect 463 56490 503 56566
rect 575 56490 629 56566
rect 701 56490 749 56566
rect 821 56490 866 56566
rect 463 56454 866 56490
rect 25028 56695 25428 59262
rect 25028 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 25028 56577 25428 56619
rect 25028 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 463 55506 863 56454
rect 25028 55571 25428 56501
rect 25027 55546 25428 55571
rect 463 55481 864 55506
rect 463 55405 503 55481
rect 575 55405 629 55481
rect 701 55405 749 55481
rect 821 55405 864 55481
rect 463 55363 864 55405
rect 463 55287 503 55363
rect 575 55287 629 55363
rect 701 55287 749 55363
rect 821 55287 864 55363
rect 25027 55470 25068 55546
rect 25140 55470 25194 55546
rect 25266 55470 25314 55546
rect 25386 55470 25428 55546
rect 25027 55428 25428 55470
rect 25027 55352 25068 55428
rect 25140 55352 25194 55428
rect 25266 55352 25314 55428
rect 25386 55352 25428 55428
rect 25027 55316 25428 55352
rect 463 55251 864 55287
rect 463 55109 863 55251
rect 463 55060 864 55109
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 463 53299 863 54650
rect 463 53223 504 53299
rect 576 53223 626 53299
rect 698 53223 752 53299
rect 824 53223 863 53299
rect 463 53152 863 53223
rect 463 53076 504 53152
rect 576 53076 626 53152
rect 698 53076 752 53152
rect 824 53076 863 53152
rect 463 53015 863 53076
rect 463 52939 504 53015
rect 576 52939 626 53015
rect 698 52939 752 53015
rect 824 52939 863 53015
rect 463 52729 863 52939
rect 463 52704 864 52729
rect 463 52628 503 52704
rect 575 52628 629 52704
rect 701 52628 749 52704
rect 821 52628 864 52704
rect 463 52586 864 52628
rect 463 52510 503 52586
rect 575 52510 629 52586
rect 701 52510 749 52586
rect 821 52510 864 52586
rect 463 52474 864 52510
rect 25028 52630 25428 55316
rect 25028 52554 25068 52630
rect 25140 52554 25194 52630
rect 25266 52554 25314 52630
rect 25386 52554 25428 52630
rect 25028 52512 25428 52554
rect 463 51522 863 52474
rect 25028 52436 25068 52512
rect 25140 52436 25194 52512
rect 25266 52436 25314 52512
rect 25386 52436 25428 52512
rect 463 51497 866 51522
rect 463 51421 503 51497
rect 575 51421 629 51497
rect 701 51421 749 51497
rect 821 51421 866 51497
rect 25028 51472 25428 52436
rect 463 51379 866 51421
rect 463 51303 503 51379
rect 575 51303 629 51379
rect 701 51303 749 51379
rect 821 51303 866 51379
rect 463 51267 866 51303
rect 25027 51447 25428 51472
rect 25027 51371 25068 51447
rect 25140 51371 25194 51447
rect 25266 51371 25314 51447
rect 25386 51371 25428 51447
rect 25027 51329 25428 51371
rect 463 51060 863 51267
rect 25027 51253 25068 51329
rect 25140 51253 25194 51329
rect 25266 51253 25314 51329
rect 25386 51253 25428 51329
rect 25027 51217 25428 51253
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 863 51060
rect 463 50913 863 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 863 50913
rect 463 50776 863 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 863 50776
rect 463 49301 863 50700
rect 463 49225 504 49301
rect 576 49225 626 49301
rect 698 49225 752 49301
rect 824 49225 863 49301
rect 463 49154 863 49225
rect 463 49078 504 49154
rect 576 49078 626 49154
rect 698 49078 752 49154
rect 824 49078 863 49154
rect 463 49017 863 49078
rect 463 48941 504 49017
rect 576 48941 626 49017
rect 698 48941 752 49017
rect 824 48941 863 49017
rect 463 48756 863 48941
rect 463 48731 864 48756
rect 463 48655 503 48731
rect 575 48655 629 48731
rect 701 48655 749 48731
rect 821 48655 864 48731
rect 463 48613 864 48655
rect 463 48537 503 48613
rect 575 48537 629 48613
rect 701 48537 749 48613
rect 821 48537 864 48613
rect 463 48501 864 48537
rect 25028 48575 25428 51217
rect 463 47569 863 48501
rect 25028 48499 25068 48575
rect 25140 48499 25194 48575
rect 25266 48499 25314 48575
rect 25386 48499 25428 48575
rect 25028 48457 25428 48499
rect 25028 48381 25068 48457
rect 25140 48381 25194 48457
rect 25266 48381 25314 48457
rect 25386 48381 25428 48457
rect 463 47544 864 47569
rect 463 47468 503 47544
rect 575 47468 629 47544
rect 701 47468 749 47544
rect 821 47468 864 47544
rect 463 47426 864 47468
rect 463 47350 503 47426
rect 575 47350 629 47426
rect 701 47350 749 47426
rect 821 47350 864 47426
rect 463 47314 864 47350
rect 25028 47440 25428 48381
rect 25028 47364 25068 47440
rect 25140 47364 25194 47440
rect 25266 47364 25314 47440
rect 25386 47364 25428 47440
rect 25028 47322 25428 47364
rect 463 47060 863 47314
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 45301 863 46700
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44747 863 44941
rect 25028 47246 25068 47322
rect 25140 47246 25194 47322
rect 25266 47246 25314 47322
rect 25386 47246 25428 47322
rect 463 44722 864 44747
rect 463 44646 503 44722
rect 575 44646 629 44722
rect 701 44646 749 44722
rect 821 44646 864 44722
rect 463 44604 864 44646
rect 463 44528 503 44604
rect 575 44528 629 44604
rect 701 44528 749 44604
rect 821 44528 864 44604
rect 463 44492 864 44528
rect 25028 44681 25428 47246
rect 25028 44605 25068 44681
rect 25140 44605 25194 44681
rect 25266 44605 25314 44681
rect 25386 44605 25428 44681
rect 25028 44563 25428 44605
rect 463 43594 863 44492
rect 25028 44487 25068 44563
rect 25140 44487 25194 44563
rect 25266 44487 25314 44563
rect 25386 44487 25428 44563
rect 463 43569 864 43594
rect 463 43493 503 43569
rect 575 43493 629 43569
rect 701 43493 749 43569
rect 821 43493 864 43569
rect 463 43451 864 43493
rect 463 43375 503 43451
rect 575 43375 629 43451
rect 701 43375 749 43451
rect 821 43375 864 43451
rect 463 43339 864 43375
rect 25028 43528 25428 44487
rect 25028 43452 25068 43528
rect 25140 43452 25194 43528
rect 25266 43452 25314 43528
rect 25386 43452 25428 43528
rect 25028 43410 25428 43452
rect 463 43060 863 43339
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 41300 863 42700
rect 463 41224 504 41300
rect 576 41224 626 41300
rect 698 41224 752 41300
rect 824 41224 863 41300
rect 463 41153 863 41224
rect 463 41077 504 41153
rect 576 41077 626 41153
rect 698 41077 752 41153
rect 824 41077 863 41153
rect 463 41016 863 41077
rect 463 40940 504 41016
rect 576 40940 626 41016
rect 698 40940 752 41016
rect 824 40940 863 41016
rect 463 40509 863 40940
rect 463 40433 503 40509
rect 575 40433 629 40509
rect 701 40433 749 40509
rect 821 40433 863 40509
rect 463 40391 863 40433
rect 463 40315 503 40391
rect 575 40315 629 40391
rect 701 40315 749 40391
rect 821 40315 863 40391
rect 463 35131 863 40315
rect 25028 43334 25068 43410
rect 25140 43334 25194 43410
rect 25266 43334 25314 43410
rect 25386 43334 25428 43410
rect 25028 40412 25428 43334
rect 25028 40336 25068 40412
rect 25140 40336 25194 40412
rect 25266 40336 25314 40412
rect 25386 40336 25428 40412
rect 25028 40294 25428 40336
rect 25028 40218 25068 40294
rect 25140 40218 25194 40294
rect 25266 40218 25314 40294
rect 25386 40218 25428 40294
rect 2306 35942 2868 40002
rect 2246 35925 2868 35942
rect 2246 35861 2249 35925
rect 2313 35861 2337 35925
rect 2401 35861 2868 35925
rect 2246 35845 2868 35861
rect 2246 35781 2249 35845
rect 2313 35781 2337 35845
rect 2401 35781 2868 35845
rect 2246 35775 2868 35781
rect 2306 35774 2868 35775
rect 4119 35905 4490 40000
rect 4119 35841 4192 35905
rect 4256 35841 4280 35905
rect 4344 35841 4490 35905
rect 4119 35825 4490 35841
rect 4119 35761 4192 35825
rect 4256 35761 4280 35825
rect 4344 35761 4490 35825
rect 4119 35754 4490 35761
rect 463 35051 478 35131
rect 562 35051 592 35131
rect 676 35051 706 35131
rect 790 35051 863 35131
rect 463 34043 863 35051
rect 25028 34998 25428 40218
rect 24527 34972 25428 34998
rect 24527 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 24527 34852 25428 34892
rect 24527 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 24527 34743 25428 34772
rect 463 33963 478 34043
rect 562 33963 592 34043
rect 676 33963 706 34043
rect 790 33963 863 34043
rect 463 32955 863 33963
rect 25028 34392 25428 34743
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 25028 34245 25428 34316
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 24527 33476 24927 33502
rect 24527 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 24927 33476
rect 24527 33356 24927 33396
rect 24527 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 24927 33356
rect 24527 33247 24927 33276
rect 463 32875 478 32955
rect 562 32875 592 32955
rect 676 32875 706 32955
rect 790 32875 863 32955
rect 463 28360 863 32875
rect 25028 32632 25428 34032
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 2306 32463 2738 32476
rect 2306 32399 2536 32463
rect 2600 32399 2624 32463
rect 2688 32399 2738 32463
rect 463 28302 866 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 866 28302
rect 463 28184 866 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 866 28184
rect 463 28072 866 28108
rect 463 28000 863 28072
rect 2306 28000 2738 32399
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 31943 25428 32272
rect 24514 31917 25428 31943
rect 24514 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25428 31917
rect 24514 31797 25428 31837
rect 24514 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25428 31797
rect 24514 31688 25428 31717
rect 25028 28360 25428 31688
rect 25025 28302 25428 28360
rect 25025 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 25025 28184 25428 28226
rect 25025 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 25025 28072 25428 28108
rect 463 27760 946 28000
rect 463 27520 863 27760
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 863 27520
rect 463 27402 863 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 863 27402
rect 463 27061 863 27326
rect 25028 27520 25428 28072
rect 25028 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 25028 27402 25428 27444
rect 25028 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 953 27120 1155 27121
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 25294 863 26701
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24668 862 24885
rect 944 24681 946 24880
rect 463 24608 863 24668
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 863 24608
rect 463 24490 863 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 863 24490
rect 463 24238 863 24414
rect 25028 24559 25428 27326
rect 25028 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 25028 24441 25428 24483
rect 25028 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 463 24209 946 24238
rect 25028 24232 25428 24365
rect 462 23979 946 24209
rect 463 23760 946 23979
rect 24946 23766 25428 24232
rect 463 23604 863 23760
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 863 23604
rect 463 23486 863 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 863 23486
rect 25028 23467 25428 23766
rect 463 23060 863 23410
rect 25027 23442 25428 23467
rect 25027 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25428 23442
rect 25027 23324 25428 23366
rect 25027 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25428 23324
rect 25027 23212 25428 23248
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 21300 863 22700
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20651 863 20940
rect 463 20626 864 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 864 20626
rect 463 20508 864 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 864 20508
rect 463 20396 864 20432
rect 25028 20599 25428 23212
rect 25028 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 25028 20481 25428 20523
rect 25028 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 463 20239 863 20396
rect 463 19759 947 20239
rect 25028 20232 25428 20405
rect 24946 19767 25428 20232
rect 463 19569 863 19759
rect 463 19544 864 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 864 19544
rect 463 19426 864 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 864 19426
rect 463 19314 864 19350
rect 25028 19424 25428 19767
rect 25028 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 463 19060 863 19314
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 17301 863 18700
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16694 863 16941
rect 25028 19306 25428 19348
rect 25028 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 463 16669 864 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 864 16669
rect 25028 16608 25428 19230
rect 463 16551 864 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 864 16551
rect 463 16439 864 16475
rect 25027 16583 25428 16608
rect 25027 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25428 16583
rect 25027 16465 25428 16507
rect 463 16240 863 16439
rect 25027 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25428 16465
rect 25027 16353 25428 16389
rect 463 15760 946 16240
rect 25028 16233 25428 16353
rect 24946 15768 25428 16233
rect 463 15593 863 15760
rect 463 15568 864 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 864 15568
rect 463 15450 864 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 864 15450
rect 25028 15437 25428 15768
rect 463 15338 864 15374
rect 25027 15412 25428 15437
rect 463 15060 863 15338
rect 25027 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25428 15412
rect 25027 15294 25428 15336
rect 25027 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25428 15294
rect 25027 15182 25428 15218
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 13300 863 14700
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12727 863 12940
rect 463 12702 865 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 865 12702
rect 25028 12676 25428 15182
rect 463 12584 865 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 865 12584
rect 463 12472 865 12508
rect 25027 12651 25428 12676
rect 25027 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25428 12651
rect 25027 12533 25428 12575
rect 463 12239 863 12472
rect 25027 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25428 12533
rect 25027 12421 25428 12457
rect 463 11759 946 12239
rect 25028 12232 25428 12421
rect 24946 11766 25428 12232
rect 463 11511 863 11759
rect 463 11486 866 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 866 11486
rect 25028 11462 25428 11766
rect 463 11368 866 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 866 11368
rect 463 11256 866 11292
rect 25027 11437 25428 11462
rect 25027 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25428 11437
rect 25027 11319 25428 11361
rect 463 11060 863 11256
rect 25027 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25428 11319
rect 25027 11207 25428 11243
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 9300 863 10700
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8646 863 8940
rect 463 8621 864 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 864 8621
rect 463 8503 864 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 864 8503
rect 463 8391 864 8427
rect 25028 8594 25428 11207
rect 25028 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 25028 8476 25428 8518
rect 25028 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 463 8238 863 8391
rect 463 7998 947 8238
rect 25028 8233 25428 8400
rect 463 7758 946 7998
rect 24946 7766 25428 8233
rect 463 7524 863 7758
rect 463 7499 864 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 864 7499
rect 25028 7462 25428 7766
rect 463 7381 864 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 864 7381
rect 463 7269 864 7305
rect 25027 7437 25428 7462
rect 25027 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25428 7437
rect 25027 7319 25428 7361
rect 463 7061 863 7269
rect 25027 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25428 7319
rect 25027 7207 25428 7243
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 5299 863 6701
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4639 863 4939
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 863 4639
rect 463 4521 863 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 863 4521
rect 463 4238 863 4445
rect 25028 4594 25428 7207
rect 25028 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 25028 4476 25428 4518
rect 25028 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 463 4000 946 4238
rect 25028 4233 25428 4400
rect 463 3760 947 4000
rect 24946 3766 25428 4233
rect 463 3528 863 3760
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 25028 3462 25428 3766
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3061 863 3334
rect 25027 3437 25428 3462
rect 25027 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25428 3437
rect 25027 3319 25428 3361
rect 25027 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25428 3319
rect 25027 3207 25428 3243
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 1300 863 2701
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 730 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 25028 594 25428 3207
rect 25028 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 25028 476 25428 518
rect 463 239 863 475
rect 25028 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 463 0 947 239
rect 25028 233 25428 400
rect 24946 0 25428 233
rect 25502 35726 25902 68000
rect 25502 35646 25535 35726
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 25502 35606 25902 35646
rect 25502 35526 25534 35606
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 25502 33476 25902 35526
rect 25502 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 25502 33356 25902 33396
rect 25502 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 25502 0 25902 33276
rect 25970 66071 26370 68000
rect 25970 65995 26010 66071
rect 26082 65995 26136 66071
rect 26208 65995 26256 66071
rect 26328 65995 26370 66071
rect 25970 65953 26370 65995
rect 25970 65877 26010 65953
rect 26082 65877 26136 65953
rect 26208 65877 26256 65953
rect 26328 65877 26370 65953
rect 25970 62058 26370 65877
rect 25970 61982 26010 62058
rect 26082 61982 26136 62058
rect 26208 61982 26256 62058
rect 26328 61982 26370 62058
rect 25970 61940 26370 61982
rect 25970 61864 26010 61940
rect 26082 61864 26136 61940
rect 26208 61864 26256 61940
rect 26328 61864 26370 61940
rect 25970 58057 26370 61864
rect 25970 57981 26010 58057
rect 26082 57981 26136 58057
rect 26208 57981 26256 58057
rect 26328 57981 26370 58057
rect 25970 57939 26370 57981
rect 25970 57863 26010 57939
rect 26082 57863 26136 57939
rect 26208 57863 26256 57939
rect 26328 57863 26370 57939
rect 25970 54096 26370 57863
rect 25970 54020 26010 54096
rect 26082 54020 26136 54096
rect 26208 54020 26256 54096
rect 26328 54020 26370 54096
rect 25970 53978 26370 54020
rect 25970 53902 26010 53978
rect 26082 53902 26136 53978
rect 26208 53902 26256 53978
rect 26328 53902 26370 53978
rect 25970 50079 26370 53902
rect 25970 50003 26010 50079
rect 26082 50003 26136 50079
rect 26208 50003 26256 50079
rect 26328 50003 26370 50079
rect 25970 49961 26370 50003
rect 25970 49885 26010 49961
rect 26082 49885 26136 49961
rect 26208 49885 26256 49961
rect 26328 49885 26370 49961
rect 25970 46158 26370 49885
rect 25970 46082 26010 46158
rect 26082 46082 26136 46158
rect 26208 46082 26256 46158
rect 26328 46082 26370 46158
rect 25970 46040 26370 46082
rect 25970 45964 26010 46040
rect 26082 45964 26136 46040
rect 26208 45964 26256 46040
rect 26328 45964 26370 46040
rect 25970 41900 26370 45964
rect 25970 41824 26010 41900
rect 26082 41824 26136 41900
rect 26208 41824 26256 41900
rect 26328 41824 26370 41900
rect 25970 41782 26370 41824
rect 25970 41706 26010 41782
rect 26082 41706 26136 41782
rect 26208 41706 26256 41782
rect 26328 41706 26370 41782
rect 25970 26130 26370 41706
rect 25970 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 25970 26012 26370 26054
rect 25970 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 25970 21971 26370 25936
rect 25970 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 25970 21853 26370 21895
rect 25970 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 25970 18181 26370 21777
rect 25970 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 25970 18063 26370 18105
rect 25970 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 25970 14074 26370 17987
rect 25970 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 25970 13956 26370 13998
rect 25970 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 25970 10256 26370 13880
rect 25970 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 25970 10138 26370 10180
rect 25970 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 25970 6292 26370 10062
rect 25970 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 25970 6174 26370 6216
rect 25970 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 25970 2280 26370 6098
rect 25970 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 25970 2162 26370 2204
rect 25970 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 25970 0 26370 2086
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0
array 0 3 4000 0 0 4000
timestamp 1663849571
transform 1 0 8527 0 1 31332
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 5 4000 0 6 4000
timestamp 1663849571
transform 1 0 946 0 1 0
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_3
array 0 5 4000 0 6 4000
timestamp 1663849571
transform 1 0 946 0 1 40000
box 0 0 4000 4000
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_0
timestamp 1663599054
transform 1 0 2655 0 1 35031
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_1
timestamp 1663599054
transform 1 0 2210 0 1 35031
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_2
timestamp 1663599054
transform 1 0 2612 0 1 32975
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_3
timestamp 1663599054
transform 1 0 2132 0 1 32975
box -187 -76 187 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_4
timestamp 1663599054
transform 1 0 1779 0 -1 35031
box -187 -76 187 76
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_0
timestamp 1664545144
transform 1 0 2655 0 1 34693
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_1
timestamp 1664545144
transform 1 0 2210 0 1 34692
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_2
timestamp 1664545144
transform 1 0 2612 0 1 33213
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_3
timestamp 1664545144
transform 1 0 2132 0 1 33213
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_4
timestamp 1664545144
transform 1 0 1779 0 -1 34794
box -224 -36 223 138
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 4169 0 -1 35091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_1
timestamp 1662439860
transform -1 0 3617 0 -1 35091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_2
timestamp 1662439860
transform -1 0 4169 0 1 32915
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_3
timestamp 1662439860
transform -1 0 3617 0 1 32915
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1961 0 1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_1
timestamp 1662439860
transform 1 0 1961 0 -1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_2
timestamp 1662439860
transform 1 0 2881 0 1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_3
timestamp 1662439860
transform 1 0 3801 0 1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_4
timestamp 1662439860
transform 1 0 2881 0 -1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_5
timestamp 1662439860
transform 1 0 3801 0 -1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 4721 0 -1 35091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1662439860
transform -1 0 4721 0 1 32915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1662439860
transform -1 0 4445 0 -1 35091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1662439860
transform -1 0 4445 0 1 32915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1662439860
transform 1 0 1409 0 -1 34003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 1961 0 1 34003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1662439860
transform 1 0 1685 0 -1 34003
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1593 0 1 34003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1662439860
transform -1 0 3065 0 -1 35091
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1662439860
transform -1 0 3065 0 1 32915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1662439860
transform 1 0 1317 0 -1 34003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1662439860
transform 1 0 1501 0 1 32915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1662439860
transform 1 0 1420 0 -1 35092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1662439860
transform 1 0 4721 0 1 34003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1662439860
transform 1 0 4721 0 -1 34003
box -38 -48 130 592
<< labels >>
flabel metal4 s 0 0 400 68000 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 463 0 863 68000 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 25502 0 25902 68000 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 25028 0 25428 68000 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 2306 35775 2467 36000 0 FreeSans 480 90 0 0 mimtop1
flabel locali 1339 34217 1373 34269 0 FreeSans 800 0 0 0 clk
port 3 nsew signal input
flabel metal1 2919 33023 2956 33058 0 FreeSans 320 180 0 0 phi2
flabel metal1 2900 34829 2937 34876 0 FreeSans 320 180 0 0 phi1_n
flabel metal1 2927 33131 2964 33178 0 FreeSans 320 180 0 0 phi2_n
flabel metal1 2899 34946 2935 34981 0 FreeSans 320 180 0 0 phi1
flabel metal4 2493 28001 2737 28321 0 FreeSans 480 90 0 0 mimtop2
flabel metal4 25970 0 26370 64000 0 FreeSans 1600 90 0 0 vcm
port 4 nsew signal output
flabel metal4 4189 35754 4348 36000 0 FreeSans 480 90 0 0 mimbot1
<< properties >>
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
