magic
tech sky130A
timestamp 1666978453
<< metal1 >>
rect 12 10 4950 3471
<< properties >>
string FIXED_BBOX 0 0 5000 3500
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
