VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO emptybox_45_45
  CLASS BLOCK ;
  FOREIGN emptybox_45_45 ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.000 BY 45.000 ;
  OBS
      LAYER met1 ;
        RECT 0 0 45 45 ;
  END
END emptybox_45_45
END LIBRARY

