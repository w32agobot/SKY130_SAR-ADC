** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_top_postlayout_tb.sch
**.subckt adc_top_postlayout_tb
V_VDD_1 VDD GND pwl 0 0 {boot} 1.8
V_VCM_2 vmid GND pwl 0 0 {boot} 0.9
V_VCM_1 inp vmid pwl 0 0 {boot} {vdiff/2}
V_VCM_3 vmid inn pwl 0 0 {boot} {vdiff/2}
V_VCM clk_vcm GND 0 pulse(0 1.8 {0.5/fclk} 1n 1n {0.5/fclk} {1/fclk})
V1 rst_n GND pwl 0 0 390025n 0 390026n 1.8
V31 start_conv GND pwl 0 0 400025n 0 400026n 1.8 400525n 1.8 400526n 0 401300n 0 401326n 1.8 401825n
+ 1.8 401826n 0 402600n 0 402626n 1.8 403125n 1.8 403126n 0 403900n 0 403926n 1.8 404425n 1.8 404426n 0
V4 dlyctrl1_4 GND pwl 0 0 {boot} {bit4}
V5 dlyctrl1_3 GND pwl 0 0 {boot} {bit3}
V6 dlyctrl1_2 GND pwl 0 0 {boot} {bit2}
V7 dlyctrl1_1 GND pwl 0 0 {boot} {bit1}
V8 dlyctrl1_0 GND pwl 0 0 {boot} {bit0}
V2 avg_mode2 GND pwl 0 0 {boot} {avg2}
V3 avg_mode1 GND pwl 0 0 {boot} {avg1}
V25 avg_mode0 GND pwl 0 0 {boot} {avg0}
V19 dlyctrl4_5 GND pwl 0 0 {boot} {ed_bit5}
V20 dlyctrl4_4 GND pwl 0 0 {boot} {ed_bit4}
V21 dlyctrl4_3 GND pwl 0 0 {boot} {ed_bit3}
V22 dlyctrl4_2 GND pwl 0 0 {boot} {ed_bit2}
V23 dlyctrl4_1 GND pwl 0 0 {boot} {ed_bit1}
V24 dlyctrl4_0 GND pwl 0 0 {boot} {ed_bit0}
V26 en_dly_contr GND pwl 0 0 {boot} {dlyctrl}
V27 osr_mode2 GND pwl 0 0 {boot} {osr2}
V28 osr_mode1 GND pwl 0 0 {boot} {osr1}
V29 osr_mode0 GND pwl 0 0 {boot} {osr0}
V30 nc0 GND 0
x1 result0 result1 result2 result3 result4 result5 result6 result7 result8 result9 result10 result11
+ result12 result13 result14 result15 VDD GND conv_finished rst_n start_conv clk_vcm inp inn avg_mode0
+ avg_mode1 avg_mode2 osr_mode0 osr_mode1 osr_mode2 row_mode col_mode nc0 nc1 dlyctrl4_0 dlyctrl4_1 dlyctrl4_2
+ dlyctrl4_3 dlyctrl4_4 dlyctrl4_5 dlyctrl1_0 dlyctrl1_1 dlyctrl1_2 dlyctrl1_3 dlyctrl1_4 dlyctrl2_0 dlyctrl2_1
+ dlyctrl2_2 dlyctrl2_3 dlyctrl2_4 dlyctrl3_0 dlyctrl3_1 dlyctrl3_2 dlyctrl3_3 dlyctrl3_4 en_dly_contr net1[15]
+ net1[14] net1[13] net1[12] net1[11] net1[10] net1[9] net1[8] net1[7] net1[6] net1[5] net1[4] net1[3] net1[2]
+ net1[1] net1[0] ctopp ctopn vcm clk_dig clk_comp clk_ena ndecision_finish comp_latch conv_finished_osr
+ adc_top_postlayout
V9 dlyctrl2_4 GND pwl 0 0 {boot} {bit4}
V10 dlyctrl2_3 GND pwl 0 0 {boot} {bit3}
V11 dlyctrl2_2 GND pwl 0 0 {boot} {bit2}
V12 dlyctrl2_1 GND pwl 0 0 {boot} {bit1}
V13 dlyctrl2_0 GND pwl 0 0 {boot} {bit0}
V14 dlyctrl3_4 GND pwl 0 0 {boot} {bit4}
V15 dlyctrl3_3 GND pwl 0 0 {boot} {bit3}
V16 dlyctrl3_2 GND pwl 0 0 {boot} {bit2}
V17 dlyctrl3_1 GND pwl 0 0 {boot} {bit1}
V18 dlyctrl3_0 GND pwl 0 0 {boot} {bit0}
V32 GND 0 0
V33 row_mode GND pwl 0 0 {boot} {rowmode}
V34 col_mode GND pwl 0 0 {boot} {colmode}
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt





* xyce commands
.include ../../spice/adc_top.gds.C.noD.merge.postlayout.spice

****************
* Misc
****************
.param fclk=32768
.param vdiff=200m
.param boot=100n

****************
* Delay Config
****************
.param dlyctrl = 1.8

* delay 1-3
.param bit0 = 1.8
.param bit1 = 0
.param bit2 = 0
.param bit3 = 0
.param bit4 = 0

* edgedetect pulse
.param ed_bit0 = 0
.param ed_bit1 = 1.8
.param ed_bit2 = 1.8
.param ed_bit3 = 0
.param ed_bit4 = 0
.param ed_bit5 = 0

****************
* Averaging Config
****************
.param avg0 = 1.8
.param avg1 = 0
.param avg2 = 0

****************
* OSR Config
****************
.param osr0 = 1.8
.param osr1 = 0
.param osr2 = 0


****************
* Row Column
* sequential or symmetric
****************
.param rowmode = 1.8
.param colmode = 1.8


****************
* XYCE Simulation Control
****************

*.options linsol type=klu
*.OPTIONS TIMEINT BREAKPOINTS=610us,611us,612us
.OPTIONS TIMEINT ABSTOL=1e-8 RELTOL=1e-4
.tran 1n 420u uic

.print tran format=raw file=adc_top_postlayout_tb.raw         v(x1:ctopp) v(x1:ctopn) v(x1:vcm)
+ v(x1:clk_ena) v(x1:ndecision_finish) v(x1:comp_latch) v(VDD) v(rst_n) v(start_conv) v(clk_vcm) v(inp) v(inn)
+ v(conv_finished) v(conv_finished_osr) v(x1:clk_dig) v(x1:clk_comp) v(result*) v(dlyctrl*) v(avg_mode*) v(osr_mode*)
+ v(en_dly_contr) i(v_vdd_1) v(x1:sh_switch_pmat) v(x1:sh_switch_pmat_n) v(x1:sample_pmat_n) v(x1:sample_pmat_n_int)
+ v(x1:sample_pmat_int)
.print tran format=std file=adc_top_postlayout_tb.ascii       v(x1:ctopp) v(x1:ctopn) v(x1:vcm)
+ v(x1:clk_ena) v(x1:ndecision_finish) v(x1:comp_latch) v(VDD) v(rst_n) v(start_conv) v(clk_vcm) v(inp) v(inn)
+ v(conv_finished) v(conv_finished_osr) v(x1:clk_dig) v(x1:clk_comp) v(result*) v(dlyctrl*) v(avg_mode*) v(osr_mode*)
+ v(en_dly_contr) i(v_vdd_1) v(x1:sh_switch_pmat) v(x1:sh_switch_pmat_n) v(x1:sample_pmat_n) v(x1:sample_pmat_n_int)
+ v(x1:sample_pmat_int)
.print tran format=csv file=adc_top_postlayout_tb.csv         v(x1:ctopp) v(x1:ctopn) v(x1:vcm)
+ v(x1:clk_ena) v(x1:ndecision_finish) v(x1:comp_latch) v(VDD) v(rst_n) v(start_conv) v(clk_vcm) v(inp) v(inn)
+ v(conv_finished) v(conv_finished_osr) v(x1:clk_dig) v(x1:clk_comp) v(result*) v(dlyctrl*) v(avg_mode*) v(osr_mode*)
+ v(en_dly_contr) i(v_vdd_1)  v(x1:sh_switch_pmat) v(x1:sh_switch_pmat_n) v(x1:sample_pmat_n) v(x1:sample_pmat_n_int)
+ v(x1:sample_pmat_int)
.print tran format=gnuplot file=adc_top_postlayout_tb.gnu.dat v(x1:ctopp) v(x1:ctopn) v(x1:vcm)
+ v(x1:clk_ena) v(x1:ndecision_finish) v(x1:comp_latch) v(VDD) v(rst_n) v(start_conv) v(clk_vcm) v(inp) v(inn)
+ v(conv_finished) v(conv_finished_osr) v(x1:clk_dig) v(x1:clk_comp) v(result*) v(dlyctrl*) v(avg_mode*) v(osr_mode*)
+ v(en_dly_contr) i(v_vdd_1)  v(x1:sh_switch_pmat) v(x1:sh_switch_pmat_n) v(x1:sample_pmat_n) v(x1:sample_pmat_n_int)
+ v(x1:sample_pmat_int)








**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
