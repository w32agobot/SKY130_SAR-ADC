magic
tech sky130A
timestamp 1660640026
<< checkpaint >>
rect -310 988 1617 1110
rect -661 -612 1617 988
rect -661 -734 1266 -612
<< metal2 >>
rect 8 220 622 280
rect 8 192 13 220
rect 41 192 77 220
rect 105 192 141 220
rect 169 192 205 220
rect 233 192 269 220
rect 297 192 333 220
rect 361 192 397 220
rect 425 192 461 220
rect 489 192 525 220
rect 553 192 589 220
rect 617 192 622 220
rect 8 134 622 192
rect 8 106 13 134
rect 41 106 77 134
rect 105 106 141 134
rect 169 106 205 134
rect 233 106 269 134
rect 297 106 333 134
rect 361 106 397 134
rect 425 106 461 134
rect 489 106 525 134
rect 553 106 589 134
rect 617 106 622 134
rect 8 48 622 106
rect 8 20 13 48
rect 41 20 77 48
rect 105 20 141 48
rect 169 20 205 48
rect 233 20 269 48
rect 297 20 333 48
rect 361 20 397 48
rect 425 20 461 48
rect 489 20 525 48
rect 553 20 589 48
rect 617 20 622 48
rect 8 -40 622 20
<< via2 >>
rect 13 192 41 220
rect 77 192 105 220
rect 141 192 169 220
rect 205 192 233 220
rect 269 192 297 220
rect 333 192 361 220
rect 397 192 425 220
rect 461 192 489 220
rect 525 192 553 220
rect 589 192 617 220
rect 13 106 41 134
rect 77 106 105 134
rect 141 106 169 134
rect 205 106 233 134
rect 269 106 297 134
rect 333 106 361 134
rect 397 106 425 134
rect 461 106 489 134
rect 525 106 553 134
rect 589 106 617 134
rect 13 20 41 48
rect 77 20 105 48
rect 141 20 169 48
rect 205 20 233 48
rect 269 20 297 48
rect 333 20 361 48
rect 397 20 425 48
rect 461 20 489 48
rect 525 20 553 48
rect 589 20 617 48
<< metal3 >>
rect 10 220 44 259
rect 10 192 13 220
rect 41 192 44 220
rect 10 134 44 192
rect 10 106 13 134
rect 41 106 44 134
rect 10 48 44 106
rect 10 20 13 48
rect 41 20 44 48
rect 10 -19 44 20
rect 74 220 108 259
rect 74 192 77 220
rect 105 192 108 220
rect 74 134 108 192
rect 74 106 77 134
rect 105 106 108 134
rect 74 48 108 106
rect 74 20 77 48
rect 105 20 108 48
rect 74 -19 108 20
rect 138 220 172 259
rect 138 192 141 220
rect 169 192 172 220
rect 138 134 172 192
rect 138 106 141 134
rect 169 106 172 134
rect 138 48 172 106
rect 138 20 141 48
rect 169 20 172 48
rect 138 -19 172 20
rect 202 220 236 259
rect 202 192 205 220
rect 233 192 236 220
rect 202 134 236 192
rect 202 106 205 134
rect 233 106 236 134
rect 202 48 236 106
rect 202 20 205 48
rect 233 20 236 48
rect 202 -19 236 20
rect 266 220 300 259
rect 266 192 269 220
rect 297 192 300 220
rect 266 134 300 192
rect 266 106 269 134
rect 297 106 300 134
rect 266 48 300 106
rect 266 20 269 48
rect 297 20 300 48
rect 266 -19 300 20
rect 330 220 364 259
rect 330 192 333 220
rect 361 192 364 220
rect 330 134 364 192
rect 330 106 333 134
rect 361 106 364 134
rect 330 48 364 106
rect 330 20 333 48
rect 361 20 364 48
rect 330 -19 364 20
rect 394 220 428 259
rect 394 192 397 220
rect 425 192 428 220
rect 394 134 428 192
rect 394 106 397 134
rect 425 106 428 134
rect 394 48 428 106
rect 394 20 397 48
rect 425 20 428 48
rect 394 -19 428 20
rect 458 220 492 259
rect 458 192 461 220
rect 489 192 492 220
rect 458 134 492 192
rect 458 106 461 134
rect 489 106 492 134
rect 458 48 492 106
rect 458 20 461 48
rect 489 20 492 48
rect 458 -19 492 20
rect 522 220 556 259
rect 522 192 525 220
rect 553 192 556 220
rect 522 134 556 192
rect 522 106 525 134
rect 553 106 556 134
rect 522 48 556 106
rect 522 20 525 48
rect 553 20 556 48
rect 522 -19 556 20
rect 586 220 620 259
rect 586 192 589 220
rect 617 192 620 220
rect 586 134 620 192
rect 586 106 589 134
rect 617 106 620 134
rect 586 48 620 106
rect 586 20 589 48
rect 617 20 620 48
rect 586 -19 620 20
<< metal4 >>
rect -6 295 636 310
rect 12 -25 42 265
rect 76 -55 106 295
rect 140 -55 170 295
rect 204 -55 234 295
rect 268 -55 298 295
rect 332 -55 362 295
rect 396 -55 426 295
rect 460 -55 490 295
rect 524 -55 554 295
rect 588 -25 618 265
rect -6 -70 636 -55
<< end >>
