* SPICE3 file created from extract.ext - technology: sky130A

C0 bot_8 dummy_bot 8.02fF
C1 bot_1 top_1 34.30fF
C2 dummy_bot dummy-top 294.60fF
C3 bot_8 top_8 33.34fF
C4 dummy_bot top_8 2.41fF
C5 top_8 dummy-top 3.20fF
C6 dummy_bot top_2 2.25fF
C7 dummy_bot top_4 2.32fF
C8 m3_15766_216# bot_1 2.49fF
C9 dummy-top top_2 3.05fF
C10 dummy_bot bot_2 9.02fF
C11 dummy-top top_4 3.20fF
C12 dummy_bot bot_4 9.02fF
C13 dummy_bot bot_1 9.01fF
C14 bot_2 top_2 34.91fF
C15 dummy_bot top_1 2.17fF
C16 bot_4 top_4 36.16fF
C17 dummy-top top_1 2.96fF
C18 dummy-top VSUBS 6.70fF
C19 bot_1 VSUBS 3.90fF
C20 bot_2 VSUBS 3.90fF
C21 bot_4 VSUBS 3.90fF
C22 bot_8 VSUBS 3.05fF
C23 dummy_bot VSUBS 41.48fF
